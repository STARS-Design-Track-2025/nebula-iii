* NGSPICE file created from team_05.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_40_12 abstract view
.subckt sky130_ef_sc_hd__decap_40_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_4 abstract view
.subckt sky130_fd_sc_hd__fill_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_8 abstract view
.subckt sky130_fd_sc_hd__fill_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_1 abstract view
.subckt sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_1 abstract view
.subckt sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

.subckt team_05 ACK_I ADR_O[0] ADR_O[10] ADR_O[11] ADR_O[12] ADR_O[13] ADR_O[14] ADR_O[15]
+ ADR_O[16] ADR_O[17] ADR_O[18] ADR_O[19] ADR_O[1] ADR_O[20] ADR_O[21] ADR_O[22] ADR_O[23]
+ ADR_O[24] ADR_O[25] ADR_O[26] ADR_O[27] ADR_O[28] ADR_O[29] ADR_O[2] ADR_O[30] ADR_O[31]
+ ADR_O[3] ADR_O[4] ADR_O[5] ADR_O[6] ADR_O[7] ADR_O[8] ADR_O[9] CYC_O DAT_I[0] DAT_I[10]
+ DAT_I[11] DAT_I[12] DAT_I[13] DAT_I[14] DAT_I[15] DAT_I[16] DAT_I[17] DAT_I[18]
+ DAT_I[19] DAT_I[1] DAT_I[20] DAT_I[21] DAT_I[22] DAT_I[23] DAT_I[24] DAT_I[25] DAT_I[26]
+ DAT_I[27] DAT_I[28] DAT_I[29] DAT_I[2] DAT_I[30] DAT_I[31] DAT_I[3] DAT_I[4] DAT_I[5]
+ DAT_I[6] DAT_I[7] DAT_I[8] DAT_I[9] DAT_O[0] DAT_O[10] DAT_O[11] DAT_O[12] DAT_O[13]
+ DAT_O[14] DAT_O[15] DAT_O[16] DAT_O[17] DAT_O[18] DAT_O[19] DAT_O[1] DAT_O[20] DAT_O[21]
+ DAT_O[22] DAT_O[23] DAT_O[24] DAT_O[25] DAT_O[26] DAT_O[27] DAT_O[28] DAT_O[29]
+ DAT_O[2] DAT_O[30] DAT_O[31] DAT_O[3] DAT_O[4] DAT_O[5] DAT_O[6] DAT_O[7] DAT_O[8]
+ DAT_O[9] SEL_O[0] SEL_O[1] SEL_O[2] SEL_O[3] STB_O WE_O clk en gpio_in[0] gpio_in[10]
+ gpio_in[11] gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17]
+ gpio_in[18] gpio_in[19] gpio_in[1] gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23]
+ gpio_in[24] gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2]
+ gpio_in[30] gpio_in[31] gpio_in[32] gpio_in[33] gpio_in[3] gpio_in[4] gpio_in[5]
+ gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9] gpio_oeb[0] gpio_oeb[10] gpio_oeb[11]
+ gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15] gpio_oeb[16] gpio_oeb[17] gpio_oeb[18]
+ gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21] gpio_oeb[22] gpio_oeb[23] gpio_oeb[24]
+ gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28] gpio_oeb[29] gpio_oeb[2] gpio_oeb[30]
+ gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[3] gpio_oeb[4] gpio_oeb[5] gpio_oeb[6]
+ gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12]
+ gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19]
+ gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25]
+ gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31]
+ gpio_out[32] gpio_out[33] gpio_out[3] gpio_out[4] gpio_out[5] gpio_out[6] gpio_out[7]
+ gpio_out[8] gpio_out[9] nrst vccd1 vssd1
X_05903_ top.sram_interface.CB_write_counter\[1\] _02452_ _02857_ top.CB_write_complete
+ vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__a31o_1
X_09671_ net785 net625 vssd1 vssd1 vccd1 vccd1 _00285_ sky130_fd_sc_hd__and2_1
X_06883_ top.findLeastValue.val2\[42\] net150 net123 _03583_ vssd1 vssd1 vccd1 vccd1
+ _01984_ sky130_fd_sc_hd__o22a_1
X_08622_ top.cb_syn.num_lefts\[4\] _04829_ top.cb_syn.num_lefts\[5\] vssd1 vssd1 vccd1
+ vccd1 _04839_ sky130_fd_sc_hd__a21o_1
X_05834_ net452 _02843_ _02844_ _02780_ vssd1 vssd1 vccd1 vccd1 _02845_ sky130_fd_sc_hd__a211o_1
XANTENNA__05545__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06928__S net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08553_ net1306 top.cb_syn.char_path_n\[23\] net229 vssd1 vssd1 vccd1 vccd1 _01541_
+ sky130_fd_sc_hd__mux2_1
X_05765_ top.translation.resEn top.translation.totalEn vssd1 vssd1 vccd1 vccd1 _02786_
+ sky130_fd_sc_hd__or2_1
X_08484_ net1075 top.cb_syn.char_path_n\[92\] net234 vssd1 vssd1 vccd1 vccd1 _01610_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_85_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05560__A3 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07504_ _04091_ _04092_ _04093_ _04094_ _04072_ _04071_ vssd1 vssd1 vccd1 vccd1 _04095_
+ sky130_fd_sc_hd__mux4_1
X_07435_ _04026_ _04030_ net404 vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__mux2_1
X_05696_ net18 net417 net359 top.WB.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1 _02362_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__05848__B2 top.WB.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09039__A1 top.WB.CPU_DAT_O\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07366_ net499 _03553_ _03975_ vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_33_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09105_ _05123_ _05124_ _03323_ vssd1 vssd1 vccd1 vccd1 _00044_ sky130_fd_sc_hd__or3b_1
XANTENNA__08798__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07297_ _03797_ _03930_ vssd1 vssd1 vccd1 vccd1 _03931_ sky130_fd_sc_hd__nand2_1
X_06317_ top.hist_data_o\[10\] top.hist_data_o\[9\] _03179_ vssd1 vssd1 vccd1 vccd1
+ _03180_ sky130_fd_sc_hd__and3_1
XFILLER_108_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_06248_ top.cw1\[3\] top.cw1\[2\] top.cw1\[1\] top.cw1\[0\] vssd1 vssd1 vccd1 vccd1
+ _03115_ sky130_fd_sc_hd__and4_1
X_09036_ net1371 top.WB.CPU_DAT_O\[21\] net291 vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout796_A net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06179_ _02946_ _03048_ vssd1 vssd1 vccd1 vccd1 _03049_ sky130_fd_sc_hd__nor2_1
XFILLER_89_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold362 top.hTree.tree_reg\[63\] vssd1 vssd1 vccd1 vccd1 net1315 sky130_fd_sc_hd__dlygate4sd3_1
Xhold340 top.hTree.node_reg\[43\] vssd1 vssd1 vccd1 vccd1 net1293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold351 top.cb_syn.char_path\[45\] vssd1 vssd1 vccd1 vccd1 net1304 sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 net63 vssd1 vssd1 vccd1 vccd1 net1326 sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 top.path\[47\] vssd1 vssd1 vccd1 vccd1 net1337 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07347__X _03966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06025__A1 top.WB.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold395 top.cb_syn.char_path\[42\] vssd1 vssd1 vccd1 vccd1 net1348 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09938_ net787 net627 vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__and2_1
XANTENNA__07773__A1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout842 net879 vssd1 vssd1 vccd1 vccd1 net842 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout584_X net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout820 net823 vssd1 vssd1 vccd1 vccd1 net820 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout831 net835 vssd1 vssd1 vccd1 vccd1 net831 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08970__A0 top.WB.CPU_DAT_O\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout875 net876 vssd1 vssd1 vccd1 vccd1 net875 sky130_fd_sc_hd__buf_1
Xfanout853 net857 vssd1 vssd1 vccd1 vccd1 net853 sky130_fd_sc_hd__clkbuf_2
Xfanout864 net865 vssd1 vssd1 vccd1 vccd1 net864 sky130_fd_sc_hd__clkbuf_2
XFILLER_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09869_ net778 net618 vssd1 vssd1 vccd1 vccd1 _00483_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout849_X net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05536__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11831_ clknet_leaf_114_clk _02347_ _01186_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08338__B _02506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11762_ clknet_leaf_114_clk _02295_ _01117_ vssd1 vssd1 vccd1 vccd1 top.compVal\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11693_ clknet_leaf_61_clk _02226_ _01048_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_14_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05839__B2 top.WB.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10713_ clknet_leaf_3_clk _01312_ _00132_ vssd1 vssd1 vccd1 vccd1 top.path\[89\]
+ sky130_fd_sc_hd__dfrtp_1
X_10644_ clknet_leaf_49_clk _00039_ _00063_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.word_cnt\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10575_ net810 net650 vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__and2_1
XANTENNA__08789__B1 top.translation.index\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06264__B2 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06016__A1 top.WB.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11127_ clknet_leaf_30_clk _01675_ _00482_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[29\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08961__A0 top.WB.CPU_DAT_O\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11058_ clknet_leaf_26_clk _01606_ _00413_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[88\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05527__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10009_ net818 net658 vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__and2_1
XANTENNA__06781__B_N _03546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05542__A3 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05550_ net1432 net145 _02646_ net177 vssd1 vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__a22o_1
XFILLER_32_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05481_ top.WB.curr_state\[0\] _02544_ net212 vssd1 vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_50_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07220_ _03845_ _03872_ vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__nand2_1
XFILLER_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07151_ _03782_ _03808_ vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__or2_1
X_06102_ top.TRN_char_index\[3\] _02974_ vssd1 vssd1 vccd1 vccd1 _02975_ sky130_fd_sc_hd__and2_1
XFILLER_105_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07082_ top.findLeastValue.val1\[6\] top.findLeastValue.val2\[6\] vssd1 vssd1 vccd1
+ vccd1 _03740_ sky130_fd_sc_hd__or2_1
XANTENNA__10018__B net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09807__B net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06033_ top.hist_data_o\[2\] top.WB.CPU_DAT_O\[2\] net355 vssd1 vssd1 vccd1 vccd1
+ _02177_ sky130_fd_sc_hd__mux2_1
XANTENNA__06007__A1 top.WB.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08401__C1 top.cb_syn.end_cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout127 _03549_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__08952__A0 top.WB.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout138 net140 vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__buf_4
Xfanout116 net117 vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__clkbuf_2
X_07984_ _02513_ top.cb_syn.zero_count\[3\] top.cb_syn.zero_count\[4\] _02512_ vssd1
+ vssd1 vccd1 vccd1 _04487_ sky130_fd_sc_hd__a22o_1
XFILLER_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05773__D top.findLeastValue.least1\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout149 net151 vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__clkbuf_4
X_06935_ top.findLeastValue.val2\[16\] net146 net120 _03609_ vssd1 vssd1 vccd1 vccd1
+ _01958_ sky130_fd_sc_hd__o22a_1
X_09723_ net735 net575 vssd1 vssd1 vccd1 vccd1 _00337_ sky130_fd_sc_hd__and2_1
X_09654_ net798 net638 vssd1 vssd1 vccd1 vccd1 _00268_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout377_A net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06866_ net497 _03571_ _03577_ vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__o21ba_1
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08605_ net534 net540 top.cb_syn.curr_state\[8\] vssd1 vssd1 vccd1 vccd1 _04824_
+ sky130_fd_sc_hd__or3_1
X_05817_ _02821_ _02826_ top.sram_interface.counter_HTREE\[0\] vssd1 vssd1 vccd1 vccd1
+ _02834_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_38_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout544_A net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09585_ net822 net662 vssd1 vssd1 vccd1 vccd1 _00199_ sky130_fd_sc_hd__and2_1
X_06797_ top.findLeastValue.val1\[33\] net133 net117 top.compVal\[33\] vssd1 vssd1
+ vccd1 vccd1 _02041_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout165_X net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05748_ _02539_ net172 vssd1 vssd1 vccd1 vccd1 _02783_ sky130_fd_sc_hd__nor2_2
X_08536_ net1238 top.cb_syn.char_path_n\[40\] net226 vssd1 vssd1 vccd1 vccd1 _01558_
+ sky130_fd_sc_hd__mux2_1
X_05679_ top.cb_syn.char_path\[0\] net560 net315 top.cb_syn.char_path\[96\] vssd1
+ vssd1 vccd1 vccd1 _02754_ sky130_fd_sc_hd__a22o_1
X_08467_ net1313 top.cb_syn.char_path_n\[109\] net220 vssd1 vssd1 vccd1 vccd1 _01627_
+ sky130_fd_sc_hd__mux2_1
X_07418_ _04014_ _04016_ net354 vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__mux2_1
XFILLER_50_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_08398_ top.cb_syn.char_path_n\[9\] net393 net330 top.cb_syn.char_path_n\[10\] _02504_
+ vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_98_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_93_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07349_ _03763_ _03765_ vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__or2_1
X_10360_ net864 net704 vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__and2_1
X_10291_ net724 net564 vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__and2_1
X_09019_ top.WB.CPU_DAT_O\[6\] net1198 net320 vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__mux2_1
XANTENNA__06797__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_05_900 vssd1 vssd1 vccd1 vccd1 team_05_900/HI gpio_out[15] sky130_fd_sc_hd__conb_1
Xteam_05_911 vssd1 vssd1 vccd1 vccd1 team_05_911/HI gpio_out[26] sky130_fd_sc_hd__conb_1
Xhold170 top.path\[11\] vssd1 vssd1 vccd1 vccd1 net1123 sky130_fd_sc_hd__dlygate4sd3_1
Xteam_05_922 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] team_05_922/LO sky130_fd_sc_hd__conb_1
XANTENNA__08943__A0 top.WB.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold181 top.cb_syn.char_path\[3\] vssd1 vssd1 vccd1 vccd1 net1134 sky130_fd_sc_hd__dlygate4sd3_1
Xteam_05_944 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] team_05_944/LO sky130_fd_sc_hd__conb_1
Xteam_05_933 vssd1 vssd1 vccd1 vccd1 gpio_oeb[13] team_05_933/LO sky130_fd_sc_hd__conb_1
Xhold192 top.path\[65\] vssd1 vssd1 vccd1 vccd1 net1145 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_31_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout650 net651 vssd1 vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__clkbuf_2
Xfanout694 net695 vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__clkbuf_2
Xfanout683 net718 vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__clkbuf_2
Xfanout661 net663 vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__buf_1
Xfanout672 net674 vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__clkbuf_2
XANTENNA__05509__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05524__A3 _02583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_46_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11814_ clknet_leaf_47_clk net452 _01169_ vssd1 vssd1 vccd1 vccd1 top.WB.prev_BUSY_O
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08783__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11745_ clknet_leaf_94_clk _02278_ _01100_ vssd1 vssd1 vccd1 vccd1 top.compVal\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11676_ clknet_leaf_60_clk _02209_ _01031_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10627_ net805 net645 vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_104_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10558_ net870 net710 vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_58_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06788__A2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10489_ net830 net670 vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__and2_1
XANTENNA__08934__A0 top.WB.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_119_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07715__X _04278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06720_ _02421_ top.findLeastValue.val2\[29\] top.findLeastValue.val2\[28\] _02422_
+ vssd1 vssd1 vccd1 vccd1 _03508_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_69_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06651_ _03436_ _03438_ _03439_ vssd1 vssd1 vccd1 vccd1 _03440_ sky130_fd_sc_hd__nor3_1
X_05602_ _02454_ net459 net362 vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__and3_1
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_35_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09370_ net976 net238 net215 _04306_ vssd1 vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__a22o_1
X_06582_ _02434_ top.findLeastValue.val1\[15\] vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__and2_1
X_05533_ top.cb_syn.char_path\[88\] net553 net544 top.cb_syn.char_path\[56\] vssd1
+ vssd1 vccd1 vccd1 _02632_ sky130_fd_sc_hd__a22o_1
X_08321_ top.cb_syn.char_path_n\[9\] net378 net337 top.cb_syn.char_path_n\[7\] net182
+ vssd1 vssd1 vccd1 vccd1 _04688_ sky130_fd_sc_hd__a221o_1
X_05464_ net451 top.findLeastValue.wipe_the_char_2 net546 vssd1 vssd1 vccd1 vccd1
+ _02572_ sky130_fd_sc_hd__and3_2
XANTENNA__07673__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08252_ top.cb_syn.char_path_n\[43\] net195 _04653_ vssd1 vssd1 vccd1 vccd1 _01689_
+ sky130_fd_sc_hd__o21a_1
X_07203_ top.findLeastValue.val1\[45\] top.findLeastValue.val2\[45\] vssd1 vssd1 vccd1
+ vccd1 _03861_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_4_12_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_12_0_clk sky130_fd_sc_hd__clkbuf_8
X_05395_ top.cb_syn.end_cnt\[4\] vssd1 vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__inv_2
X_08183_ top.cb_syn.char_path_n\[78\] net374 net334 top.cb_syn.char_path_n\[76\] net179
+ vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__a221o_1
X_07134_ _03789_ _03790_ vssd1 vssd1 vccd1 vccd1 _03792_ sky130_fd_sc_hd__nor2_1
XANTENNA__07520__S0 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06779__A2 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07065_ _03722_ vssd1 vssd1 vccd1 vccd1 _03723_ sky130_fd_sc_hd__inv_2
X_06016_ net1704 top.WB.CPU_DAT_O\[19\] net357 vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_93_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06242__A top.findLeastValue.histo_index\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08925__A0 top.WB.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10760__Q top.cb_syn.h_element\[54\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07967_ top.findLeastValue.alternator_timer\[2\] top.findLeastValue.alternator_timer\[1\]
+ top.findLeastValue.alternator_timer\[0\] _04474_ vssd1 vssd1 vccd1 vccd1 _04475_
+ sky130_fd_sc_hd__a31oi_1
XANTENNA_fanout282_X net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09706_ net850 net690 vssd1 vssd1 vccd1 vccd1 _00320_ sky130_fd_sc_hd__and2_1
XANTENNA__06951__A2 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06918_ top.compVal\[24\] top.findLeastValue.val1\[24\] net163 vssd1 vssd1 vccd1
+ vccd1 _03601_ sky130_fd_sc_hd__mux2_1
XFILLER_114_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09350__B1 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07898_ net440 net1546 net251 top.findLeastValue.sum\[9\] _04424_ vssd1 vssd1 vccd1
+ vccd1 _01814_ sky130_fd_sc_hd__a221o_1
X_09637_ net801 net641 vssd1 vssd1 vccd1 vccd1 _00251_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout547_X net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05506__A3 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06849_ top.findLeastValue.least1\[0\] net504 _03424_ vssd1 vssd1 vccd1 vccd1 _03564_
+ sky130_fd_sc_hd__mux2_1
X_09568_ net843 net683 vssd1 vssd1 vccd1 vccd1 _00182_ sky130_fd_sc_hd__and2_1
XFILLER_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08519_ net1255 top.cb_syn.char_path_n\[57\] net232 vssd1 vssd1 vccd1 vccd1 _01575_
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_13_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09499_ net756 net596 vssd1 vssd1 vccd1 vccd1 _00113_ sky130_fd_sc_hd__and2_1
X_11530_ clknet_leaf_5_clk _02078_ _00885_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_102_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwire325 _05035_ vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__clkbuf_2
X_11461_ clknet_leaf_94_clk _02009_ _00816_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[1\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__06219__B2 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10412_ net794 net634 vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__and2_1
XANTENNA__05690__A2 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11392_ clknet_leaf_82_clk _01940_ _00747_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[44\]
+ sky130_fd_sc_hd__dfrtp_1
X_10343_ net854 net694 vssd1 vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__and2_1
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07511__S0 _04072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09169__B1 _02581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10274_ net727 net567 vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__and2_1
XFILLER_105_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08392__A1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout480 net481 vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__buf_4
Xfanout491 net492 vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_105_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11728_ clknet_leaf_121_clk _02261_ _01083_ vssd1 vssd1 vccd1 vccd1 top.path\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_104_Right_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11659_ clknet_leaf_14_clk _02192_ _01014_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05681__A2 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07958__A1 top.findLeastValue.least2\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07502__S0 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08870_ top.translation.index\[3\] _05048_ vssd1 vssd1 vccd1 vccd1 _05049_ sky130_fd_sc_hd__or2_1
XFILLER_69_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08383__A1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07821_ net484 _04361_ vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__or2_1
XANTENNA__07605__B _04187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07752_ net430 _04306_ _04307_ net260 vssd1 vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__o211a_1
X_07683_ net492 _04251_ vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__nand2_1
XANTENNA__07489__A3 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06703_ top.compVal\[22\] _02490_ _02491_ top.compVal\[21\] vssd1 vssd1 vccd1 vccd1
+ _03491_ sky130_fd_sc_hd__a22o_1
X_09422_ net966 _05291_ net245 vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06936__S net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07894__A0 top.findLeastValue.sum\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06634_ _03388_ _03413_ _03422_ vssd1 vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__a21oi_4
X_09353_ net1024 net241 net217 _04374_ vssd1 vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__a22o_1
X_08304_ top.cb_syn.char_path_n\[17\] net197 _04679_ vssd1 vssd1 vccd1 vccd1 _01663_
+ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout242_A net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06565_ _02440_ top.findLeastValue.val1\[9\] top.findLeastValue.val1\[8\] _02441_
+ vssd1 vssd1 vccd1 vccd1 _03354_ sky130_fd_sc_hd__o22a_1
X_09284_ _04000_ _04011_ _04034_ vssd1 vssd1 vccd1 vccd1 top.dut.bit_buf_next\[2\]
+ sky130_fd_sc_hd__o21a_1
X_05516_ top.cb_syn.char_path\[27\] net559 net314 top.cb_syn.char_path\[123\] vssd1
+ vssd1 vccd1 vccd1 _02618_ sky130_fd_sc_hd__a22o_1
X_06496_ net1630 _03283_ vssd1 vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__nor2_1
X_05447_ top.cb_syn.setup _02527_ _02554_ vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__or3_2
X_08235_ top.cb_syn.char_path_n\[52\] net375 net335 top.cb_syn.char_path_n\[50\] net180
+ vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout507_A net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08166_ top.cb_syn.char_path_n\[86\] net208 _04610_ vssd1 vssd1 vccd1 vccd1 _01732_
+ sky130_fd_sc_hd__o21a_1
X_05378_ top.findLeastValue.val2\[35\] vssd1 vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout128_X net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07117_ _03770_ _03772_ _03774_ vssd1 vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__a21o_1
X_08097_ top.cb_syn.char_path_n\[121\] net383 net342 top.cb_syn.char_path_n\[119\]
+ net187 vssd1 vssd1 vccd1 vccd1 _04576_ sky130_fd_sc_hd__a221o_1
Xclkload90 clknet_leaf_83_clk vssd1 vssd1 vccd1 vccd1 clkload90/X sky130_fd_sc_hd__clkbuf_8
X_07048_ net496 top.findLeastValue.val2\[25\] _03705_ vssd1 vssd1 vccd1 vccd1 _03706_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout876_A net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout497_X net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout664_X net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08999_ top.WB.CPU_DAT_O\[26\] net1137 net318 vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__mux2_1
XANTENNA__09323__B1 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10961_ clknet_leaf_58_clk net920 _00316_ vssd1 vssd1 vccd1 vccd1 top.controller.fin_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10892_ clknet_leaf_110_clk _01469_ _00247_ vssd1 vssd1 vccd1 vccd1 top.translation.resEn
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_26_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08834__C1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11513_ clknet_leaf_70_clk _02061_ _00868_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least1\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_11444_ clknet_leaf_67_clk _01992_ _00799_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.histo_index\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__05663__A2 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08362__A top.cb_syn.end_cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11375_ clknet_leaf_104_clk _01923_ _00730_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_98_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10326_ net766 net606 vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__and2_1
X_10257_ net858 net698 vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__and2_1
XFILLER_105_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10188_ net862 net702 vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__and2_1
XFILLER_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07628__A0 top.findLeastValue.least1\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_06350_ top.hist_data_o\[24\] _03196_ _03191_ vssd1 vssd1 vccd1 vccd1 _03206_ sky130_fd_sc_hd__o21ba_1
XANTENNA__08825__C1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06281_ top.cb_syn.curr_index\[2\] _02558_ _03143_ net463 _03146_ vssd1 vssd1 vccd1
+ vccd1 _03147_ sky130_fd_sc_hd__a221o_1
X_05301_ top.compVal\[41\] vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__inv_2
X_08020_ _04519_ _04521_ vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__and2_1
XANTENNA__05654__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold703 top.translation.index\[6\] vssd1 vssd1 vccd1 vccd1 net1656 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_77_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold714 top.histogram.sram_out\[3\] vssd1 vssd1 vccd1 vccd1 net1667 sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 top.compVal\[6\] vssd1 vssd1 vccd1 vccd1 net1689 sky130_fd_sc_hd__dlygate4sd3_1
Xhold725 top.findLeastValue.sum\[8\] vssd1 vssd1 vccd1 vccd1 net1678 sky130_fd_sc_hd__dlygate4sd3_1
X_09971_ net783 net623 vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__and2_1
XFILLER_89_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold758 top.findLeastValue.sum\[34\] vssd1 vssd1 vccd1 vccd1 net1711 sky130_fd_sc_hd__dlygate4sd3_1
Xhold769 top.histogram.total\[6\] vssd1 vssd1 vccd1 vccd1 net1722 sky130_fd_sc_hd__dlygate4sd3_1
Xhold747 top.compVal\[40\] vssd1 vssd1 vccd1 vccd1 net1700 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08922_ net456 net546 vssd1 vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__nand2_1
XANTENNA__10026__B net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08356__B2 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout192_A net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08853_ _04925_ _05033_ net325 _02786_ net473 vssd1 vssd1 vccd1 vccd1 _05036_ sky130_fd_sc_hd__a2111o_1
X_05996_ net1717 _02904_ vssd1 vssd1 vccd1 vccd1 _02923_ sky130_fd_sc_hd__nor2_1
X_07804_ top.findLeastValue.sum\[27\] top.hTree.tree_reg\[27\] net285 vssd1 vssd1
+ vccd1 vccd1 _04349_ sky130_fd_sc_hd__mux2_1
X_08784_ top.path\[116\] net409 net327 top.path\[117\] _02522_ vssd1 vssd1 vccd1 vccd1
+ _04967_ sky130_fd_sc_hd__o221a_1
X_07735_ top.hTree.tree_reg\[41\] top.findLeastValue.sum\[41\] net250 vssd1 vssd1
+ vccd1 vccd1 _04294_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout457_A net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09117__C_N _05087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09405_ net979 net241 _05279_ _05280_ vssd1 vssd1 vccd1 vccd1 _01449_ sky130_fd_sc_hd__a22o_1
X_07666_ net267 _04237_ _04238_ net1163 net445 vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__a32o_1
XFILLER_53_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07597_ net1451 _04182_ _04144_ vssd1 vssd1 vccd1 vccd1 _01873_ sky130_fd_sc_hd__mux2_1
XFILLER_13_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_06617_ top.compVal\[32\] _02469_ _03392_ vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07619__B1 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06548_ _03330_ _03336_ vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__nor2_1
X_09336_ net1028 net236 net214 _04442_ vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__a22o_1
X_09267_ top.cb_syn.zero_count\[0\] top.cb_syn.zero_count\[1\] top.cb_syn.zero_count\[2\]
+ top.cb_syn.zero_count\[3\] vssd1 vssd1 vccd1 vccd1 _05221_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_23_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08218_ top.cb_syn.char_path_n\[60\] net208 _04636_ vssd1 vssd1 vccd1 vccd1 _01706_
+ sky130_fd_sc_hd__o21a_1
X_06479_ _03291_ _03297_ vssd1 vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__nor2_1
X_09198_ top.hTree.state\[4\] net264 _05162_ net1535 vssd1 vssd1 vccd1 vccd1 _00023_
+ sky130_fd_sc_hd__a22o_1
X_08149_ top.cb_syn.char_path_n\[95\] net388 net346 top.cb_syn.char_path_n\[93\] net192
+ vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__a221o_1
X_11160_ clknet_leaf_18_clk _01708_ _00515_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout879_X net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11091_ clknet_leaf_25_clk _01639_ _00446_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[121\]
+ sky130_fd_sc_hd__dfrtp_1
X_10111_ net813 net653 vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__and2_1
X_10042_ net820 net660 vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__and2_1
Xhold30 top.hTree.node_reg\[7\] vssd1 vssd1 vccd1 vccd1 net983 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 top.hTree.node_reg\[8\] vssd1 vssd1 vccd1 vccd1 net994 sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 top.sram_interface.init_counter\[23\] vssd1 vssd1 vccd1 vccd1 net1016 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 top.sram_interface.init_counter\[16\] vssd1 vssd1 vccd1 vccd1 net1027 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 top.hTree.node_reg\[48\] vssd1 vssd1 vccd1 vccd1 net1005 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 net110 vssd1 vssd1 vccd1 vccd1 net1038 sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 net48 vssd1 vssd1 vccd1 vccd1 net1049 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input18_A DAT_I[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10944_ clknet_leaf_33_clk _01499_ _00299_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.num_lefts\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07858__B1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10875_ clknet_leaf_41_clk _00006_ _00230_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.curr_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_42_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09075__A2 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08807__C1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06308__C net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05636__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_5 top.findLeastValue.histo_index\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11427_ clknet_leaf_85_clk _01975_ _00782_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[33\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_113_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11358_ clknet_leaf_97_clk _01906_ _00713_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[10\]
+ sky130_fd_sc_hd__dfrtp_2
X_10309_ net812 net652 vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__and2_1
X_11289_ clknet_leaf_84_clk _01837_ _00644_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05850_ top.compVal\[17\] net168 net154 top.WB.CPU_DAT_O\[17\] vssd1 vssd1 vccd1
+ vccd1 _02292_ sky130_fd_sc_hd__a22o_1
X_07520_ top.cb_syn.char_path_n\[124\] top.cb_syn.char_path_n\[123\] top.cb_syn.char_path_n\[122\]
+ top.cb_syn.char_path_n\[121\] net401 net352 vssd1 vssd1 vccd1 vccd1 _04111_ sky130_fd_sc_hd__mux4_1
X_05781_ _02796_ _02800_ vssd1 vssd1 vccd1 vccd1 _02801_ sky130_fd_sc_hd__nor2_2
XFILLER_35_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07451_ net1649 top.dut.out_valid_next _04002_ _04028_ _04043_ vssd1 vssd1 vccd1
+ vccd1 _01880_ sky130_fd_sc_hd__o221a_1
X_07382_ _03984_ _03985_ vssd1 vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__and2_1
X_06402_ net1467 net299 _03237_ _03238_ vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__a22o_1
X_09121_ net548 net468 net414 top.sram_interface.word_cnt\[14\] net461 vssd1 vssd1
+ vccd1 vccd1 _05137_ sky130_fd_sc_hd__a32o_1
X_06333_ net1157 _03195_ net303 vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_123_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_123_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_20_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06264_ net1429 net145 _03130_ net160 vssd1 vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__a22o_1
XANTENNA__06074__X _02949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09052_ net1390 top.WB.CPU_DAT_O\[5\] net293 vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__mux2_1
X_08003_ _02499_ top.cb_syn.zeroes\[7\] top.cb_syn.zeroes\[6\] _02500_ _04505_ vssd1
+ vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__a221o_1
X_06195_ net501 _03012_ net498 vssd1 vssd1 vccd1 vccd1 _03064_ sky130_fd_sc_hd__a21oi_1
Xhold500 top.hTree.tree_reg\[62\] vssd1 vssd1 vccd1 vccd1 net1453 sky130_fd_sc_hd__dlygate4sd3_1
Xhold511 top.hist_data_o\[16\] vssd1 vssd1 vccd1 vccd1 net1464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold533 top.dut.out\[4\] vssd1 vssd1 vccd1 vccd1 net1486 sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 top.cb_syn.curr_index\[1\] vssd1 vssd1 vccd1 vccd1 net1475 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout205_A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold544 top.hTree.nullSumIndex\[3\] vssd1 vssd1 vccd1 vccd1 net1497 sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 top.header_synthesis.count\[7\] vssd1 vssd1 vccd1 vccd1 net1519 sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 top.hist_addr\[5\] vssd1 vssd1 vccd1 vccd1 net1530 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold588 top.hTree.tree_reg\[32\] vssd1 vssd1 vccd1 vccd1 net1541 sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 top.hist_data_o\[3\] vssd1 vssd1 vccd1 vccd1 net1508 sky130_fd_sc_hd__dlygate4sd3_1
X_09954_ net769 net609 vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__and2_1
Xhold599 top.histogram.total\[29\] vssd1 vssd1 vccd1 vccd1 net1552 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08905_ top.cb_syn.max_index\[5\] _05065_ top.cb_syn.max_index\[6\] vssd1 vssd1 vccd1
+ vccd1 _05074_ sky130_fd_sc_hd__a21oi_1
X_09885_ net739 net579 vssd1 vssd1 vccd1 vccd1 _00499_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout574_A net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08836_ _05015_ _05018_ vssd1 vssd1 vccd1 vccd1 _05019_ sky130_fd_sc_hd__nor2_1
XANTENNA__07780__S net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05979_ top.sram_interface.init_counter\[8\] top.sram_interface.init_counter\[7\]
+ _02914_ vssd1 vssd1 vccd1 vccd1 _02915_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout362_X net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06760__B1 _03547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08767_ top.path\[82\] top.path\[83\] net526 vssd1 vssd1 vccd1 vccd1 _04950_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout741_A net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08698_ _04876_ _04885_ _04892_ _04875_ net1668 vssd1 vssd1 vccd1 vccd1 _01482_ sky130_fd_sc_hd__a32o_1
X_07718_ net444 net1525 net255 top.findLeastValue.sum\[45\] _04280_ vssd1 vssd1 vccd1
+ vccd1 _01850_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_0_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07649_ top.hTree.tree_reg\[57\] net394 net285 vssd1 vssd1 vccd1 vccd1 _04224_ sky130_fd_sc_hd__and3_1
XFILLER_53_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10660_ clknet_leaf_118_clk _01259_ _00079_ vssd1 vssd1 vccd1 vccd1 top.path\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_09319_ net436 _05250_ _05252_ _05253_ vssd1 vssd1 vccd1 vccd1 _05254_ sky130_fd_sc_hd__a22o_1
X_10591_ net747 net587 vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_114_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_114_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__05967__C _02760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05618__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06144__B net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11212_ clknet_leaf_23_clk _01760_ _00567_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[114\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput53 net53 vssd1 vssd1 vccd1 vccd1 ADR_O[18] sky130_fd_sc_hd__buf_2
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 ADR_O[2] sky130_fd_sc_hd__buf_2
X_11143_ clknet_leaf_6_clk _01691_ _00498_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[45\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_8_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 DAT_O[11] sky130_fd_sc_hd__buf_2
Xoutput97 net97 vssd1 vssd1 vccd1 vccd1 DAT_O[31] sky130_fd_sc_hd__buf_2
Xoutput86 net86 vssd1 vssd1 vccd1 vccd1 DAT_O[21] sky130_fd_sc_hd__buf_2
X_11074_ clknet_leaf_10_clk _01622_ _00429_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[104\]
+ sky130_fd_sc_hd__dfrtp_1
X_10025_ net822 net662 vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__and2_1
XANTENNA__07543__X _04134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10927_ clknet_leaf_30_clk _01482_ _00282_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.zeroes\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_55_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10858_ clknet_leaf_78_clk _01444_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[50\]
+ sky130_fd_sc_hd__dfxtp_1
X_10789_ clknet_leaf_52_clk _00029_ _00208_ vssd1 vssd1 vccd1 vccd1 top.histogram.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_105_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_105_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_117_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09205__C1 top.CB_write_complete vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06054__B net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07767__C1 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout309 _02762_ vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__buf_2
X_06951_ top.findLeastValue.val2\[8\] net149 net122 _03617_ vssd1 vssd1 vccd1 vccd1
+ _01950_ sky130_fd_sc_hd__o22a_1
X_09670_ net781 net621 vssd1 vssd1 vccd1 vccd1 _00284_ sky130_fd_sc_hd__and2_1
X_05902_ _02857_ _02875_ vssd1 vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__nand2_1
X_08621_ _04836_ _04838_ vssd1 vssd1 vccd1 vccd1 _01505_ sky130_fd_sc_hd__and2_1
X_06882_ top.compVal\[42\] top.findLeastValue.val1\[42\] net165 vssd1 vssd1 vccd1
+ vccd1 _03583_ sky130_fd_sc_hd__mux2_1
X_05833_ net556 _02843_ vssd1 vssd1 vccd1 vccd1 _02844_ sky130_fd_sc_hd__nor2_1
XFILLER_27_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08552_ net1232 top.cb_syn.char_path_n\[24\] net229 vssd1 vssd1 vccd1 vccd1 _01542_
+ sky130_fd_sc_hd__mux2_1
X_05764_ net473 _02784_ vssd1 vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__or2_1
X_08483_ net1155 top.cb_syn.char_path_n\[93\] net234 vssd1 vssd1 vccd1 vccd1 _01611_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_85_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07503_ top.cb_syn.char_path_n\[48\] top.cb_syn.char_path_n\[47\] top.cb_syn.char_path_n\[46\]
+ top.cb_syn.char_path_n\[45\] net400 net351 vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__mux4_1
X_07434_ top.dut.bit_buf\[3\] net41 net721 vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__mux2_1
XANTENNA__05848__A2 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05695_ net19 net415 net308 top.WB.CPU_DAT_O\[25\] vssd1 vssd1 vccd1 vccd1 _02363_
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout155_A net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06944__S net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07365_ top.cw1\[5\] net167 vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_4_8_0_clk_X clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout322_A net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09104_ top.sram_interface.word_cnt\[1\] _05116_ _02818_ vssd1 vssd1 vccd1 vccd1
+ _05124_ sky130_fd_sc_hd__a21bo_1
X_07296_ top.findLeastValue.val1\[20\] top.findLeastValue.val2\[20\] _03923_ vssd1
+ vssd1 vccd1 vccd1 _03930_ sky130_fd_sc_hd__a21oi_1
X_06316_ top.hist_data_o\[8\] _03178_ vssd1 vssd1 vccd1 vccd1 _03179_ sky130_fd_sc_hd__and2_1
X_06247_ _03001_ _03113_ vssd1 vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__nand2_1
X_09035_ net1059 top.WB.CPU_DAT_O\[22\] net291 vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout208_X net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06178_ top.sram_interface.init_counter\[6\] _02945_ vssd1 vssd1 vccd1 vccd1 _03048_
+ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout691_A net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold341 top.cb_syn.char_path\[85\] vssd1 vssd1 vccd1 vccd1 net1294 sky130_fd_sc_hd__dlygate4sd3_1
Xhold352 top.path\[43\] vssd1 vssd1 vccd1 vccd1 net1305 sky130_fd_sc_hd__dlygate4sd3_1
Xhold330 net100 vssd1 vssd1 vccd1 vccd1 net1283 sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 top.hTree.nulls\[58\] vssd1 vssd1 vccd1 vccd1 net1327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 top.path\[61\] vssd1 vssd1 vccd1 vccd1 net1338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold363 top.cb_syn.char_path\[75\] vssd1 vssd1 vccd1 vccd1 net1316 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 top.cb_syn.char_path\[8\] vssd1 vssd1 vccd1 vccd1 net1349 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout843 net878 vssd1 vssd1 vccd1 vccd1 net843 sky130_fd_sc_hd__clkbuf_2
X_09937_ net791 net631 vssd1 vssd1 vccd1 vccd1 _00551_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_5_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout810 net811 vssd1 vssd1 vccd1 vccd1 net810 sky130_fd_sc_hd__clkbuf_2
Xfanout832 net834 vssd1 vssd1 vccd1 vccd1 net832 sky130_fd_sc_hd__clkbuf_2
Xfanout821 net823 vssd1 vssd1 vccd1 vccd1 net821 sky130_fd_sc_hd__buf_1
Xfanout876 net877 vssd1 vssd1 vccd1 vccd1 net876 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout854 net855 vssd1 vssd1 vccd1 vccd1 net854 sky130_fd_sc_hd__clkbuf_2
Xfanout865 net866 vssd1 vssd1 vccd1 vccd1 net865 sky130_fd_sc_hd__clkbuf_2
X_09868_ net778 net618 vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__and2_1
X_09799_ net775 net615 vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__and2_1
XFILLER_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout744_X net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05536__A1 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08819_ top.path\[4\] net410 net328 top.path\[5\] net522 vssd1 vssd1 vccd1 vccd1
+ _05002_ sky130_fd_sc_hd__o221a_1
XFILLER_18_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11830_ clknet_leaf_100_clk _02346_ _01185_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_26_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11761_ clknet_leaf_114_clk _02294_ _01116_ vssd1 vssd1 vccd1 vccd1 top.compVal\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05839__A2 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10712_ clknet_leaf_3_clk _01311_ _00131_ vssd1 vssd1 vccd1 vccd1 top.path\[88\]
+ sky130_fd_sc_hd__dfrtp_1
X_11692_ clknet_leaf_62_clk _02225_ _01047_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10643_ clknet_leaf_49_clk _00052_ _00062_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.word_cnt\[9\]
+ sky130_fd_sc_hd__dfrtp_2
X_10574_ net814 net654 vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__and2_1
XANTENNA__08789__A1 top.translation.index\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06264__A2 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_5_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11126_ clknet_leaf_29_clk _01674_ _00481_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[28\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_96_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11057_ clknet_leaf_20_clk _01605_ _00412_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[87\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_37_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10008_ net818 net658 vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__and2_1
XFILLER_91_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_17_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06049__B net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05480_ top.WB.curr_state\[0\] net212 vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_50_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07150_ _03798_ _03806_ _03807_ vssd1 vssd1 vccd1 vccd1 _03808_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_30_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06101_ top.TRN_char_index\[1\] top.TRN_char_index\[0\] top.TRN_char_index\[2\] vssd1
+ vssd1 vccd1 vccd1 _02974_ sky130_fd_sc_hd__o21a_1
XFILLER_9_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07081_ top.findLeastValue.val1\[6\] top.findLeastValue.val2\[6\] vssd1 vssd1 vccd1
+ vccd1 _03739_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_10_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06032_ net1508 top.WB.CPU_DAT_O\[3\] net355 vssd1 vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__mux2_1
XANTENNA__06004__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout117 _03552_ vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__clkbuf_4
Xfanout128 net129 vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__clkbuf_4
Xfanout139 net140 vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__buf_4
X_07983_ _02515_ top.cb_syn.zero_count\[1\] top.cb_syn.zeroes\[0\] _02531_ vssd1 vssd1
+ vccd1 vccd1 _04486_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__06963__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09722_ net735 net575 vssd1 vssd1 vccd1 vccd1 _00336_ sky130_fd_sc_hd__and2_1
XANTENNA__08165__C1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06934_ top.compVal\[16\] top.findLeastValue.val1\[16\] net161 vssd1 vssd1 vccd1
+ vccd1 _03609_ sky130_fd_sc_hd__mux2_1
X_09653_ net784 net624 vssd1 vssd1 vccd1 vccd1 _00267_ sky130_fd_sc_hd__and2_1
XFILLER_95_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06865_ net497 _03571_ _03568_ vssd1 vssd1 vccd1 vccd1 _03577_ sky130_fd_sc_hd__a21bo_1
XANTENNA_fanout272_A _03864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_08604_ net1263 _04823_ _04536_ vssd1 vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__a21o_1
X_05816_ _02828_ _02830_ _02833_ vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__and3b_1
X_09584_ net845 net685 vssd1 vssd1 vccd1 vccd1 _00198_ sky130_fd_sc_hd__and2_1
XANTENNA__05415__Y _02523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_118_Right_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_06796_ top.findLeastValue.val1\[34\] net133 net117 top.compVal\[34\] vssd1 vssd1
+ vccd1 vccd1 _02042_ sky130_fd_sc_hd__o22a_1
X_08535_ net1091 top.cb_syn.char_path_n\[41\] net225 vssd1 vssd1 vccd1 vccd1 _01559_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout537_A top.cb_syn.curr_state\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05747_ net452 top.sram_interface.word_cnt\[5\] _02781_ _02529_ _02780_ vssd1 vssd1
+ vccd1 vccd1 _02782_ sky130_fd_sc_hd__a221o_2
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05678_ top.cb_syn.char_path\[64\] net554 net545 top.cb_syn.char_path\[32\] vssd1
+ vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__a22o_1
XFILLER_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08466_ net1203 top.cb_syn.char_path_n\[110\] net220 vssd1 vssd1 vccd1 vccd1 _01628_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09050__S net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07417_ _03992_ _04015_ net404 vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__mux2_1
XANTENNA__07691__B2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08397_ _02506_ top.cb_syn.char_path_n\[12\] _04755_ net509 vssd1 vssd1 vccd1 vccd1
+ _04756_ sky130_fd_sc_hd__o211a_1
X_07348_ top.findLeastValue.sum\[6\] net274 _03966_ vssd1 vssd1 vccd1 vccd1 _01902_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_98_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07279_ _03683_ _03916_ vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__nand2_1
XFILLER_117_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10290_ net724 net564 vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__and2_1
X_09018_ top.WB.CPU_DAT_O\[7\] net1345 net320 vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__mux2_1
Xteam_05_912 vssd1 vssd1 vccd1 vccd1 team_05_912/HI gpio_out[27] sky130_fd_sc_hd__conb_1
Xhold171 top.header_synthesis.header\[5\] vssd1 vssd1 vccd1 vccd1 net1124 sky130_fd_sc_hd__dlygate4sd3_1
Xteam_05_901 vssd1 vssd1 vccd1 vccd1 team_05_901/HI gpio_out[16] sky130_fd_sc_hd__conb_1
Xhold160 top.cb_syn.char_path\[10\] vssd1 vssd1 vccd1 vccd1 net1113 sky130_fd_sc_hd__dlygate4sd3_1
Xteam_05_923 vssd1 vssd1 vccd1 vccd1 gpio_oeb[3] team_05_923/LO sky130_fd_sc_hd__conb_1
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold182 top.cb_syn.char_path\[90\] vssd1 vssd1 vccd1 vccd1 net1135 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 top.cb_syn.char_path\[17\] vssd1 vssd1 vccd1 vccd1 net1146 sky130_fd_sc_hd__dlygate4sd3_1
Xteam_05_945 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] team_05_945/LO sky130_fd_sc_hd__conb_1
Xteam_05_934 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] team_05_934/LO sky130_fd_sc_hd__conb_1
Xfanout640 net646 vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout651 net664 vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__buf_1
XANTENNA__05757__B2 top.WB.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout684 net685 vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06849__S _03424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout662 net663 vssd1 vssd1 vccd1 vccd1 net662 sky130_fd_sc_hd__clkbuf_2
XANTENNA_hold749_A top.findLeastValue.sum\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout673 net674 vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__buf_1
Xfanout695 net696 vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__clkbuf_2
XFILLER_58_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08171__A2 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11813_ clknet_leaf_97_clk _02330_ _01168_ vssd1 vssd1 vccd1 vccd1 top.compVal\[45\]
+ sky130_fd_sc_hd__dfrtp_2
X_11744_ clknet_leaf_94_clk _02277_ _01099_ vssd1 vssd1 vccd1 vccd1 top.compVal\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_11675_ clknet_leaf_60_clk _02208_ _01030_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10626_ net805 net645 vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__and2_1
X_10557_ net870 net710 vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__and2_1
XANTENNA__08631__B1 _04826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09196__A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10488_ net830 net670 vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__and2_1
XANTENNA__07737__A2 _04294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06945__B1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11109_ clknet_leaf_3_clk _01657_ _00464_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08698__B1 _04875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08162__A2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06650_ _03427_ _03429_ _03432_ _03434_ vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_69_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08974__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05601_ _02687_ _02688_ vssd1 vssd1 vccd1 vccd1 _02689_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_82_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06581_ _02434_ top.findLeastValue.val1\[15\] top.findLeastValue.val1\[14\] _02435_
+ vssd1 vssd1 vccd1 vccd1 _03370_ sky130_fd_sc_hd__o22a_1
X_05532_ net1122 net144 _02631_ net177 vssd1 vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__a22o_1
X_08320_ top.cb_syn.char_path_n\[9\] net199 _04687_ vssd1 vssd1 vccd1 vccd1 _01655_
+ sky130_fd_sc_hd__o21a_1
X_05463_ net460 net541 _02566_ _02569_ _02570_ vssd1 vssd1 vccd1 vccd1 _02571_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10955__D top.controller.fin_TRN vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08251_ top.cb_syn.char_path_n\[44\] net373 net333 top.cb_syn.char_path_n\[42\] net178
+ vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__a221o_1
X_07202_ _03855_ _03857_ _03859_ vssd1 vssd1 vccd1 vccd1 _03860_ sky130_fd_sc_hd__a21o_1
X_05394_ top.cb_syn.count\[3\] vssd1 vssd1 vccd1 vccd1 _02502_ sky130_fd_sc_hd__inv_2
X_08182_ top.cb_syn.char_path_n\[78\] net196 _04618_ vssd1 vssd1 vccd1 vccd1 _01724_
+ sky130_fd_sc_hd__o21a_1
X_07133_ top.findLeastValue.val1\[19\] top.findLeastValue.val2\[19\] vssd1 vssd1 vccd1
+ vccd1 _03791_ sky130_fd_sc_hd__nand2_1
XANTENNA__07520__S1 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07064_ _03715_ _03718_ _03721_ vssd1 vssd1 vccd1 vccd1 _03722_ sky130_fd_sc_hd__and3_1
X_06015_ net1477 top.WB.CPU_DAT_O\[20\] net357 vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_93_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout487_A net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07966_ _02763_ _04473_ _02765_ vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__a21oi_1
XFILLER_75_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09705_ net850 net690 vssd1 vssd1 vccd1 vccd1 _00319_ sky130_fd_sc_hd__and2_1
XANTENNA__09045__S net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06917_ top.findLeastValue.val2\[25\] net148 net124 _03600_ vssd1 vssd1 vccd1 vccd1
+ _01967_ sky130_fd_sc_hd__o22a_1
X_09636_ net801 net641 vssd1 vssd1 vccd1 vccd1 _00250_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_94_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_94_clk sky130_fd_sc_hd__clkbuf_8
X_07897_ net425 _04422_ _04423_ net258 vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__o211a_1
X_06848_ _02479_ net152 net126 _03563_ vssd1 vssd1 vccd1 vccd1 _01999_ sky130_fd_sc_hd__a2bb2o_1
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09567_ net843 net683 vssd1 vssd1 vccd1 vccd1 _00181_ sky130_fd_sc_hd__and2_1
X_06779_ top.findLeastValue.least1\[1\] net136 net118 net503 vssd1 vssd1 vccd1 vccd1
+ _02057_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout442_X net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout821_A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08518_ net1249 top.cb_syn.char_path_n\[58\] net232 vssd1 vssd1 vccd1 vccd1 _01576_
+ sky130_fd_sc_hd__mux2_1
X_09498_ net749 net589 vssd1 vssd1 vccd1 vccd1 _00112_ sky130_fd_sc_hd__and2_1
XANTENNA__08616__C net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08449_ net1518 top.cb_syn.char_path_n\[127\] net232 vssd1 vssd1 vccd1 vccd1 _01645_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_102_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11460_ clknet_leaf_93_clk _02008_ _00815_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__06219__A2 _02595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10411_ net795 net635 vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11391_ clknet_leaf_82_clk _01939_ _00746_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[43\]
+ sky130_fd_sc_hd__dfrtp_1
X_10342_ net871 net711 vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__and2_1
XANTENNA__07511__S1 _04071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09169__A1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10273_ net727 net567 vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__and2_1
Xfanout470 top.controller.state_reg\[2\] vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__clkbuf_4
Xfanout481 top.controller.state_reg\[1\] vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__clkbuf_2
Xfanout492 net493 vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__clkbuf_2
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_85_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_19_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08794__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_14_Left_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11727_ clknet_leaf_121_clk _02260_ _01082_ vssd1 vssd1 vccd1 vccd1 top.path\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11658_ clknet_leaf_108_clk _02191_ _01013_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11589_ clknet_leaf_45_clk _02137_ _00944_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10609_ net752 net592 vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_40_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07502__S1 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_23_Left_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07820_ top.findLeastValue.sum\[24\] _04361_ net395 vssd1 vssd1 vccd1 vccd1 _04362_
+ sky130_fd_sc_hd__mux2_1
XFILLER_96_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07751_ net488 _04305_ vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__or2_1
XFILLER_84_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_76_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_clk sky130_fd_sc_hd__clkbuf_8
X_06702_ _03489_ _03487_ _03488_ vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__or3b_1
XANTENNA_clkbuf_leaf_92_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07682_ _02475_ net396 _04250_ vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__o21a_1
XANTENNA__08766__S0 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09421_ top.hTree.nulls\[61\] _04207_ net406 vssd1 vssd1 vccd1 vccd1 _05291_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_32_Left_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06633_ _03403_ _03421_ _03391_ vssd1 vssd1 vccd1 vccd1 _03422_ sky130_fd_sc_hd__a21boi_2
XANTENNA__07621__B net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09352_ net1424 net240 net217 _04378_ vssd1 vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__a22o_1
X_06564_ _02438_ top.findLeastValue.val1\[11\] top.findLeastValue.val1\[10\] _02439_
+ vssd1 vssd1 vccd1 vccd1 _03353_ sky130_fd_sc_hd__o22a_1
X_05515_ top.cb_syn.char_path\[91\] net553 net544 top.cb_syn.char_path\[59\] vssd1
+ vssd1 vccd1 vccd1 _02617_ sky130_fd_sc_hd__a22o_1
XFILLER_80_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08303_ top.cb_syn.char_path_n\[18\] net375 net335 top.cb_syn.char_path_n\[16\] net180
+ vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__a221o_1
XANTENNA__05422__A net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09283_ top.dut.bits_in_buf_next\[1\] _04000_ _04037_ vssd1 vssd1 vccd1 vccd1 top.dut.bit_buf_next\[1\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout235_A _04805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06495_ net1490 _03284_ vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__xor2_1
XANTENNA__08733__A top.header_synthesis.enable vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_30_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05446_ top.CB_write_complete top.CB_read_complete vssd1 vssd1 vccd1 vccd1 _02554_
+ sky130_fd_sc_hd__or2_1
X_08234_ top.cb_syn.char_path_n\[52\] net197 _04644_ vssd1 vssd1 vccd1 vccd1 _01698_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__06952__S net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08165_ top.cb_syn.char_path_n\[87\] net387 net346 top.cb_syn.char_path_n\[85\] net191
+ vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__a221o_1
X_05377_ top.findLeastValue.val2\[37\] vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__inv_2
XFILLER_109_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07116_ _03773_ vssd1 vssd1 vccd1 vccd1 _03774_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_41_Left_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08096_ top.cb_syn.char_path_n\[121\] net206 _04575_ vssd1 vssd1 vccd1 vccd1 _01767_
+ sky130_fd_sc_hd__o21a_1
Xclkload80 clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 clkload80/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_45_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload91 clknet_leaf_85_clk vssd1 vssd1 vccd1 vccd1 clkload91/Y sky130_fd_sc_hd__clkinv_2
X_07047_ net496 top.findLeastValue.val2\[25\] top.findLeastValue.val2\[24\] top.findLeastValue.val1\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout771_A net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout392_X net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__09020__A0 top.WB.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06909__B1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08998_ top.WB.CPU_DAT_O\[27\] net1297 net317 vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_67_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_clk sky130_fd_sc_hd__clkbuf_8
X_07949_ net1500 _04464_ _04461_ vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_50_Left_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08126__A2 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10960_ clknet_leaf_59_clk net957 _00315_ vssd1 vssd1 vccd1 vccd1 top.controller.fin_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_103_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08757__S0 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09619_ net798 net638 vssd1 vssd1 vccd1 vccd1 _00233_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout824_X net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07885__A1 top.findLeastValue.sum\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10891_ clknet_leaf_110_clk _01468_ _00246_ vssd1 vssd1 vccd1 vccd1 top.translation.index\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_clkbuf_leaf_118_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11512_ clknet_leaf_70_clk _02060_ _00867_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least1\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__05648__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_11443_ clknet_leaf_68_clk _01991_ _00798_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.histo_index\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_109_142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07496__S0 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11374_ clknet_leaf_79_clk _01922_ _00729_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_115_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10325_ net766 net606 vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__and2_1
XANTENNA__05820__B1 _02581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10256_ net862 net702 vssd1 vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__and2_1
XANTENNA__09011__A0 top.WB.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10187_ net862 net702 vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_58_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09314__B2 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_11_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_11_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_66_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06280_ _03127_ _03145_ _03144_ net460 vssd1 vssd1 vccd1 vccd1 _03146_ sky130_fd_sc_hd__a2bb2o_1
X_05300_ top.compVal\[43\] vssd1 vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__inv_2
Xhold715 top.cb_syn.zeroes\[1\] vssd1 vssd1 vccd1 vccd1 net1668 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06064__B1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold704 top.cw2\[5\] vssd1 vssd1 vccd1 vccd1 net1657 sky130_fd_sc_hd__dlygate4sd3_1
Xhold737 top.histogram.state\[2\] vssd1 vssd1 vccd1 vccd1 net1690 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07487__S0 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold726 top.hTree.state\[8\] vssd1 vssd1 vccd1 vccd1 net1679 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold748 top.cb_syn.i\[5\] vssd1 vssd1 vccd1 vccd1 net1701 sky130_fd_sc_hd__dlygate4sd3_1
X_09970_ net783 net623 vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__and2_1
Xhold759 top.compVal\[2\] vssd1 vssd1 vccd1 vccd1 net1712 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08921_ _02525_ _05072_ vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09002__A0 top.WB.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08852_ top.TRN_char_index\[5\] top.TRN_char_index\[2\] _03123_ _05034_ vssd1 vssd1
+ vccd1 vccd1 _05035_ sky130_fd_sc_hd__nor4_2
XFILLER_97_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08356__A2 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07803_ net443 net1575 net254 top.findLeastValue.sum\[28\] _04348_ vssd1 vssd1 vccd1
+ vccd1 _01833_ sky130_fd_sc_hd__a221o_1
X_05995_ _02913_ _02922_ vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_49_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout185_A net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08783_ top.path\[118\] top.path\[119\] net526 vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__mux2_1
XFILLER_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05778__D_N top.findLeastValue.least2\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07734_ top.findLeastValue.sum\[41\] top.hTree.tree_reg\[41\] _04197_ vssd1 vssd1
+ vccd1 vccd1 _04293_ sky130_fd_sc_hd__mux2_1
X_07665_ net485 _04235_ vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__or2_1
XFILLER_53_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout352_A net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09404_ top.hTree.nulls\[55\] net407 net244 vssd1 vssd1 vccd1 vccd1 _05280_ sky130_fd_sc_hd__o21a_1
XFILLER_25_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06616_ _02411_ top.findLeastValue.val1\[38\] top.findLeastValue.val1\[34\] _02414_
+ _03390_ vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__a221o_1
X_07596_ top.cb_syn.max_index\[2\] _04136_ _04178_ _04181_ vssd1 vssd1 vccd1 vccd1
+ _04182_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout140_X net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09335_ net999 net239 net219 _04446_ vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__a22o_1
X_06547_ top.compVal\[28\] _02470_ _03331_ _03335_ vssd1 vssd1 vccd1 vccd1 _03336_
+ sky130_fd_sc_hd__o22a_1
X_09266_ _05219_ vssd1 vssd1 vccd1 vccd1 _05220_ sky130_fd_sc_hd__inv_2
XANTENNA__06535__X _03325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06478_ net1721 _03290_ net1469 vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_23_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05429_ net471 vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__inv_2
X_08217_ top.cb_syn.char_path_n\[61\] net387 net348 top.cb_syn.char_path_n\[59\] net193
+ vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__a221o_1
XFILLER_119_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09197_ net962 net265 _05179_ net491 vssd1 vssd1 vccd1 vccd1 _00017_ sky130_fd_sc_hd__a22o_1
XFILLER_107_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08148_ top.cb_syn.char_path_n\[95\] net208 _04601_ vssd1 vssd1 vccd1 vccd1 _01741_
+ sky130_fd_sc_hd__o21a_1
X_08079_ _04133_ _04563_ _04555_ _02931_ _04562_ vssd1 vssd1 vccd1 vccd1 _04566_ sky130_fd_sc_hd__a2111o_1
X_11090_ clknet_leaf_24_clk _01638_ _00445_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[120\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08402__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10110_ net813 net653 vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__and2_1
XFILLER_88_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10041_ net820 net660 vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__and2_1
Xhold20 top.sram_interface.init_counter\[12\] vssd1 vssd1 vccd1 vccd1 net973 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 top.hTree.node_reg\[34\] vssd1 vssd1 vccd1 vccd1 net984 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 top.sram_interface.init_counter\[17\] vssd1 vssd1 vccd1 vccd1 net1017 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_110_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold53 top.hTree.node_reg\[33\] vssd1 vssd1 vccd1 vccd1 net1006 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 top.hTree.node_reg\[9\] vssd1 vssd1 vccd1 vccd1 net995 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_90_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold97 top.hTree.node_reg\[14\] vssd1 vssd1 vccd1 vccd1 net1050 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold731_A top.findLeastValue.sum\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xhold75 top.hTree.node_reg\[4\] vssd1 vssd1 vccd1 vccd1 net1028 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 top.hTree.node_reg\[44\] vssd1 vssd1 vccd1 vccd1 net1039 sky130_fd_sc_hd__dlygate4sd3_1
X_10943_ clknet_leaf_36_clk _01498_ _00298_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.cb_length\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07542__A net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05581__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07858__A1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07307__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05614__X _02700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07858__B2 top.findLeastValue.sum\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10874_ clknet_leaf_36_clk _00005_ _00229_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.curr_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06833__A2 net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_11426_ clknet_leaf_86_clk _01974_ _00781_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[32\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA_6 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11357_ clknet_leaf_97_clk _01905_ _00712_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[9\]
+ sky130_fd_sc_hd__dfrtp_2
X_10308_ net824 net664 vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__and2_1
X_11288_ clknet_leaf_84_clk net1409 _00643_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_72_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10239_ net833 net673 vssd1 vssd1 vccd1 vccd1 _00853_ sky130_fd_sc_hd__and2_1
XFILLER_79_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05780_ top.findLeastValue.least2\[8\] _02799_ vssd1 vssd1 vccd1 vccd1 _02800_ sky130_fd_sc_hd__nand2_1
X_07450_ _03986_ top.dut.bits_in_buf_next\[0\] _04037_ _04042_ vssd1 vssd1 vccd1 vccd1
+ _04043_ sky130_fd_sc_hd__a31o_1
XANTENNA__08982__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07381_ _02405_ top.dut.bits_in_buf\[0\] top.dut.bits_in_buf\[1\] vssd1 vssd1 vccd1
+ vccd1 _03985_ sky130_fd_sc_hd__o21ai_1
X_06401_ net299 _03177_ vssd1 vssd1 vccd1 vccd1 _03238_ sky130_fd_sc_hd__nor2_1
X_09120_ top.sram_interface.TRN_counter\[2\] net463 _05121_ _05130_ _05113_ vssd1
+ vssd1 vccd1 vccd1 _05136_ sky130_fd_sc_hd__a221o_1
XANTENNA__08274__A1 top.cb_syn.char_path_n\[32\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06332_ top.hist_data_o\[31\] _03194_ vssd1 vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__xor2_1
X_09051_ net1361 top.WB.CPU_DAT_O\[6\] net294 vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08002_ top.cb_syn.count\[5\] _02511_ _04497_ vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__o21ai_1
X_06263_ net478 _03129_ _03126_ _03118_ vssd1 vssd1 vccd1 vccd1 _03130_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06194_ net1213 net141 _03063_ net159 vssd1 vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__a22o_1
Xhold501 net99 vssd1 vssd1 vccd1 vccd1 net1454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 top.cb_syn.h_element\[62\] vssd1 vssd1 vccd1 vccd1 net1476 sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 top.hist_data_o\[30\] vssd1 vssd1 vccd1 vccd1 net1498 sky130_fd_sc_hd__dlygate4sd3_1
Xhold512 top.hTree.tree_reg\[24\] vssd1 vssd1 vccd1 vccd1 net1465 sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 top.histogram.total\[23\] vssd1 vssd1 vccd1 vccd1 net1487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold567 top.hTree.tree_reg\[46\] vssd1 vssd1 vccd1 vccd1 net1520 sky130_fd_sc_hd__dlygate4sd3_1
Xhold556 top.hTree.tree_reg\[41\] vssd1 vssd1 vccd1 vccd1 net1509 sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 top.histogram.total\[14\] vssd1 vssd1 vccd1 vccd1 net1531 sky130_fd_sc_hd__dlygate4sd3_1
Xhold589 top.cb_syn.h_element\[53\] vssd1 vssd1 vccd1 vccd1 net1542 sky130_fd_sc_hd__dlygate4sd3_1
X_09953_ net768 net608 vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__and2_1
X_08904_ _04157_ _04187_ vssd1 vssd1 vccd1 vccd1 _05073_ sky130_fd_sc_hd__nand2_1
XANTENNA__10053__A net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09884_ net737 net577 vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_4_4_0_clk_X clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08835_ net434 _05016_ _05017_ vssd1 vssd1 vccd1 vccd1 _05018_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout567_A net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08766_ top.path\[92\] top.path\[93\] top.path\[94\] top.path\[95\] net526 net523
+ vssd1 vssd1 vccd1 vccd1 _04949_ sky130_fd_sc_hd__mux4_1
X_05978_ top.sram_interface.init_counter\[6\] top.sram_interface.init_counter\[5\]
+ top.sram_interface.init_counter\[4\] _02913_ vssd1 vssd1 vccd1 vccd1 _02914_ sky130_fd_sc_hd__and4_1
XANTENNA__06760__A1 _03424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05563__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07717_ net429 _04278_ _04279_ net260 vssd1 vssd1 vccd1 vccd1 _04280_ sky130_fd_sc_hd__o211a_1
XANTENNA__09053__S net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08697_ top.cb_syn.zeroes\[1\] top.cb_syn.zeroes\[0\] vssd1 vssd1 vccd1 vccd1 _04892_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_0_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout734_A net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07648_ net265 _04222_ _04223_ net1099 net447 vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_0_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07579_ top.cb_syn.max_index\[4\] _04148_ vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__nand2_1
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout522_X net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09318_ top.histogram.total\[28\] net408 net326 top.histogram.total\[29\] net521
+ vssd1 vssd1 vccd1 vccd1 _05253_ sky130_fd_sc_hd__o221a_1
X_10590_ net747 net587 vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__and2_1
X_09249_ net1206 _05209_ net296 vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_header\[5\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA__06815__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_110_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_11211_ clknet_leaf_23_clk _01759_ _00566_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[113\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07537__A top.cb_syn.h_element\[63\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08640__B net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11142_ clknet_leaf_6_clk _01690_ _00497_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[44\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 ADR_O[3] sky130_fd_sc_hd__buf_2
Xoutput54 net54 vssd1 vssd1 vccd1 vccd1 ADR_O[19] sky130_fd_sc_hd__buf_2
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 DAT_O[12] sky130_fd_sc_hd__buf_2
XFILLER_110_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__09174__D net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xoutput98 net98 vssd1 vssd1 vccd1 vccd1 DAT_O[3] sky130_fd_sc_hd__buf_2
X_11073_ clknet_leaf_10_clk _01621_ _00428_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[103\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_8_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput87 net87 vssd1 vssd1 vccd1 vccd1 DAT_O[22] sky130_fd_sc_hd__buf_2
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10024_ net822 net662 vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__and2_1
XANTENNA_input30_A DAT_I[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08368__A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10926_ clknet_leaf_30_clk _01481_ _00281_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.zeroes\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_55_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10857_ clknet_leaf_46_clk _01443_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10788_ clknet_leaf_53_clk _00028_ _00207_ vssd1 vssd1 vccd1 vccd1 top.histogram.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08256__A1 top.cb_syn.char_path_n\[41\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06806__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09927__A net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11409_ clknet_leaf_98_clk _01957_ _00764_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[15\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_74_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06950_ top.compVal\[8\] top.findLeastValue.val1\[8\] net164 vssd1 vssd1 vccd1 vccd1
+ _03617_ sky130_fd_sc_hd__mux2_1
XFILLER_100_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05901_ _02875_ vssd1 vssd1 vccd1 vccd1 _02876_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06881_ top.findLeastValue.val2\[43\] net150 net123 _03582_ vssd1 vssd1 vccd1 vccd1
+ _01985_ sky130_fd_sc_hd__o22a_1
X_08620_ _04832_ _04835_ top.cb_syn.num_lefts\[6\] vssd1 vssd1 vccd1 vccd1 _04838_
+ sky130_fd_sc_hd__a21o_1
X_05832_ net550 net555 vssd1 vssd1 vccd1 vccd1 _02843_ sky130_fd_sc_hd__or2_2
XANTENNA__05545__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_6_Left_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08551_ net1358 top.cb_syn.char_path_n\[25\] net229 vssd1 vssd1 vccd1 vccd1 _01543_
+ sky130_fd_sc_hd__mux2_1
XFILLER_82_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_05763_ top.controller.state_reg\[5\] net36 vssd1 vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_85_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08482_ net1171 top.cb_syn.char_path_n\[94\] net235 vssd1 vssd1 vccd1 vccd1 _01612_
+ sky130_fd_sc_hd__mux2_1
X_07502_ top.cb_syn.char_path_n\[44\] top.cb_syn.char_path_n\[43\] top.cb_syn.char_path_n\[42\]
+ top.cb_syn.char_path_n\[41\] net400 net351 vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__mux4_1
X_05694_ net20 net417 net359 top.WB.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1 _02364_
+ sky130_fd_sc_hd__a22o_1
X_07433_ top.dut.out\[3\] net297 vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout148_A net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07364_ net1610 net135 _03547_ net126 _03974_ vssd1 vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__a32o_1
XANTENNA__05430__A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09103_ net454 _02853_ _05122_ _05120_ vssd1 vssd1 vccd1 vccd1 _05123_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_33_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout315_A net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08798__A2 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07295_ _03928_ _03929_ top.findLeastValue.sum\[22\] net274 vssd1 vssd1 vccd1 vccd1
+ _01918_ sky130_fd_sc_hd__a2bb2o_1
X_06315_ top.hist_data_o\[7\] top.hist_data_o\[6\] _03177_ vssd1 vssd1 vccd1 vccd1
+ _03178_ sky130_fd_sc_hd__and3_2
X_06246_ top.cw2\[3\] _03000_ vssd1 vssd1 vccd1 vccd1 _03113_ sky130_fd_sc_hd__nand2_1
XANTENNA__06960__S net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09034_ net1370 top.WB.CPU_DAT_O\[23\] net291 vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__mux2_1
Xhold320 top.path\[75\] vssd1 vssd1 vccd1 vccd1 net1273 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06177_ _03042_ _03044_ _03046_ net424 vssd1 vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__a31o_1
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold353 top.cb_syn.char_path\[23\] vssd1 vssd1 vccd1 vccd1 net1306 sky130_fd_sc_hd__dlygate4sd3_1
Xhold342 _01603_ vssd1 vssd1 vccd1 vccd1 net1295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold331 top.cb_syn.char_path\[118\] vssd1 vssd1 vccd1 vccd1 net1284 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09048__S net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout800 net806 vssd1 vssd1 vccd1 vccd1 net800 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout684_A net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold386 top.cb_syn.char_path\[53\] vssd1 vssd1 vccd1 vccd1 net1339 sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 net83 vssd1 vssd1 vccd1 vccd1 net1328 sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 top.histogram.sram_out\[17\] vssd1 vssd1 vccd1 vccd1 net1317 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09936_ net791 net631 vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__and2_1
Xfanout822 net823 vssd1 vssd1 vccd1 vccd1 net822 sky130_fd_sc_hd__clkbuf_2
Xhold397 top.path\[41\] vssd1 vssd1 vccd1 vccd1 net1350 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout811 net824 vssd1 vssd1 vccd1 vccd1 net811 sky130_fd_sc_hd__buf_1
Xfanout833 net834 vssd1 vssd1 vccd1 vccd1 net833 sky130_fd_sc_hd__buf_1
Xfanout855 net856 vssd1 vssd1 vccd1 vccd1 net855 sky130_fd_sc_hd__clkbuf_2
Xfanout866 net877 vssd1 vssd1 vccd1 vccd1 net866 sky130_fd_sc_hd__clkbuf_2
Xfanout844 net845 vssd1 vssd1 vccd1 vccd1 net844 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout877 net878 vssd1 vssd1 vccd1 vccd1 net877 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout851_A net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09867_ net779 net619 vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout472_X net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08183__B1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09798_ net775 net615 vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__and2_1
XANTENNA__07930__A0 top.findLeastValue.sum\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08818_ top.path\[6\] top.path\[7\] net528 vssd1 vssd1 vccd1 vccd1 _05001_ sky130_fd_sc_hd__mux2_1
X_08749_ net435 _04931_ vssd1 vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__or2_1
X_11760_ clknet_leaf_101_clk _02293_ _01115_ vssd1 vssd1 vccd1 vccd1 top.compVal\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10711_ clknet_leaf_2_clk _01310_ _00130_ vssd1 vssd1 vccd1 vccd1 top.path\[87\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_26_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11691_ clknet_leaf_62_clk _02224_ _01046_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_52_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10642_ clknet_leaf_74_clk _00051_ _00061_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.word_cnt\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10573_ net814 net654 vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__and2_1
XANTENNA__06171__A top.findLeastValue.histo_index\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11125_ clknet_leaf_29_clk _01673_ _00480_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_79_Left_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11056_ clknet_leaf_20_clk _01604_ _00411_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[86\]
+ sky130_fd_sc_hd__dfrtp_1
X_10007_ net818 net658 vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__and2_1
XANTENNA__05527__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__09421__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10909_ clknet_leaf_31_clk top.header_synthesis.next_zero_count\[4\] _00264_ vssd1
+ vssd1 vccd1 vccd1 top.cb_syn.zero_count\[4\] sky130_fd_sc_hd__dfrtp_1
X_11889_ clknet_leaf_53_clk top.dut.bits_in_buf_next\[0\] _01244_ vssd1 vssd1 vccd1
+ vccd1 top.dut.bits_in_buf\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09426__B1 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06100_ top.TRN_char_index\[5\] top.TRN_char_index\[4\] _02971_ vssd1 vssd1 vccd1
+ vccd1 _02973_ sky130_fd_sc_hd__and3_1
X_07080_ top.findLeastValue.val1\[7\] top.findLeastValue.val2\[7\] vssd1 vssd1 vccd1
+ vccd1 _03738_ sky130_fd_sc_hd__or2_1
XANTENNA__07452__A2 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06031_ net1619 top.WB.CPU_DAT_O\[4\] net355 vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08401__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07982_ top.cb_syn.zero_count\[4\] _02512_ top.cb_syn.zeroes\[5\] _02533_ vssd1 vssd1
+ vccd1 vccd1 _04485_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout118 _03551_ vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__clkbuf_4
Xfanout129 net132 vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__clkbuf_4
XFILLER_113_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09392__A net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06933_ top.findLeastValue.val2\[17\] net146 net120 _03608_ vssd1 vssd1 vccd1 vccd1
+ _01959_ sky130_fd_sc_hd__o22a_1
X_09721_ net740 net580 vssd1 vssd1 vccd1 vccd1 _00335_ sky130_fd_sc_hd__and2_1
XFILLER_79_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08500__S net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09652_ net785 net625 vssd1 vssd1 vccd1 vccd1 _00266_ sky130_fd_sc_hd__and2_1
XFILLER_103_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_06864_ top.findLeastValue.histo_index\[7\] _03572_ _03575_ vssd1 vssd1 vccd1 vccd1
+ _01996_ sky130_fd_sc_hd__o21a_1
XFILLER_55_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08603_ _04537_ _04822_ top.cb_syn.cb_enable vssd1 vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__or3b_1
X_05815_ top.sram_interface.counter_HTREE\[1\] _02827_ vssd1 vssd1 vccd1 vccd1 _02833_
+ sky130_fd_sc_hd__or2_1
X_09583_ net845 net685 vssd1 vssd1 vccd1 vccd1 _00197_ sky130_fd_sc_hd__and2_1
XANTENNA__06020__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06795_ top.findLeastValue.val1\[35\] net133 net117 top.compVal\[35\] vssd1 vssd1
+ vccd1 vccd1 _02043_ sky130_fd_sc_hd__o22a_1
XFILLER_103_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05746_ net550 top.sram_interface.word_cnt\[2\] vssd1 vssd1 vccd1 vccd1 _02781_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout265_A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08534_ net1348 top.cb_syn.char_path_n\[42\] net225 vssd1 vssd1 vccd1 vccd1 _01560_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07640__A net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08465_ net1335 top.cb_syn.char_path_n\[111\] net221 vssd1 vssd1 vccd1 vccd1 _01629_
+ sky130_fd_sc_hd__mux2_1
X_05677_ net1243 net145 _02752_ net177 vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_18_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout432_A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07416_ top.dut.bit_buf\[6\] net35 net720 vssd1 vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__mux2_1
XANTENNA__05431__Y _02539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08396_ net514 top.cb_syn.char_path_n\[11\] vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__or2_1
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07347_ _03741_ _03768_ net270 _03965_ vssd1 vssd1 vccd1 vccd1 _03966_ sky130_fd_sc_hd__o211a_1
XFILLER_109_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09017_ top.WB.CPU_DAT_O\[8\] net1369 net319 vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__mux2_1
X_07278_ top.findLeastValue.val1\[24\] top.findLeastValue.val2\[24\] _03910_ vssd1
+ vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__a21oi_1
X_06229_ _02577_ _02956_ _03095_ _03096_ vssd1 vssd1 vccd1 vccd1 _03097_ sky130_fd_sc_hd__a31o_1
Xhold150 _00047_ vssd1 vssd1 vccd1 vccd1 net1103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 top.histogram.sram_out\[6\] vssd1 vssd1 vccd1 vccd1 net1114 sky130_fd_sc_hd__dlygate4sd3_1
Xteam_05_902 vssd1 vssd1 vccd1 vccd1 team_05_902/HI gpio_out[17] sky130_fd_sc_hd__conb_1
Xteam_05_935 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] team_05_935/LO sky130_fd_sc_hd__conb_1
Xteam_05_924 vssd1 vssd1 vccd1 vccd1 gpio_oeb[4] team_05_924/LO sky130_fd_sc_hd__conb_1
Xteam_05_913 vssd1 vssd1 vccd1 vccd1 team_05_913/HI gpio_out[28] sky130_fd_sc_hd__conb_1
Xhold183 top.cb_syn.char_path\[64\] vssd1 vssd1 vccd1 vccd1 net1136 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 top.cb_syn.char_path\[69\] vssd1 vssd1 vccd1 vccd1 net1125 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 top.cb_syn.char_path\[6\] vssd1 vssd1 vccd1 vccd1 net1147 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout641 net642 vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__clkbuf_2
Xfanout630 net631 vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__clkbuf_2
Xteam_05_946 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] team_05_946/LO sky130_fd_sc_hd__conb_1
Xfanout685 net718 vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__buf_2
Xfanout663 net664 vssd1 vssd1 vccd1 vccd1 net663 sky130_fd_sc_hd__clkbuf_2
X_09919_ net743 net583 vssd1 vssd1 vccd1 vccd1 _00533_ sky130_fd_sc_hd__and2_1
Xfanout674 net675 vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__clkbuf_2
Xfanout652 net653 vssd1 vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__clkbuf_2
Xfanout696 net697 vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__buf_2
XANTENNA__05509__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ clknet_leaf_90_clk _02329_ _01167_ vssd1 vssd1 vccd1 vccd1 top.compVal\[44\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_26_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05622__X _02707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11743_ clknet_leaf_94_clk _02276_ _01098_ vssd1 vssd1 vccd1 vccd1 top.compVal\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_11674_ clknet_leaf_72_clk _02207_ _01029_ vssd1 vssd1 vccd1 vccd1 top.hTree.write_HT_fin
+ sky130_fd_sc_hd__dfrtp_4
X_10625_ net803 net643 vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__and2_1
XANTENNA__05693__B2 top.WB.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10556_ net857 net697 vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_58_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09232__B1_N top.header_synthesis.enable vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10487_ net830 net670 vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_4_12_0_clk_X clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_87_Left_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11108_ clknet_leaf_10_clk _01656_ _00463_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[10\]
+ sky130_fd_sc_hd__dfrtp_2
X_11039_ clknet_leaf_14_clk _01587_ _00394_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[69\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05600_ top.cb_syn.char_path\[13\] net557 net312 top.cb_syn.char_path\[109\] vssd1
+ vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_82_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06580_ _03354_ _03367_ _03368_ vssd1 vssd1 vccd1 vccd1 _03369_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_35_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_96_Left_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05531_ top.hTree.node_reg\[25\] net421 _02629_ _02630_ vssd1 vssd1 vccd1 vccd1 _02631_
+ sky130_fd_sc_hd__a211o_1
XFILLER_32_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05462_ net459 top.WorR net548 vssd1 vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_15_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08250_ top.cb_syn.char_path_n\[44\] net195 _04652_ vssd1 vssd1 vccd1 vccd1 _01690_
+ sky130_fd_sc_hd__o21a_1
X_08181_ top.cb_syn.char_path_n\[79\] net374 net334 top.cb_syn.char_path_n\[77\] net179
+ vssd1 vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__a221o_1
XFILLER_20_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07201_ _03659_ _03858_ vssd1 vssd1 vccd1 vccd1 _03859_ sky130_fd_sc_hd__nand2_1
X_05393_ top.cb_syn.count\[5\] vssd1 vssd1 vccd1 vccd1 _02501_ sky130_fd_sc_hd__inv_2
XFILLER_9_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07132_ top.findLeastValue.val1\[19\] top.findLeastValue.val2\[19\] vssd1 vssd1 vccd1
+ vccd1 _03790_ sky130_fd_sc_hd__and2_1
X_07063_ _03719_ _03720_ vssd1 vssd1 vccd1 vccd1 _03721_ sky130_fd_sc_hd__nor2_1
XFILLER_114_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06014_ net1586 top.WB.CPU_DAT_O\[21\] net357 vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__mux2_1
XANTENNA__06015__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07965_ top.findLeastValue.alternator_timer\[2\] net414 _02770_ vssd1 vssd1 vccd1
+ vccd1 _04473_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout382_A net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09704_ net850 net690 vssd1 vssd1 vccd1 vccd1 _00318_ sky130_fd_sc_hd__and2_1
XFILLER_68_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06916_ top.compVal\[25\] net496 net163 vssd1 vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__mux2_1
X_09635_ net803 net643 vssd1 vssd1 vccd1 vccd1 _00249_ sky130_fd_sc_hd__and2_1
XANTENNA__10769__Q top.cb_syn.h_element\[63\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07896_ net482 _04421_ vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_4_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout647_A net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06847_ top.findLeastValue.least1\[1\] net503 _03424_ vssd1 vssd1 vccd1 vccd1 _03563_
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09566_ net795 net635 vssd1 vssd1 vccd1 vccd1 _00180_ sky130_fd_sc_hd__and2_1
XFILLER_70_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06778_ top.findLeastValue.least1\[2\] net136 net118 net502 vssd1 vssd1 vccd1 vccd1
+ _02058_ sky130_fd_sc_hd__a22o_1
X_08517_ net1078 top.cb_syn.char_path_n\[59\] net232 vssd1 vssd1 vccd1 vccd1 _01577_
+ sky130_fd_sc_hd__mux2_1
X_05729_ top.findLeastValue.alternator_timer\[1\] top.findLeastValue.alternator_timer\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout435_X net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09497_ net749 net589 vssd1 vssd1 vccd1 vccd1 _00111_ sky130_fd_sc_hd__and2_1
X_08448_ net234 vssd1 vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_102_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05675__B2 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10410_ net795 net635 vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__and2_1
X_08379_ top.cb_syn.char_path_n\[105\] net391 net330 top.cb_syn.char_path_n\[106\]
+ net508 vssd1 vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__a221o_1
XANTENNA__08405__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11390_ clknet_leaf_89_clk _01938_ _00745_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[42\]
+ sky130_fd_sc_hd__dfrtp_1
X_10341_ net869 net709 vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__and2_1
XANTENNA__10236__A net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10272_ net736 net576 vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__and2_1
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold761_A top.findLeastValue.sum\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout460 net461 vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__buf_2
Xfanout471 top.controller.state_reg\[2\] vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__clkbuf_2
Xfanout493 top.hTree.state\[0\] vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__clkbuf_2
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout482 net484 vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__clkbuf_2
XFILLER_61_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11726_ clknet_leaf_121_clk _02259_ _01081_ vssd1 vssd1 vccd1 vccd1 top.path\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11657_ clknet_leaf_108_clk _02190_ _01012_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11588_ clknet_leaf_45_clk _02136_ _00943_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10608_ net808 net648 vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_40_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10539_ net867 net707 vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__and2_1
XANTENNA__07812__C1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09935__A net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08907__A2 _05072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07750_ top.hTree.tree_reg\[38\] top.findLeastValue.sum\[38\] net250 vssd1 vssd1
+ vccd1 vccd1 _04306_ sky130_fd_sc_hd__mux2_1
X_06701_ _02426_ top.findLeastValue.val2\[23\] vssd1 vssd1 vccd1 vccd1 _03489_ sky130_fd_sc_hd__nor2_1
XANTENNA__09332__A2 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07681_ net396 _04249_ vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__nand2_1
XANTENNA__08766__S1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09420_ net996 net242 _05289_ _05290_ vssd1 vssd1 vccd1 vccd1 _01454_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_48_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06632_ _03414_ _03419_ _03420_ top.findLeastValue.val1\[44\] _02407_ vssd1 vssd1
+ vccd1 vccd1 _03421_ sky130_fd_sc_hd__a32o_1
X_09351_ net1011 net240 net216 _04382_ vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__a22o_1
X_06563_ _02432_ top.findLeastValue.val1\[17\] top.findLeastValue.val1\[16\] _02433_
+ vssd1 vssd1 vccd1 vccd1 _03352_ sky130_fd_sc_hd__o22a_1
X_05514_ net1219 net139 _02616_ net175 vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__a22o_1
X_09282_ top.dut.bits_in_buf\[1\] top.dut.bits_in_buf_next\[0\] _04000_ _04041_ vssd1
+ vssd1 vccd1 vccd1 top.dut.bit_buf_next\[0\] sky130_fd_sc_hd__o31a_1
X_08302_ top.cb_syn.char_path_n\[18\] net198 _04678_ vssd1 vssd1 vccd1 vccd1 _01664_
+ sky130_fd_sc_hd__o21a_1
XFILLER_21_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08233_ top.cb_syn.char_path_n\[53\] net375 net343 top.cb_syn.char_path_n\[51\] net188
+ vssd1 vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__a221o_1
XANTENNA__08843__A1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06494_ _03285_ _03303_ vssd1 vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__nor2_1
X_05445_ top.CB_write_complete top.CB_read_complete vssd1 vssd1 vccd1 vccd1 _02553_
+ sky130_fd_sc_hd__nor2_2
XANTENNA_fanout228_A _04805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05657__B2 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout130_A net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08164_ top.cb_syn.char_path_n\[87\] net208 _04609_ vssd1 vssd1 vccd1 vccd1 _01733_
+ sky130_fd_sc_hd__o21a_1
X_05376_ top.findLeastValue.val2\[40\] vssd1 vssd1 vccd1 vccd1 _02484_ sky130_fd_sc_hd__inv_2
XFILLER_118_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08095_ top.cb_syn.char_path_n\[122\] net385 net344 top.cb_syn.char_path_n\[120\]
+ net189 vssd1 vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__a221o_1
X_07115_ top.findLeastValue.val1\[8\] top.findLeastValue.val2\[8\] vssd1 vssd1 vccd1
+ vccd1 _03773_ sky130_fd_sc_hd__xor2_1
XFILLER_119_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload70 clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 clkload70/Y sky130_fd_sc_hd__clkinv_8
X_07046_ _03685_ _03703_ vssd1 vssd1 vccd1 vccd1 _03704_ sky130_fd_sc_hd__or2_1
Xclkload92 clknet_leaf_86_clk vssd1 vssd1 vccd1 vccd1 clkload92/X sky130_fd_sc_hd__clkbuf_4
Xclkload81 clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 clkload81/X sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout597_A net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09056__S net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08997_ top.WB.CPU_DAT_O\[28\] net1107 net318 vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__mux2_1
XANTENNA__09308__C1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout764_A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07948_ top.findLeastValue.least1\[5\] top.findLeastValue.least2\[5\] _04462_ vssd1
+ vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__mux2_1
XANTENNA__05593__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_fanout552_X net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08757__S1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07879_ top.findLeastValue.sum\[12\] top.hTree.tree_reg\[12\] net283 vssd1 vssd1
+ vccd1 vccd1 _04409_ sky130_fd_sc_hd__mux2_1
X_09618_ net802 net642 vssd1 vssd1 vccd1 vccd1 _00232_ sky130_fd_sc_hd__and2_1
XFILLER_16_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10890_ clknet_leaf_110_clk _01467_ _00245_ vssd1 vssd1 vccd1 vccd1 top.translation.index\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_104_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09549_ net729 net569 vssd1 vssd1 vccd1 vccd1 _00163_ sky130_fd_sc_hd__and2_1
XFILLER_34_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05900__X _02875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06845__A0 top.findLeastValue.least1\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11511_ clknet_leaf_69_clk _02059_ _00866_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least1\[3\]
+ sky130_fd_sc_hd__dfrtp_2
X_11442_ clknet_leaf_67_clk _01990_ _00797_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.histo_index\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_109_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__10962__Q top.cb_syn.char_index\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11373_ clknet_leaf_81_clk _01921_ _00728_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07496__S1 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10324_ net766 net606 vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_115_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10255_ net866 net706 vssd1 vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__and2_1
X_10186_ net865 net705 vssd1 vssd1 vccd1 vccd1 _00800_ sky130_fd_sc_hd__and2_1
XANTENNA_clkload6_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06836__B1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11709_ clknet_leaf_117_clk _02242_ _01064_ vssd1 vssd1 vccd1 vccd1 top.path\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05639__B2 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09250__A1 top.cb_syn.char_index\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07487__S1 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold705 top.cb_syn.end_cnt\[2\] vssd1 vssd1 vccd1 vccd1 net1658 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_77_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold716 top.compVal\[29\] vssd1 vssd1 vccd1 vccd1 net1669 sky130_fd_sc_hd__dlygate4sd3_1
Xhold727 top.findLeastValue.sum\[27\] vssd1 vssd1 vccd1 vccd1 net1680 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_77_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold738 top.compVal\[17\] vssd1 vssd1 vccd1 vccd1 net1691 sky130_fd_sc_hd__dlygate4sd3_1
Xhold749 top.findLeastValue.sum\[13\] vssd1 vssd1 vccd1 vccd1 net1702 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08920_ _05081_ _05084_ _05083_ vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__o21ai_1
X_08851_ top.TRN_char_index\[6\] top.TRN_sram_complete top.TRN_char_index\[3\] top.TRN_char_index\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05034_ sky130_fd_sc_hd__or4bb_1
X_07802_ net429 _04346_ _04347_ net261 vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__o211a_1
X_05994_ top.sram_interface.init_counter\[3\] _02905_ vssd1 vssd1 vccd1 vccd1 _02922_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__05575__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08782_ top.path\[124\] net409 _04964_ vssd1 vssd1 vccd1 vccd1 _04965_ sky130_fd_sc_hd__o21a_1
X_07733_ net444 net1352 net255 top.findLeastValue.sum\[42\] _04292_ vssd1 vssd1 vccd1
+ vccd1 _01847_ sky130_fd_sc_hd__a221o_1
X_07664_ net485 _04236_ vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__nand2_1
XANTENNA__05590__A3 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_09403_ net406 _04236_ vssd1 vssd1 vccd1 vccd1 _05279_ sky130_fd_sc_hd__nand2_1
X_06615_ top.compVal\[38\] _02463_ _02464_ top.compVal\[37\] vssd1 vssd1 vccd1 vccd1
+ _03404_ sky130_fd_sc_hd__a22o_1
XANTENNA__09069__A1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout345_A net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07595_ net537 _04177_ _04180_ net531 vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__a22o_1
XANTENNA__07619__A2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09334_ net1032 net239 net218 _04450_ vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__a22o_1
X_06546_ net494 _02471_ _02472_ top.compVal\[26\] _03334_ vssd1 vssd1 vccd1 vccd1
+ _03335_ sky130_fd_sc_hd__o221a_1
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09265_ top.cb_syn.zero_count\[0\] top.cb_syn.zero_count\[1\] top.cb_syn.zero_count\[3\]
+ top.cb_syn.zero_count\[2\] vssd1 vssd1 vccd1 vccd1 _05219_ sky130_fd_sc_hd__and4_1
X_06477_ net1516 _03291_ vssd1 vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__xor2_1
XANTENNA_clkbuf_4_0_0_clk_X clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout133_X net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05428_ net549 vssd1 vssd1 vccd1 vccd1 _02536_ sky130_fd_sc_hd__inv_2
X_08216_ top.cb_syn.char_path_n\[61\] net209 _04635_ vssd1 vssd1 vccd1 vccd1 _01707_
+ sky130_fd_sc_hd__o21a_1
X_09196_ net257 _05178_ _02802_ vssd1 vssd1 vccd1 vccd1 _05179_ sky130_fd_sc_hd__or3b_1
XFILLER_119_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08147_ top.cb_syn.char_path_n\[96\] net388 net347 top.cb_syn.char_path_n\[94\] net192
+ vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__a221o_1
X_05359_ top.findLeastValue.val1\[34\] vssd1 vssd1 vccd1 vccd1 _02467_ sky130_fd_sc_hd__inv_2
X_08078_ _04133_ _04563_ _04555_ _02931_ _04562_ vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__06055__B2 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07029_ top.findLeastValue.val1\[31\] top.findLeastValue.val2\[31\] vssd1 vssd1 vccd1
+ vccd1 _03687_ sky130_fd_sc_hd__nand2_1
X_10040_ net836 net676 vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__and2_1
Xhold10 _01869_ vssd1 vssd1 vccd1 vccd1 net963 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout767_X net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold21 top.hTree.node_reg\[35\] vssd1 vssd1 vccd1 vccd1 net974 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 top.hTree.node_reg\[37\] vssd1 vssd1 vccd1 vccd1 net985 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_110_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold43 top.hTree.node_reg\[60\] vssd1 vssd1 vccd1 vccd1 net996 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 top.hTree.node_reg\[46\] vssd1 vssd1 vccd1 vccd1 net1007 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 top.hTree.tree_reg\[50\] vssd1 vssd1 vccd1 vccd1 net1018 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 net51 vssd1 vssd1 vccd1 vccd1 net1051 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 net66 vssd1 vssd1 vccd1 vccd1 net1040 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 net49 vssd1 vssd1 vccd1 vccd1 net1029 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07307__A1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10942_ clknet_leaf_33_clk _01497_ _00297_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.cb_length\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_3_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07307__B2 top.findLeastValue.sum\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10873_ clknet_leaf_35_clk _00004_ _00228_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.curr_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_42_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_502 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__06818__B1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_91_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06046__A1 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_7 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11425_ clknet_leaf_90_clk _01973_ _00780_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[31\]
+ sky130_fd_sc_hd__dfstp_2
X_11356_ clknet_leaf_97_clk _01904_ _00711_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_10307_ net803 net643 vssd1 vssd1 vccd1 vccd1 _00921_ sky130_fd_sc_hd__and2_1
XFILLER_113_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08991__A0 top.WB.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11287_ clknet_leaf_80_clk _01835_ _00642_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10238_ net833 net673 vssd1 vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__and2_1
XFILLER_86_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05557__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10169_ net840 net680 vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__and2_1
XANTENNA__05572__A3 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_44_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06400_ top.hist_data_o\[5\] _03175_ vssd1 vssd1 vccd1 vccd1 _03237_ sky130_fd_sc_hd__or2_1
X_07380_ _02405_ top.dut.bits_in_buf\[0\] top.dut.bits_in_buf\[1\] vssd1 vssd1 vccd1
+ vccd1 _03984_ sky130_fd_sc_hd__or3_1
XFILLER_22_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06331_ top.hist_data_o\[30\] top.hist_data_o\[29\] _03193_ vssd1 vssd1 vccd1 vccd1
+ _03194_ sky130_fd_sc_hd__and3_1
XANTENNA__06809__B1 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06262_ top.cb_syn.char_index\[1\] top.cb_syn.char_index\[0\] net561 _03128_ vssd1
+ vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__a31o_1
XANTENNA__08274__A2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09050_ net1087 top.WB.CPU_DAT_O\[7\] net294 vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08001_ _02499_ top.cb_syn.zeroes\[7\] _04497_ vssd1 vssd1 vccd1 vccd1 _04504_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_59_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06193_ _03062_ _03051_ _03047_ _03057_ vssd1 vssd1 vccd1 vccd1 _03063_ sky130_fd_sc_hd__or4bb_1
Xhold502 top.cb_syn.char_path\[113\] vssd1 vssd1 vccd1 vccd1 net1455 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_102_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold535 top.cb_syn.check_right vssd1 vssd1 vccd1 vccd1 net1488 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08431__C1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold524 top.hist_data_o\[20\] vssd1 vssd1 vccd1 vccd1 net1477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 _01829_ vssd1 vssd1 vccd1 vccd1 net1466 sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 top.cb_syn.curr_index\[3\] vssd1 vssd1 vccd1 vccd1 net1521 sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 top.histogram.sram_out\[22\] vssd1 vssd1 vccd1 vccd1 net1499 sky130_fd_sc_hd__dlygate4sd3_1
X_09952_ net768 net608 vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__and2_1
Xhold579 top.hTree.node_reg\[26\] vssd1 vssd1 vccd1 vccd1 net1532 sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 _01846_ vssd1 vssd1 vccd1 vccd1 net1510 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08982__A0 top.WB.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__05428__A net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08903_ top.cb_syn.max_index\[7\] _05070_ _05072_ vssd1 vssd1 vccd1 vccd1 _01393_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__10053__B net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_117_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06023__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09883_ net737 net577 vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__and2_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08834_ top.path\[36\] net410 net328 top.path\[37\] net522 vssd1 vssd1 vccd1 vccd1
+ _05017_ sky130_fd_sc_hd__o221a_1
XANTENNA__06958__S net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08765_ net433 _04946_ _04947_ vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__o21a_1
X_05977_ top.sram_interface.init_counter\[3\] _02902_ _02911_ vssd1 vssd1 vccd1 vccd1
+ _02913_ sky130_fd_sc_hd__and3_1
X_07716_ net488 _04277_ vssd1 vssd1 vccd1 vccd1 _04279_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_28_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08696_ _04877_ _04885_ _04891_ _04875_ top.cb_syn.zeroes\[2\] vssd1 vssd1 vccd1
+ vccd1 _01483_ sky130_fd_sc_hd__a32o_1
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07647_ net491 _04220_ vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout250_X net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout727_A net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07578_ net532 top.cb_syn.h_element\[49\] net539 top.cb_syn.h_element\[58\] _04135_
+ vssd1 vssd1 vccd1 vccd1 _04166_ sky130_fd_sc_hd__a221o_1
XANTENNA__05720__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07789__S net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06529_ _03319_ vssd1 vssd1 vccd1 vccd1 _03320_ sky130_fd_sc_hd__inv_2
X_09317_ net432 _05251_ vssd1 vssd1 vccd1 vccd1 _05252_ sky130_fd_sc_hd__or2_1
XFILLER_41_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout515_X net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09248_ top.header_synthesis.header\[5\] top.cb_syn.char_index\[5\] net518 vssd1
+ vssd1 vccd1 vccd1 _05209_ sky130_fd_sc_hd__mux2_1
X_09179_ _04536_ _05169_ _05170_ vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__or3_1
Xclkbuf_4_10_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_10_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08921__B _05072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11210_ clknet_leaf_7_clk _01758_ _00565_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[112\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06028__A1 top.WB.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__08973__A0 top.WB.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11141_ clknet_leaf_4_clk _01689_ _00496_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[43\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 ADR_O[4] sky130_fd_sc_hd__buf_2
Xoutput55 net55 vssd1 vssd1 vccd1 vccd1 ADR_O[20] sky130_fd_sc_hd__buf_2
XFILLER_1_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput88 net88 vssd1 vssd1 vccd1 vccd1 DAT_O[23] sky130_fd_sc_hd__buf_2
X_11072_ clknet_leaf_12_clk _01620_ _00427_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[102\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_8_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput99 net99 vssd1 vssd1 vccd1 vccd1 DAT_O[4] sky130_fd_sc_hd__buf_2
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 DAT_O[13] sky130_fd_sc_hd__buf_2
XFILLER_102_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05539__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10023_ net820 net660 vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__and2_1
XANTENNA__06200__B2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input23_A DAT_I[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05554__A3 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10925_ clknet_leaf_38_clk _01480_ _00280_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.left_check
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_55_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10856_ clknet_leaf_78_clk _01442_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05711__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10787_ clknet_leaf_47_clk _01386_ _00206_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__09205__A1 top.CB_read_complete vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09927__B net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06019__A1 top.WB.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11408_ clknet_leaf_99_clk _01956_ _00763_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[14\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07767__A1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08964__A0 top.WB.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11339_ clknet_leaf_53_clk _01887_ _00694_ vssd1 vssd1 vccd1 vccd1 top.dut.out\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09943__A net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05900_ _02554_ _02867_ _02870_ _02874_ _02863_ vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__a311o_2
X_06880_ top.compVal\[43\] top.findLeastValue.val1\[43\] net164 vssd1 vssd1 vccd1
+ vccd1 _03582_ sky130_fd_sc_hd__mux2_1
X_05831_ _02840_ _02842_ vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__and2_1
XANTENNA__05535__X _02634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08550_ net1120 top.cb_syn.char_path_n\[26\] net231 vssd1 vssd1 vccd1 vccd1 _01544_
+ sky130_fd_sc_hd__mux2_1
XFILLER_54_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05950__A0 top.WB.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05762_ top.compVal\[32\] net173 _02783_ top.WB.CPU_DAT_O\[0\] vssd1 vssd1 vccd1
+ vccd1 _02317_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_85_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08481_ net1111 top.cb_syn.char_path_n\[95\] net233 vssd1 vssd1 vccd1 vccd1 _01613_
+ sky130_fd_sc_hd__mux2_1
X_07501_ top.cb_syn.char_path_n\[40\] top.cb_syn.char_path_n\[39\] top.cb_syn.char_path_n\[38\]
+ top.cb_syn.char_path_n\[37\] net399 net350 vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__mux4_1
X_05693_ net21 net415 net308 top.WB.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1 _02365_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07750__X _04306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07432_ net1486 net297 _03999_ _04028_ _04025_ vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__a221o_1
XANTENNA__05702__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07363_ top.cw1\[6\] net167 _03553_ top.findLeastValue.histo_index\[6\] vssd1 vssd1
+ vccd1 vccd1 _03974_ sky130_fd_sc_hd__a22o_1
X_09102_ top.sram_interface.zero_cnt\[2\] _02449_ _02450_ _02763_ vssd1 vssd1 vccd1
+ vccd1 _05122_ sky130_fd_sc_hd__nor4_1
XTAP_TAPCELL_ROW_33_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06018__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06314_ _03174_ _03176_ vssd1 vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__and2_1
X_07294_ net269 _03925_ vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout210_A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06245_ net502 net412 _03111_ net549 _02573_ vssd1 vssd1 vccd1 vccd1 _03112_ sky130_fd_sc_hd__o2111a_1
X_09033_ net1228 top.WB.CPU_DAT_O\[24\] net292 vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_107_Left_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06176_ _02536_ _02573_ _02996_ _03045_ vssd1 vssd1 vccd1 vccd1 _03046_ sky130_fd_sc_hd__or4_1
Xhold310 top.cb_syn.end_check vssd1 vssd1 vccd1 vccd1 net1263 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout308_A net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08955__A0 top.WB.CPU_DAT_O\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold343 top.hTree.nulls\[52\] vssd1 vssd1 vccd1 vccd1 net1296 sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 top.cb_syn.char_path\[103\] vssd1 vssd1 vccd1 vccd1 net1285 sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 top.path\[84\] vssd1 vssd1 vccd1 vccd1 net1274 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07758__A1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold354 net45 vssd1 vssd1 vccd1 vccd1 net1307 sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 top.cb_syn.char_path\[114\] vssd1 vssd1 vccd1 vccd1 net1329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold387 top.hTree.nulls\[59\] vssd1 vssd1 vccd1 vccd1 net1340 sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 top.path\[103\] vssd1 vssd1 vccd1 vccd1 net1318 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout801 net802 vssd1 vssd1 vccd1 vccd1 net801 sky130_fd_sc_hd__clkbuf_2
X_09935_ net791 net631 vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__and2_1
Xfanout823 net824 vssd1 vssd1 vccd1 vccd1 net823 sky130_fd_sc_hd__clkbuf_2
Xhold398 net76 vssd1 vssd1 vccd1 vccd1 net1351 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout834 net835 vssd1 vssd1 vccd1 vccd1 net834 sky130_fd_sc_hd__clkbuf_2
Xfanout812 net813 vssd1 vssd1 vccd1 vccd1 net812 sky130_fd_sc_hd__clkbuf_2
Xfanout856 net857 vssd1 vssd1 vccd1 vccd1 net856 sky130_fd_sc_hd__buf_2
Xfanout867 net877 vssd1 vssd1 vccd1 vccd1 net867 sky130_fd_sc_hd__clkbuf_2
X_09866_ net777 net617 vssd1 vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__and2_1
Xfanout845 net878 vssd1 vssd1 vccd1 vccd1 net845 sky130_fd_sc_hd__buf_2
XFILLER_58_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout878 net879 vssd1 vssd1 vccd1 vccd1 net878 sky130_fd_sc_hd__buf_2
XFILLER_112_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_08817_ net436 _04999_ _04998_ vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_116_Left_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout465_X net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout844_A net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09797_ net774 net614 vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__and2_1
XANTENNA__05536__A3 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05941__A0 top.WB.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08748_ top.path\[70\] top.path\[71\] net527 vssd1 vssd1 vccd1 vccd1 _04931_ sky130_fd_sc_hd__mux2_1
X_08679_ top.cb_syn.zeroes\[4\] _04878_ vssd1 vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__nand2_1
XFILLER_26_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ clknet_leaf_1_clk _01309_ _00129_ vssd1 vssd1 vccd1 vccd1 top.path\[86\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11690_ clknet_leaf_62_clk _02223_ _01045_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08408__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10641_ clknet_leaf_65_clk _00050_ _00060_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.word_cnt\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10572_ net752 net592 vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__and2_1
XANTENNA__08946__A0 top.WB.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08410__A2 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11124_ clknet_leaf_29_clk _01672_ _00479_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11055_ clknet_leaf_20_clk net1295 _00410_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[85\]
+ sky130_fd_sc_hd__dfrtp_1
X_10006_ net820 net660 vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__and2_1
XANTENNA__05932__A0 top.WB.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10908_ clknet_leaf_31_clk top.header_synthesis.next_zero_count\[3\] _00263_ vssd1
+ vssd1 vccd1 vccd1 top.cb_syn.zero_count\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_72_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11888_ clknet_leaf_37_clk top.header_synthesis.next_write_num_lefts _01243_ vssd1
+ vssd1 vccd1 vccd1 top.header_synthesis.write_num_lefts sky130_fd_sc_hd__dfrtp_1
X_10839_ clknet_leaf_79_clk _01425_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_80_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05463__A2 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06030_ net1496 top.WB.CPU_DAT_O\[5\] net355 vssd1 vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__mux2_1
XANTENNA__08937__A0 top.WB.CPU_DAT_O\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08988__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07981_ _02509_ top.cb_syn.zero_count\[7\] top.cb_syn.zero_count\[6\] _02510_ vssd1
+ vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__o22a_1
XFILLER_99_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout119 _03551_ vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06932_ top.compVal\[17\] top.findLeastValue.val1\[17\] net161 vssd1 vssd1 vccd1
+ vccd1 _03608_ sky130_fd_sc_hd__mux2_1
XANTENNA__06963__A2 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09720_ net740 net580 vssd1 vssd1 vccd1 vccd1 _00334_ sky130_fd_sc_hd__and2_1
X_09651_ net785 net625 vssd1 vssd1 vccd1 vccd1 _00265_ sky130_fd_sc_hd__and2_1
XFILLER_94_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06863_ top.findLeastValue.histo_index\[8\] _03575_ _03576_ _03574_ vssd1 vssd1 vccd1
+ vccd1 _01997_ sky130_fd_sc_hd__a22o_1
XANTENNA__05518__A3 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08602_ _02929_ _04801_ _04800_ _04543_ vssd1 vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__o211a_1
X_05814_ _02829_ _02832_ vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__nor2_1
XFILLER_67_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09582_ net793 net633 vssd1 vssd1 vccd1 vccd1 _00196_ sky130_fd_sc_hd__and2_1
X_06794_ top.findLeastValue.val1\[36\] net131 net115 top.compVal\[36\] vssd1 vssd1
+ vccd1 vccd1 _02044_ sky130_fd_sc_hd__o22a_1
XFILLER_82_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05745_ net556 _02779_ net424 vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__a21o_1
X_08533_ net1457 top.cb_syn.char_path_n\[43\] net220 vssd1 vssd1 vccd1 vccd1 _01561_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout258_A net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08464_ net1331 top.cb_syn.char_path_n\[112\] net222 vssd1 vssd1 vccd1 vccd1 _01630_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_18_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05676_ top.histogram.sram_out\[1\] net364 net419 top.hTree.node_reg\[1\] _02751_
+ vssd1 vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__a221o_1
X_07415_ _03989_ _03991_ _03987_ vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__mux2_1
XANTENNA__10059__A net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08395_ top.cb_syn.char_path_n\[6\] net330 _04753_ vssd1 vssd1 vccd1 vccd1 _04754_
+ sky130_fd_sc_hd__a21o_1
XFILLER_11_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07346_ _03741_ _03768_ vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__nand2_1
XANTENNA__09848__A net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07523__S0 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07277_ net1661 net273 _03864_ _03915_ vssd1 vssd1 vccd1 vccd1 _01922_ sky130_fd_sc_hd__a22o_1
X_09016_ top.WB.CPU_DAT_O\[9\] net1446 net319 vssd1 vssd1 vccd1 vccd1 _01296_ sky130_fd_sc_hd__mux2_1
X_06228_ _02957_ net561 vssd1 vssd1 vccd1 vccd1 _03096_ sky130_fd_sc_hd__and2b_1
XANTENNA__08928__A0 top.WB.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_05_903 vssd1 vssd1 vccd1 vccd1 team_05_903/HI gpio_out[18] sky130_fd_sc_hd__conb_1
X_06159_ top.TRN_char_index\[5\] _02972_ vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__nor2_1
Xhold151 top.cb_syn.char_path\[71\] vssd1 vssd1 vccd1 vccd1 net1104 sky130_fd_sc_hd__dlygate4sd3_1
Xhold140 top.path\[19\] vssd1 vssd1 vccd1 vccd1 net1093 sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 top.histogram.sram_out\[4\] vssd1 vssd1 vccd1 vccd1 net1115 sky130_fd_sc_hd__dlygate4sd3_1
Xteam_05_925 vssd1 vssd1 vccd1 vccd1 gpio_oeb[5] team_05_925/LO sky130_fd_sc_hd__conb_1
Xteam_05_936 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] team_05_936/LO sky130_fd_sc_hd__conb_1
XANTENNA__09583__A net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold173 top.cb_syn.char_path\[4\] vssd1 vssd1 vccd1 vccd1 net1126 sky130_fd_sc_hd__dlygate4sd3_1
Xteam_05_914 vssd1 vssd1 vccd1 vccd1 team_05_914/HI gpio_out[29] sky130_fd_sc_hd__conb_1
Xhold195 top.histogram.sram_out\[9\] vssd1 vssd1 vccd1 vccd1 net1148 sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 top.path\[90\] vssd1 vssd1 vccd1 vccd1 net1137 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout620 net626 vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__clkbuf_2
Xfanout642 net646 vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__buf_1
Xfanout631 net646 vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__clkbuf_2
Xteam_05_947 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] team_05_947/LO sky130_fd_sc_hd__conb_1
X_09918_ net742 net582 vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__and2_1
XANTENNA__09353__B1 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout664 net719 vssd1 vssd1 vccd1 vccd1 net664 sky130_fd_sc_hd__buf_2
Xfanout653 net664 vssd1 vssd1 vccd1 vccd1 net653 sky130_fd_sc_hd__clkbuf_2
Xfanout675 net719 vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__clkbuf_2
Xfanout697 net718 vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__clkbuf_2
Xfanout686 net689 vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__clkbuf_2
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__07903__A1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09849_ net741 net581 vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__and2_1
XANTENNA__07903__B2 top.findLeastValue.sum\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ clknet_leaf_90_clk _02328_ _01166_ vssd1 vssd1 vccd1 vccd1 top.compVal\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07667__B1 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11742_ clknet_leaf_94_clk _02275_ _01097_ vssd1 vssd1 vccd1 vccd1 top.compVal\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_41_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11673_ clknet_leaf_43_clk _02206_ _01028_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10624_ net805 net645 vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__and2_1
X_10555_ net844 net684 vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__and2_1
XANTENNA__11796__Q top.controller.state_reg\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10486_ net835 net675 vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_118_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08919__B1 _05072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09493__A net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11107_ clknet_leaf_10_clk _01655_ _00462_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11038_ clknet_leaf_14_clk _01586_ _00393_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[68\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05530_ net456 top.hTree.node_reg\[57\] _02583_ net365 top.histogram.sram_out\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02630_ sky130_fd_sc_hd__a32o_1
X_05461_ net453 top.histogram.wr_r_en\[1\] top.histogram.wr_r_en\[0\] net366 vssd1
+ vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_15_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05392_ top.cb_syn.count\[6\] vssd1 vssd1 vccd1 vccd1 _02500_ sky130_fd_sc_hd__inv_2
X_08180_ top.cb_syn.char_path_n\[79\] net197 _04617_ vssd1 vssd1 vccd1 vccd1 _01725_
+ sky130_fd_sc_hd__o21a_1
XFILLER_32_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07200_ top.findLeastValue.val1\[44\] top.findLeastValue.val2\[44\] vssd1 vssd1 vccd1
+ vccd1 _03858_ sky130_fd_sc_hd__or2_1
X_07131_ top.findLeastValue.val1\[19\] top.findLeastValue.val2\[19\] vssd1 vssd1 vccd1
+ vccd1 _03789_ sky130_fd_sc_hd__nor2_1
XANTENNA__06094__C1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07062_ top.findLeastValue.val1\[12\] top.findLeastValue.val2\[12\] vssd1 vssd1 vccd1
+ vccd1 _03720_ sky130_fd_sc_hd__nor2_1
X_06013_ net1587 top.WB.CPU_DAT_O\[22\] net358 vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_93_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08511__S net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07964_ top.findLeastValue.alternator_timer\[1\] top.findLeastValue.alternator_timer\[0\]
+ _03566_ top.findLeastValue.alternator_timer\[2\] vssd1 vssd1 vccd1 vccd1 _04472_
+ sky130_fd_sc_hd__a31o_1
X_09703_ net801 net641 vssd1 vssd1 vccd1 vccd1 _00317_ sky130_fd_sc_hd__and2_1
X_06915_ top.findLeastValue.val2\[26\] net148 net121 _03599_ vssd1 vssd1 vccd1 vccd1
+ _01968_ sky130_fd_sc_hd__o22a_1
X_07895_ top.hTree.tree_reg\[9\] top.findLeastValue.sum\[9\] net247 vssd1 vssd1 vccd1
+ vccd1 _04422_ sky130_fd_sc_hd__mux2_1
XANTENNA__09335__B1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout375_A net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06846_ _02478_ net152 net126 _03562_ vssd1 vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09634_ net759 net599 vssd1 vssd1 vccd1 vccd1 _00248_ sky130_fd_sc_hd__and2_1
XANTENNA__06966__S net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07361__A2 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09565_ net794 net634 vssd1 vssd1 vccd1 vccd1 _00179_ sky130_fd_sc_hd__and2_1
X_06777_ top.findLeastValue.least1\[3\] net136 net118 top.findLeastValue.histo_index\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout542_A net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08516_ net1368 top.cb_syn.char_path_n\[60\] net231 vssd1 vssd1 vccd1 vccd1 _01578_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07370__B net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05728_ top.findLeastValue.histo_index\[8\] _02547_ vssd1 vssd1 vccd1 vccd1 _02763_
+ sky130_fd_sc_hd__or2_2
XFILLER_70_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09496_ net755 net595 vssd1 vssd1 vccd1 vccd1 _00110_ sky130_fd_sc_hd__and2_1
XFILLER_23_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08447_ _04133_ _04562_ vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__nor2_1
XANTENNA__05602__C net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout330_X net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05659_ net1454 net138 _02737_ net176 vssd1 vssd1 vccd1 vccd1 _02374_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout807_A net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05675__A2 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08378_ top.cb_syn.char_path_n\[107\] top.cb_syn.char_path_n\[108\] net514 vssd1
+ vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__mux2_1
X_07329_ net269 _03944_ _03953_ net274 net1682 vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__a32o_1
X_10340_ net874 net714 vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__and2_1
X_10271_ net726 net566 vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__and2_1
XANTENNA__10236__B net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout450 _02404_ vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__clkbuf_4
Xfanout461 net462 vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__clkbuf_2
XFILLER_93_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xfanout472 net477 vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__clkbuf_4
Xfanout483 net484 vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout494 top.compVal\[27\] vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__buf_2
XANTENNA__09252__S net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06876__S net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_11725_ clknet_leaf_120_clk _02258_ _01080_ vssd1 vssd1 vccd1 vccd1 top.path\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05666__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11656_ clknet_leaf_108_clk _02189_ _01011_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11587_ clknet_leaf_15_clk _02135_ _00942_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10607_ net729 net569 vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_40_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10538_ net867 net707 vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__and2_1
XFILLER_6_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05823__C1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09935__B net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10469_ net729 net569 vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__and2_1
XFILLER_111_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_111_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06700_ _02430_ top.findLeastValue.val2\[19\] vssd1 vssd1 vccd1 vccd1 _03488_ sky130_fd_sc_hd__nand2_1
XANTENNA__07879__A0 top.findLeastValue.sum\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05543__X _02641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07680_ top.findLeastValue.least2\[5\] top.hTree.tree_reg\[51\] net281 vssd1 vssd1
+ vccd1 vccd1 _04249_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06631_ _03393_ _03418_ _03411_ vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06087__A top.cb_syn.char_index\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09350_ net987 net240 net216 _04386_ vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__a22o_1
X_06562_ _03344_ _03346_ _03349_ _03345_ vssd1 vssd1 vccd1 vccd1 _03351_ sky130_fd_sc_hd__or4b_1
X_09281_ net1670 _05228_ _05230_ _05213_ vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_zero_count\[7\]
+ sky130_fd_sc_hd__a22o_1
X_05513_ top.histogram.sram_out\[28\] net365 _02614_ _02615_ vssd1 vssd1 vccd1 vccd1
+ _02616_ sky130_fd_sc_hd__a211o_1
X_08301_ top.cb_syn.char_path_n\[19\] net375 net335 top.cb_syn.char_path_n\[17\] net180
+ vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__a221o_1
XANTENNA__06303__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08232_ top.cb_syn.char_path_n\[53\] net205 _04643_ vssd1 vssd1 vccd1 vccd1 _01699_
+ sky130_fd_sc_hd__o21a_1
X_06493_ top.histogram.total\[17\] _03284_ net1489 vssd1 vssd1 vccd1 vccd1 _03303_
+ sky130_fd_sc_hd__a21oi_1
X_05444_ _02549_ net368 _02551_ net468 vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__o211a_1
XANTENNA__06759__C_N _03545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08163_ top.cb_syn.char_path_n\[88\] net387 net346 top.cb_syn.char_path_n\[86\] net191
+ vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__a221o_1
X_05375_ top.findLeastValue.val2\[42\] vssd1 vssd1 vccd1 vccd1 _02483_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout123_A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08094_ top.cb_syn.char_path_n\[122\] net206 _04574_ vssd1 vssd1 vccd1 vccd1 _01768_
+ sky130_fd_sc_hd__o21a_1
X_07114_ _03764_ _03767_ _03771_ _03740_ _03739_ vssd1 vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__o2111ai_2
XFILLER_109_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload60 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 clkload60/Y sky130_fd_sc_hd__bufinv_16
Xclkload71 clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 clkload71/Y sky130_fd_sc_hd__clkinv_2
X_07045_ _03695_ _03696_ _03698_ _03702_ vssd1 vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__or4_1
XANTENNA__08359__A1 _02504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload93 clknet_leaf_87_clk vssd1 vssd1 vccd1 vccd1 clkload93/Y sky130_fd_sc_hd__inv_6
Xclkload82 clknet_leaf_91_clk vssd1 vssd1 vccd1 vccd1 clkload82/Y sky130_fd_sc_hd__inv_4
XANTENNA_fanout492_A net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__07365__B net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08996_ top.WB.CPU_DAT_O\[29\] net1282 net317 vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__mux2_1
XFILLER_102_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07947_ net1547 _04463_ _04461_ vssd1 vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__mux2_1
XANTENNA__06790__B1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout757_A net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07878_ net440 net1595 net252 top.findLeastValue.sum\[13\] _04408_ vssd1 vssd1 vccd1
+ vccd1 _01818_ sky130_fd_sc_hd__a221o_1
X_09617_ net798 net638 vssd1 vssd1 vccd1 vccd1 _00231_ sky130_fd_sc_hd__and2_1
X_06829_ top.findLeastValue.val1\[1\] net130 net114 net1693 vssd1 vssd1 vccd1 vccd1
+ _02009_ sky130_fd_sc_hd__o22a_1
XFILLER_28_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08819__C1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09548_ net733 net573 vssd1 vssd1 vccd1 vccd1 _00162_ sky130_fd_sc_hd__and2_1
XANTENNA__08295__B1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11510_ clknet_leaf_69_clk _02058_ _00865_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least1\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08834__A2 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09479_ net723 net563 vssd1 vssd1 vccd1 vccd1 _00093_ sky130_fd_sc_hd__and2_1
XANTENNA__05648__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11441_ clknet_leaf_67_clk _01989_ _00796_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.histo_index\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_109_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11372_ clknet_leaf_80_clk _01920_ _00727_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_109_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10323_ net766 net606 vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_115_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05820__A2 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10254_ net862 net702 vssd1 vssd1 vccd1 vccd1 _00868_ sky130_fd_sc_hd__and2_1
XANTENNA__05628__X _02712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10185_ net864 net704 vssd1 vssd1 vccd1 vccd1 _00799_ sky130_fd_sc_hd__and2_1
XFILLER_38_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout280 net282 vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__clkbuf_4
Xfanout291 net292 vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08387__A _02504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08674__X _04875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08825__A2 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06836__A1 top.findLeastValue.least2\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11708_ clknet_leaf_114_clk _02241_ _01063_ vssd1 vssd1 vccd1 vccd1 top.path\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11639_ clknet_leaf_56_clk top.dut.bit_buf_next\[11\] _00994_ vssd1 vssd1 vccd1 vccd1
+ top.dut.bit_buf\[11\] sky130_fd_sc_hd__dfrtp_1
Xhold717 top.cb_syn.zero_count\[7\] vssd1 vssd1 vccd1 vccd1 net1670 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap403 _03995_ vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_77_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold706 top.findLeastValue.sum\[38\] vssd1 vssd1 vccd1 vccd1 net1659 sky130_fd_sc_hd__dlygate4sd3_1
Xhold728 top.findLeastValue.sum\[9\] vssd1 vssd1 vccd1 vccd1 net1681 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_3_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold739 top.cb_syn.cb_length\[4\] vssd1 vssd1 vccd1 vccd1 net1692 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08850_ _02791_ _05032_ vssd1 vssd1 vccd1 vccd1 _05033_ sky130_fd_sc_hd__nand2_1
X_07801_ net488 _04345_ vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__or2_1
X_05993_ _02906_ _02921_ vssd1 vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__nor2_1
XANTENNA__06772__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08781_ top.path\[125\] net327 _04963_ net433 net520 vssd1 vssd1 vccd1 vccd1 _04964_
+ sky130_fd_sc_hd__o221a_1
X_07732_ net429 _04290_ _04291_ net260 vssd1 vssd1 vccd1 vccd1 _04292_ sky130_fd_sc_hd__o211a_1
X_07663_ top.findLeastValue.least1\[0\] net248 _04234_ vssd1 vssd1 vccd1 vccd1 _04236_
+ sky130_fd_sc_hd__a21oi_1
X_09402_ net981 net245 _05278_ vssd1 vssd1 vccd1 vccd1 _01448_ sky130_fd_sc_hd__o21a_1
X_06614_ _02406_ top.findLeastValue.val1\[45\] top.findLeastValue.val1\[44\] _02407_
+ vssd1 vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__o22a_1
X_07594_ _04179_ vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__inv_2
X_09333_ net1000 net236 net215 _04454_ vssd1 vssd1 vccd1 vccd1 _01395_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout240_A net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout338_A net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06545_ top.compVal\[24\] _03332_ _03333_ vssd1 vssd1 vccd1 vccd1 _03334_ sky130_fd_sc_hd__a21o_1
X_09264_ _05213_ _05217_ _05218_ _05214_ top.cb_syn.zero_count\[2\] vssd1 vssd1 vccd1
+ vccd1 top.header_synthesis.next_zero_count\[2\] sky130_fd_sc_hd__a32o_1
X_06476_ _03292_ net1553 vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__nor2_1
X_08215_ top.cb_syn.char_path_n\[62\] net388 net348 top.cb_syn.char_path_n\[60\] net193
+ vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__a221o_1
X_09195_ _03325_ _05059_ _05177_ vssd1 vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__and3_1
X_05427_ net485 vssd1 vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__inv_2
X_08146_ top.cb_syn.char_path_n\[96\] net209 _04600_ vssd1 vssd1 vccd1 vccd1 _01742_
+ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout126_X net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05358_ top.findLeastValue.val1\[35\] vssd1 vssd1 vccd1 vccd1 _02466_ sky130_fd_sc_hd__inv_2
X_08077_ net530 net538 vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__or2_1
X_07028_ top.findLeastValue.val1\[31\] top.findLeastValue.val2\[31\] vssd1 vssd1 vccd1
+ vccd1 _03686_ sky130_fd_sc_hd__and2_1
Xhold11 top.sram_interface.init_counter\[19\] vssd1 vssd1 vccd1 vccd1 net964 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 top.hTree.node_reg\[36\] vssd1 vssd1 vccd1 vccd1 net975 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08752__A1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout662_X net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold33 top.hTree.node_reg\[49\] vssd1 vssd1 vccd1 vccd1 net986 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 top.hTree.node_reg\[16\] vssd1 vssd1 vccd1 vccd1 net997 sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ top.WB.CPU_DAT_O\[13\] net1127 net322 vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__mux2_1
Xhold55 top.hTree.node_reg\[13\] vssd1 vssd1 vccd1 vccd1 net1008 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 net56 vssd1 vssd1 vccd1 vccd1 net1030 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 net53 vssd1 vssd1 vccd1 vccd1 net1052 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 net52 vssd1 vssd1 vccd1 vccd1 net1041 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 top.hTree.node_reg\[45\] vssd1 vssd1 vccd1 vccd1 net1019 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10941_ clknet_leaf_35_clk _01496_ _00296_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.cb_length\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_3_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10872_ clknet_leaf_41_clk _00003_ _00227_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.curr_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_31_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_117_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_117_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08807__A2 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11424_ clknet_leaf_81_clk _01972_ _00779_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[30\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_8 top.WB.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11355_ clknet_leaf_91_clk _01903_ _00710_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_10306_ net803 net643 vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__and2_1
XFILLER_98_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11286_ clknet_leaf_84_clk _01834_ _00641_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07286__A _03782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10237_ net832 net672 vssd1 vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_72_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10168_ net840 net680 vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__and2_1
XFILLER_86_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10099_ net827 net667 vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_108_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_108_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_22_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06330_ top.hist_data_o\[28\] top.hist_data_o\[27\] _03192_ vssd1 vssd1 vccd1 vccd1
+ _03193_ sky130_fd_sc_hd__and3_1
X_06261_ top.cb_syn.char_index\[1\] _03127_ _02557_ top.cb_syn.curr_index\[3\] vssd1
+ vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_20_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08000_ top.cb_syn.count\[5\] _02511_ _02512_ top.cb_syn.count\[4\] _04502_ vssd1
+ vssd1 vccd1 vccd1 _04503_ sky130_fd_sc_hd__a221oi_1
X_06192_ top.cb_syn.curr_index\[6\] _02558_ _02579_ _03059_ _03061_ vssd1 vssd1 vccd1
+ vccd1 _03062_ sky130_fd_sc_hd__a221o_1
Xhold503 top.hTree.nullSumIndex\[2\] vssd1 vssd1 vccd1 vccd1 net1456 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08431__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold525 top.histogram.total\[26\] vssd1 vssd1 vccd1 vccd1 net1478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold536 top.histogram.total\[18\] vssd1 vssd1 vccd1 vccd1 net1489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold514 top.histogram.sram_out\[5\] vssd1 vssd1 vccd1 vccd1 net1467 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold547 top.hTree.nullSumIndex\[5\] vssd1 vssd1 vccd1 vccd1 net1500 sky130_fd_sc_hd__dlygate4sd3_1
X_09951_ net738 net578 vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__and2_1
Xhold558 top.histogram.total\[25\] vssd1 vssd1 vccd1 vccd1 net1511 sky130_fd_sc_hd__dlygate4sd3_1
Xhold569 top.hTree.tree_reg\[43\] vssd1 vssd1 vccd1 vccd1 net1522 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08902_ top.hTree.finish_check _04188_ _05061_ _05071_ vssd1 vssd1 vccd1 vccd1 _05072_
+ sky130_fd_sc_hd__o211a_4
X_09882_ net736 net576 vssd1 vssd1 vccd1 vccd1 _00496_ sky130_fd_sc_hd__and2_1
XFILLER_111_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout190_A net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08833_ top.path\[38\] top.path\[39\] net528 vssd1 vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__mux2_1
X_05976_ top.sram_interface.init_counter\[3\] _02911_ vssd1 vssd1 vccd1 vccd1 _02912_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__07643__B net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08764_ top.path\[88\] net408 net327 top.path\[89\] net436 vssd1 vssd1 vccd1 vccd1
+ _04947_ sky130_fd_sc_hd__o221a_1
X_07715_ top.hTree.tree_reg\[45\] top.findLeastValue.sum\[45\] net250 vssd1 vssd1
+ vccd1 vccd1 _04278_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08695_ _02514_ _04876_ vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07646_ net491 _04221_ vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__nand2_1
XFILLER_53_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout622_A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07577_ top.cb_syn.h_element\[58\] top.cb_syn.h_element\[49\] _04145_ vssd1 vssd1
+ vccd1 vccd1 _04165_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout243_X net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05720__B2 top.WB.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06528_ top.dut.out\[2\] top.dut.out\[1\] _03318_ top.dut.out\[3\] vssd1 vssd1 vccd1
+ vccd1 _03319_ sky130_fd_sc_hd__and4b_1
X_09316_ top.histogram.total\[30\] top.histogram.total\[31\] net524 vssd1 vssd1 vccd1
+ vccd1 _05251_ sky130_fd_sc_hd__mux2_1
X_09247_ net1105 _05208_ net296 vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_header\[4\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout508_X net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout410_X net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06459_ _03268_ _03281_ vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__and2_1
XFILLER_21_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09178_ net475 _02870_ _04478_ _04804_ vssd1 vssd1 vccd1 vccd1 _05170_ sky130_fd_sc_hd__a31o_1
X_08129_ top.cb_syn.char_path_n\[105\] net378 net337 top.cb_syn.char_path_n\[103\]
+ net182 vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_112_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11140_ clknet_leaf_4_clk _01688_ _00495_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[42\]
+ sky130_fd_sc_hd__dfrtp_2
Xoutput45 net45 vssd1 vssd1 vccd1 vccd1 ADR_O[10] sky130_fd_sc_hd__buf_2
Xoutput67 net67 vssd1 vssd1 vccd1 vccd1 ADR_O[5] sky130_fd_sc_hd__buf_2
XANTENNA_fanout877_X net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput56 net56 vssd1 vssd1 vccd1 vccd1 ADR_O[21] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_112_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput89 net89 vssd1 vssd1 vccd1 vccd1 DAT_O[24] sky130_fd_sc_hd__buf_2
X_11071_ clknet_leaf_14_clk _01619_ _00426_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[101\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_8_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 DAT_O[14] sky130_fd_sc_hd__buf_2
X_10022_ net822 net662 vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__and2_1
XANTENNA__10968__Q top.cb_syn.char_index\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input16_A DAT_I[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11973_ top.translation.writeBin vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_113_Right_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10924_ clknet_leaf_34_clk _01479_ _00279_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.i\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08665__A top.cb_syn.h_element\[63\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06884__S net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07700__A2 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10855_ clknet_leaf_107_clk _01441_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_55_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05711__B2 top.WB.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10786_ clknet_leaf_76_clk _01385_ _00205_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11407_ clknet_leaf_99_clk _01955_ _00762_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[13\]
+ sky130_fd_sc_hd__dfstp_1
X_11338_ clknet_leaf_54_clk _01886_ _00693_ vssd1 vssd1 vccd1 vccd1 top.dut.out\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_74_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08177__C1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09943__B net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11269_ clknet_leaf_105_clk _01817_ _00624_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_05830_ _02835_ net290 top.sram_interface.write_counter_FLV\[0\] vssd1 vssd1 vccd1
+ vccd1 _02842_ sky130_fd_sc_hd__a21o_1
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10170__A net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07500_ top.cb_syn.char_path_n\[36\] top.cb_syn.char_path_n\[35\] top.cb_syn.char_path_n\[34\]
+ top.cb_syn.char_path_n\[33\] net399 net350 vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__mux4_1
X_05761_ top.compVal\[33\] net173 _02783_ top.WB.CPU_DAT_O\[1\] vssd1 vssd1 vccd1
+ vccd1 _02318_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_85_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08480_ net1131 top.cb_syn.char_path_n\[96\] net233 vssd1 vssd1 vccd1 vccd1 _01614_
+ sky130_fd_sc_hd__mux2_1
X_05692_ net22 net416 net308 top.WB.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 _02366_
+ sky130_fd_sc_hd__o22a_1
X_07431_ _04016_ _04027_ net354 vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__mux2_1
X_07362_ top.cw2\[7\] net135 _03547_ net119 net1694 vssd1 vssd1 vccd1 vccd1 _01895_
+ sky130_fd_sc_hd__a32o_1
XANTENNA__05702__B2 top.WB.CPU_DAT_O\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09101_ top.sram_interface.zero_cnt\[2\] _02449_ _02450_ _02763_ vssd1 vssd1 vccd1
+ vccd1 _05121_ sky130_fd_sc_hd__or4_1
X_06313_ top.hist_data_o\[5\] top.hist_data_o\[4\] vssd1 vssd1 vccd1 vccd1 _03176_
+ sky130_fd_sc_hd__and2_1
XFILLER_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07293_ _03795_ _03924_ _03805_ vssd1 vssd1 vccd1 vccd1 _03928_ sky130_fd_sc_hd__a21oi_1
X_06244_ _03109_ _02767_ _03012_ vssd1 vssd1 vccd1 vccd1 _03111_ sky130_fd_sc_hd__or3b_1
XANTENNA__08514__S net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09032_ net1251 top.WB.CPU_DAT_O\[25\] net292 vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__mux2_1
X_06175_ top.cw1\[6\] _02995_ vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__nor2_1
Xhold300 top.cb_syn.char_path\[33\] vssd1 vssd1 vccd1 vccd1 net1253 sky130_fd_sc_hd__dlygate4sd3_1
Xhold311 net77 vssd1 vssd1 vccd1 vccd1 net1264 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout203_A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold333 top.cb_syn.char_path\[47\] vssd1 vssd1 vccd1 vccd1 net1286 sky130_fd_sc_hd__dlygate4sd3_1
Xhold322 top.path\[115\] vssd1 vssd1 vccd1 vccd1 net1275 sky130_fd_sc_hd__dlygate4sd3_1
Xhold344 top.path\[91\] vssd1 vssd1 vccd1 vccd1 net1297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 net94 vssd1 vssd1 vccd1 vccd1 net1319 sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 top.cb_syn.char_path\[125\] vssd1 vssd1 vccd1 vccd1 net1330 sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 top.hTree.nulls\[55\] vssd1 vssd1 vccd1 vccd1 net1308 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout802 net806 vssd1 vssd1 vccd1 vccd1 net802 sky130_fd_sc_hd__buf_1
XFILLER_104_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09934_ net789 net629 vssd1 vssd1 vccd1 vccd1 _00548_ sky130_fd_sc_hd__and2_1
Xfanout824 net879 vssd1 vssd1 vccd1 vccd1 net824 sky130_fd_sc_hd__buf_2
Xhold388 top.path\[36\] vssd1 vssd1 vccd1 vccd1 net1341 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout813 net824 vssd1 vssd1 vccd1 vccd1 net813 sky130_fd_sc_hd__clkbuf_2
Xhold399 top.hTree.tree_reg\[42\] vssd1 vssd1 vccd1 vccd1 net1352 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout857 net878 vssd1 vssd1 vccd1 vccd1 net857 sky130_fd_sc_hd__clkbuf_2
X_09865_ net777 net617 vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__and2_1
Xfanout846 net849 vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input8_A DAT_I[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout835 net879 vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__clkbuf_2
Xfanout879 net34 vssd1 vssd1 vccd1 vccd1 net879 sky130_fd_sc_hd__clkbuf_4
Xfanout868 net877 vssd1 vssd1 vccd1 vccd1 net868 sky130_fd_sc_hd__buf_1
XANTENNA_fanout193_X net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07373__B net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08816_ top.path\[48\] top.path\[49\] top.path\[50\] top.path\[51\] net524 net523
+ vssd1 vssd1 vccd1 vccd1 _04999_ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout572_A net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06194__B2 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09796_ net774 net614 vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__and2_1
XANTENNA__09132__A1 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout458_X net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout360_X net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout837_A net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05959_ net452 top.translation.resEn net473 net36 vssd1 vssd1 vccd1 vccd1 _02897_
+ sky130_fd_sc_hd__or4b_1
XANTENNA_clkbuf_leaf_90_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08747_ net435 _04928_ _04929_ vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__o21a_1
X_08678_ _04878_ vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__inv_2
X_07629_ _04206_ _04207_ net487 vssd1 vssd1 vccd1 vccd1 _04208_ sky130_fd_sc_hd__mux2_1
XFILLER_53_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10640_ clknet_leaf_49_clk _00049_ _00059_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.word_cnt\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07531__A_N top.cb_syn.h_element\[54\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10571_ net810 net650 vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__and2_1
XFILLER_107_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05349__A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10255__A net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06957__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_11123_ clknet_leaf_25_clk _01671_ _00478_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_43_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08159__C1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11054_ clknet_leaf_20_clk _01602_ _00409_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[84\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08174__A2 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10005_ net820 net660 vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_58_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_101_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_10907_ clknet_leaf_31_clk top.header_synthesis.next_zero_count\[2\] _00262_ vssd1
+ vssd1 vccd1 vccd1 top.cb_syn.zero_count\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_72_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11887_ clknet_leaf_38_clk _02403_ _01242_ vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07685__B2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05696__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10838_ clknet_leaf_79_clk _01424_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_116_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10769_ clknet_leaf_43_clk _01368_ _00188_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[63\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_30_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08398__C1 _02504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07980_ top.cb_syn.zeroes\[2\] top.cb_syn.zero_count\[2\] vssd1 vssd1 vccd1 vccd1
+ _04483_ sky130_fd_sc_hd__xnor2_1
XFILLER_113_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06412__A2 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06931_ top.findLeastValue.val2\[18\] net146 net120 _03607_ vssd1 vssd1 vccd1 vccd1
+ _01960_ sky130_fd_sc_hd__o22a_1
XANTENNA__05620__B1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09650_ net781 net621 vssd1 vssd1 vccd1 vccd1 _00264_ sky130_fd_sc_hd__and2_1
X_08601_ _04821_ top.cb_syn.setup vssd1 vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__and2b_1
X_06862_ top.findLeastValue.startup _02773_ net288 vssd1 vssd1 vccd1 vccd1 _03576_
+ sky130_fd_sc_hd__nor3_2
XFILLER_67_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05813_ net1705 _02828_ _02830_ vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__o21ai_1
X_09581_ net793 net633 vssd1 vssd1 vccd1 vccd1 _00195_ sky130_fd_sc_hd__and2_1
X_06793_ top.findLeastValue.val1\[37\] net131 net115 top.compVal\[37\] vssd1 vssd1
+ vccd1 vccd1 _02045_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_38_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07480__Y _04071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05744_ _02775_ _02778_ vssd1 vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__nand2b_1
X_08532_ net1162 top.cb_syn.char_path_n\[44\] net220 vssd1 vssd1 vccd1 vccd1 _01562_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08463_ net1455 top.cb_syn.char_path_n\[113\] net222 vssd1 vssd1 vccd1 vccd1 _01631_
+ sky130_fd_sc_hd__mux2_1
X_07414_ net354 _04010_ _04011_ _04007_ _04012_ vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__a221o_1
X_05675_ top.hTree.node_reg\[33\] net311 _02750_ net480 vssd1 vssd1 vccd1 vccd1 _02751_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_18_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10059__B net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08394_ top.cb_syn.char_path_n\[5\] net391 _04752_ net509 net505 vssd1 vssd1 vccd1
+ vccd1 _04753_ sky130_fd_sc_hd__a221o_1
XANTENNA__08625__B1 _04826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout320_A _05088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07345_ net270 _03963_ _03964_ net275 net1687 vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__a32o_1
XANTENNA__09848__B net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_30_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_98_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout418_A _02758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07523__S1 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07276_ _03681_ _03911_ vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__xor2_1
X_06227_ top.cb_syn.char_index\[2\] top.cb_syn.char_index\[1\] vssd1 vssd1 vccd1 vccd1
+ _03095_ sky130_fd_sc_hd__or2_1
X_09015_ top.WB.CPU_DAT_O\[10\] net1223 net319 vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__mux2_1
Xhold152 top.header_synthesis.header\[3\] vssd1 vssd1 vccd1 vccd1 net1105 sky130_fd_sc_hd__dlygate4sd3_1
X_06158_ top.TRN_char_index\[5\] _02976_ vssd1 vssd1 vccd1 vccd1 _03029_ sky130_fd_sc_hd__nor2_1
Xhold130 top.cb_syn.char_path\[66\] vssd1 vssd1 vccd1 vccd1 net1083 sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 top.histogram.sram_out\[16\] vssd1 vssd1 vccd1 vccd1 net1094 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06939__B1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_05_915 vssd1 vssd1 vccd1 vccd1 team_05_915/HI gpio_out[30] sky130_fd_sc_hd__conb_1
Xteam_05_926 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] team_05_926/LO sky130_fd_sc_hd__conb_1
X_06089_ top.cb_syn.char_index\[4\] top.cb_syn.char_index\[3\] top.cb_syn.char_index\[2\]
+ top.cb_syn.char_index\[1\] vssd1 vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout787_A net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09583__B net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold163 top.hTree.finish_check vssd1 vssd1 vccd1 vccd1 net1116 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 top.histogram.sram_out\[20\] vssd1 vssd1 vccd1 vccd1 net1138 sky130_fd_sc_hd__dlygate4sd3_1
Xteam_05_904 vssd1 vssd1 vccd1 vccd1 team_05_904/HI gpio_out[19] sky130_fd_sc_hd__conb_1
Xhold174 top.path\[109\] vssd1 vssd1 vccd1 vccd1 net1127 sky130_fd_sc_hd__dlygate4sd3_1
Xteam_05_937 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] team_05_937/LO sky130_fd_sc_hd__conb_1
Xfanout621 net626 vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__buf_1
Xfanout610 net611 vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__clkbuf_2
Xfanout632 net646 vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__clkbuf_2
Xhold196 top.cb_syn.char_path\[1\] vssd1 vssd1 vccd1 vccd1 net1149 sky130_fd_sc_hd__dlygate4sd3_1
X_09917_ net742 net582 vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__and2_1
Xteam_05_948 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] team_05_948/LO sky130_fd_sc_hd__conb_1
XANTENNA__05611__B1 _02697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout643 net645 vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__clkbuf_2
XFILLER_98_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08156__A2 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout665 net675 vssd1 vssd1 vccd1 vccd1 net665 sky130_fd_sc_hd__clkbuf_2
Xfanout654 net657 vssd1 vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_97_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_97_clk sky130_fd_sc_hd__clkbuf_8
Xfanout676 net678 vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07364__B1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout687 net689 vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__clkbuf_2
Xfanout698 net699 vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__clkbuf_2
X_09848_ net744 net584 vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__and2_1
X_09779_ net765 net605 vssd1 vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__and2_1
XFILLER_18_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ clknet_leaf_90_clk _02327_ _01165_ vssd1 vssd1 vccd1 vccd1 top.compVal\[42\]
+ sky130_fd_sc_hd__dfrtp_2
X_11741_ clknet_leaf_59_clk _02274_ _01096_ vssd1 vssd1 vccd1 vccd1 top.histogram.init
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__08419__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11672_ clknet_leaf_43_clk _02205_ _01027_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10623_ net805 net645 vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_21_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07514__S1 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10554_ net828 net668 vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_58_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10485_ net831 net671 vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_118_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05850__B1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08395__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11106_ clknet_leaf_10_clk _01654_ _00461_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07294__A net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_88_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_88_clk sky130_fd_sc_hd__clkbuf_8
X_11037_ clknet_leaf_16_clk _01585_ _00392_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[67\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05669__B1 _02745_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05460_ _02417_ net466 vssd1 vssd1 vccd1 vccd1 _02568_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_15_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05391_ top.cb_syn.count\[7\] vssd1 vssd1 vccd1 vccd1 _02499_ sky130_fd_sc_hd__inv_2
XFILLER_20_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06881__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_12_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_8
X_07130_ _03786_ _03787_ vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__nand2_1
X_07061_ top.findLeastValue.val1\[12\] top.findLeastValue.val2\[12\] vssd1 vssd1 vccd1
+ vccd1 _03719_ sky130_fd_sc_hd__and2_1
XFILLER_114_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06012_ net1646 top.WB.CPU_DAT_O\[23\] net358 vssd1 vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__mux2_1
XANTENNA__05841__B1 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08386__A2 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07963_ net423 _04471_ _04470_ net287 vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_79_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_clk sky130_fd_sc_hd__clkbuf_8
X_09702_ net867 net707 vssd1 vssd1 vccd1 vccd1 _00316_ sky130_fd_sc_hd__and2_1
XFILLER_83_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06914_ top.compVal\[26\] top.findLeastValue.val1\[26\] net161 vssd1 vssd1 vccd1
+ vccd1 _03599_ sky130_fd_sc_hd__mux2_1
X_07894_ top.findLeastValue.sum\[9\] top.hTree.tree_reg\[9\] net283 vssd1 vssd1 vccd1
+ vccd1 _04421_ sky130_fd_sc_hd__mux2_1
XANTENNA__11227__Q top.cb_syn.end_cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06845_ top.findLeastValue.least1\[2\] net502 _03424_ vssd1 vssd1 vccd1 vccd1 _03562_
+ sky130_fd_sc_hd__mux2_1
X_09633_ net759 net599 vssd1 vssd1 vccd1 vccd1 _00247_ sky130_fd_sc_hd__and2_1
X_09564_ net795 net635 vssd1 vssd1 vccd1 vccd1 _00178_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout270_A net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08515_ net1400 top.cb_syn.char_path_n\[61\] net234 vssd1 vssd1 vccd1 vccd1 _01579_
+ sky130_fd_sc_hd__mux2_1
XFILLER_70_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06776_ top.findLeastValue.least1\[4\] net136 net118 net500 vssd1 vssd1 vccd1 vccd1
+ _02060_ sky130_fd_sc_hd__a22o_1
X_05727_ top.TRN_char_index\[0\] net38 net721 vssd1 vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__mux2_1
XFILLER_51_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09495_ net755 net595 vssd1 vssd1 vccd1 vccd1 _00109_ sky130_fd_sc_hd__and2_1
X_08446_ top.cb_syn.cb_enable _04800_ _04802_ _04804_ net1062 vssd1 vssd1 vccd1 vccd1
+ _01646_ sky130_fd_sc_hd__a41o_1
X_05658_ top.histogram.sram_out\[4\] net363 net419 top.hTree.node_reg\[4\] _02736_
+ vssd1 vssd1 vccd1 vccd1 _02737_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_102_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08377_ top.cb_syn.char_path_n\[109\] net391 _04735_ vssd1 vssd1 vccd1 vccd1 _04736_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_23_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05589_ _02677_ _02678_ net472 vssd1 vssd1 vccd1 vccd1 _02679_ sky130_fd_sc_hd__o21a_1
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07328_ _03721_ _03779_ _03776_ vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__or3b_1
XANTENNA_fanout323_X net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07259_ _03689_ _03690_ _03902_ vssd1 vssd1 vccd1 vccd1 _03903_ sky130_fd_sc_hd__or3b_1
XFILLER_3_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__09023__A0 top.WB.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10270_ net735 net575 vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__and2_1
XANTENNA__08377__A2 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07545__C _04134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout440 net442 vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__buf_2
Xfanout451 _02404_ vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__clkbuf_2
Xfanout462 top.controller.state_reg\[6\] vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__clkbuf_2
Xfanout484 net493 vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__clkbuf_2
Xfanout473 net477 vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__clkbuf_2
Xfanout495 top.histogram.init vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__buf_2
XFILLER_19_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07888__B2 top.findLeastValue.sum\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11724_ clknet_leaf_121_clk _02257_ _01079_ vssd1 vssd1 vccd1 vccd1 top.path\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06892__S net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11655_ clknet_leaf_110_clk _02188_ _01010_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08960__X _05087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07499__S0 _04072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11586_ clknet_leaf_15_clk _02134_ _00941_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10606_ net751 net591 vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_40_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10537_ net868 net708 vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__and2_1
XFILLER_50_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10468_ net729 net569 vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__and2_1
XANTENNA__09014__A0 top.WB.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10399_ net765 net605 vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_1_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_8
X_06630_ _03399_ _03400_ _03401_ vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_48_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06561_ _02432_ top.findLeastValue.val1\[17\] vssd1 vssd1 vccd1 vccd1 _03350_ sky130_fd_sc_hd__and2_1
XFILLER_18_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09280_ top.cb_syn.zero_count\[7\] _05227_ vssd1 vssd1 vccd1 vccd1 _05230_ sky130_fd_sc_hd__nor2_1
X_08300_ top.cb_syn.char_path_n\[19\] net198 _04677_ vssd1 vssd1 vccd1 vccd1 _01665_
+ sky130_fd_sc_hd__o21a_1
X_05512_ net462 top.hTree.node_reg\[60\] net362 net422 top.hTree.node_reg\[28\] vssd1
+ vssd1 vccd1 vccd1 _02615_ sky130_fd_sc_hd__a32o_1
X_06492_ _03286_ _03302_ vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__nor2_1
X_05443_ top.FLV_done _02548_ vssd1 vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__nand2_1
X_08231_ top.cb_syn.char_path_n\[54\] net384 net343 top.cb_syn.char_path_n\[52\] net188
+ vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__a221o_1
XANTENNA__06854__A2 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05374_ net504 vssd1 vssd1 vccd1 vccd1 _02482_ sky130_fd_sc_hd__inv_2
X_08162_ top.cb_syn.char_path_n\[88\] net208 _04608_ vssd1 vssd1 vccd1 vccd1 _01734_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__11510__Q top.findLeastValue.least1\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08093_ top.cb_syn.char_path_n\[123\] net385 net344 top.cb_syn.char_path_n\[121\]
+ net190 vssd1 vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__a221o_1
X_07113_ _03737_ _03738_ vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__and2b_1
XFILLER_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload50 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 clkload50/X sky130_fd_sc_hd__clkbuf_4
Xclkload61 clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 clkload61/Y sky130_fd_sc_hd__clkinv_1
XANTENNA__09005__A0 top.WB.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout116_A net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07044_ _03700_ _03701_ vssd1 vssd1 vccd1 vccd1 _03702_ sky130_fd_sc_hd__nand2_1
Xclkload72 clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 clkload72/X sky130_fd_sc_hd__clkbuf_8
Xclkload83 clknet_leaf_92_clk vssd1 vssd1 vccd1 vccd1 clkload83/Y sky130_fd_sc_hd__inv_4
Xclkload94 clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 clkload94/Y sky130_fd_sc_hd__inv_6
XANTENNA__07646__B _04221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_10_Left_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08764__C1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08995_ top.WB.CPU_DAT_O\[30\] net1082 net317 vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__mux2_1
XFILLER_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07946_ top.findLeastValue.least1\[6\] top.findLeastValue.least2\[6\] _04462_ vssd1
+ vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__mux2_1
XANTENNA__08758__A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05593__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07877_ net425 _04406_ _04407_ net258 vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__o211a_1
X_09616_ net801 net641 vssd1 vssd1 vccd1 vccd1 _00230_ sky130_fd_sc_hd__and2_1
X_06828_ top.findLeastValue.val1\[2\] net130 net114 net1712 vssd1 vssd1 vccd1 vccd1
+ _02010_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_104_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06759_ _03441_ _03546_ _03545_ vssd1 vssd1 vccd1 vccd1 _03547_ sky130_fd_sc_hd__or3b_4
X_09547_ net733 net573 vssd1 vssd1 vccd1 vccd1 _00161_ sky130_fd_sc_hd__and2_1
XANTENNA__09589__A net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09478_ net728 net568 vssd1 vssd1 vccd1 vccd1 _00092_ sky130_fd_sc_hd__and2_1
X_08429_ _02506_ top.cb_syn.char_path_n\[60\] _04787_ net511 vssd1 vssd1 vccd1 vccd1
+ _04788_ sky130_fd_sc_hd__o211a_1
XANTENNA__10528__A net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11440_ clknet_leaf_89_clk _01988_ _00795_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[46\]
+ sky130_fd_sc_hd__dfstp_1
Xclkload0 clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clkload0/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__06058__B1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11371_ clknet_leaf_102_clk _01919_ _00726_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[23\]
+ sky130_fd_sc_hd__dfrtp_2
X_10322_ net766 net606 vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_115_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10253_ net862 net702 vssd1 vssd1 vccd1 vccd1 _00867_ sky130_fd_sc_hd__and2_1
XFILLER_59_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10184_ net864 net704 vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__and2_1
XANTENNA__08755__C1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08668__A net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout281 net282 vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__clkbuf_2
Xfanout270 net272 vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__buf_2
Xfanout292 net294 vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06188__A top.cb_syn.char_index\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__09499__A net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11707_ clknet_leaf_114_clk _02240_ _01062_ vssd1 vssd1 vccd1 vccd1 top.path\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11638_ clknet_leaf_56_clk top.dut.bit_buf_next\[10\] _00993_ vssd1 vssd1 vccd1 vccd1
+ top.dut.bit_buf\[10\] sky130_fd_sc_hd__dfrtp_1
Xhold718 top.cb_syn.count\[5\] vssd1 vssd1 vccd1 vccd1 net1671 sky130_fd_sc_hd__dlygate4sd3_1
Xhold707 top.findLeastValue.wipe_the_char_1 vssd1 vssd1 vccd1 vccd1 net1660 sky130_fd_sc_hd__dlygate4sd3_1
X_11569_ clknet_leaf_107_clk _02117_ _00924_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_77_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold729 top.findLeastValue.sum\[12\] vssd1 vssd1 vccd1 vccd1 net1682 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10173__A net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_90_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08746__C1 _02523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07800_ top.hTree.tree_reg\[28\] top.findLeastValue.sum\[28\] net250 vssd1 vssd1
+ vccd1 vccd1 _04346_ sky130_fd_sc_hd__mux2_1
X_08780_ top.path\[126\] top.path\[127\] net526 vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__mux2_1
X_05992_ top.sram_interface.init_counter\[4\] _02913_ vssd1 vssd1 vccd1 vccd1 _02921_
+ sky130_fd_sc_hd__nor2_1
XFILLER_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06772__B2 _02767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05575__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07731_ net488 _04289_ vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__or2_1
X_07662_ top.findLeastValue.least1\[0\] top.hTree.tree_reg\[55\] net279 vssd1 vssd1
+ vccd1 vccd1 _04235_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07593_ top.cb_syn.max_index\[2\] top.cb_syn.max_index\[1\] vssd1 vssd1 vccd1 vccd1
+ _04179_ sky130_fd_sc_hd__xor2_1
X_09401_ top.hTree.nulls\[54\] _02809_ net240 _05277_ vssd1 vssd1 vccd1 vccd1 _05278_
+ sky130_fd_sc_hd__a211o_1
X_06613_ top.compVal\[37\] _02464_ vssd1 vssd1 vccd1 vccd1 _03402_ sky130_fd_sc_hd__or2_1
X_09332_ net972 net243 net218 _04458_ vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__a22o_1
X_06544_ net496 _02425_ top.compVal\[26\] _02472_ vssd1 vssd1 vccd1 vccd1 _03333_
+ sky130_fd_sc_hd__a2bb2o_1
X_09263_ _02532_ _05215_ vssd1 vssd1 vccd1 vccd1 _05218_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout233_A net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06475_ top.histogram.total\[28\] _03291_ net1552 vssd1 vssd1 vccd1 vccd1 _03296_
+ sky130_fd_sc_hd__a21oi_1
X_05426_ top.dut.out_valid vssd1 vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__inv_2
X_08214_ top.cb_syn.char_path_n\[62\] net209 _04634_ vssd1 vssd1 vccd1 vccd1 _01708_
+ sky130_fd_sc_hd__o21a_1
X_09194_ _02473_ _02799_ top.hTree.write_HT_fin vssd1 vssd1 vccd1 vccd1 _05177_ sky130_fd_sc_hd__o21a_1
X_08145_ top.cb_syn.char_path_n\[97\] net388 net347 top.cb_syn.char_path_n\[95\] net192
+ vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__a221o_1
X_05357_ top.findLeastValue.val1\[36\] vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout400_A net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08076_ net530 net538 vssd1 vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__nor2_1
XFILLER_115_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07027_ _03682_ _03683_ _03684_ vssd1 vssd1 vccd1 vccd1 _03685_ sky130_fd_sc_hd__or3_1
XFILLER_114_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold12 top.sram_interface.init_counter\[13\] vssd1 vssd1 vccd1 vccd1 net965 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout867_A net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout390_X net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold23 top.hTree.node_reg\[38\] vssd1 vssd1 vccd1 vccd1 net976 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 top.sram_interface.init_counter\[22\] vssd1 vssd1 vccd1 vccd1 net998 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_110_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold56 top.hTree.node_reg\[22\] vssd1 vssd1 vccd1 vccd1 net1009 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 top.hTree.node_reg\[18\] vssd1 vssd1 vccd1 vccd1 net987 sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ top.WB.CPU_DAT_O\[14\] net1152 net321 vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__mux2_1
Xhold89 net61 vssd1 vssd1 vccd1 vccd1 net1042 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 net57 vssd1 vssd1 vccd1 vccd1 net1031 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 top.hTree.tree_reg\[49\] vssd1 vssd1 vccd1 vccd1 net1020 sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ top.findLeastValue.sum\[2\] top.hTree.tree_reg\[2\] net282 vssd1 vssd1 vccd1
+ vccd1 _04449_ sky130_fd_sc_hd__mux2_1
X_10940_ clknet_leaf_34_clk _01495_ _00295_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.cb_length\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_56_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10871_ clknet_leaf_75_clk _01457_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout822_X net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09112__A net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06818__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_61_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11423_ clknet_leaf_82_clk _01971_ _00778_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[29\]
+ sky130_fd_sc_hd__dfstp_1
X_11354_ clknet_leaf_101_clk _01902_ _00709_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10305_ net799 net639 vssd1 vssd1 vccd1 vccd1 _00919_ sky130_fd_sc_hd__and2_1
X_11285_ clknet_leaf_80_clk net1576 _00640_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10236_ net842 net682 vssd1 vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__and2_1
XFILLER_67_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05557__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10167_ net840 net680 vssd1 vssd1 vccd1 vccd1 _00781_ sky130_fd_sc_hd__and2_1
XFILLER_47_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10098_ net827 net667 vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__and2_1
XFILLER_74_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06809__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06260_ _02508_ net561 _02577_ vssd1 vssd1 vccd1 vccd1 _03127_ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06191_ _02962_ _03060_ _02578_ vssd1 vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__and3b_1
Xhold515 top.histogram.sram_out\[25\] vssd1 vssd1 vccd1 vccd1 net1468 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05549__X _02646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold526 top.histogram.total\[7\] vssd1 vssd1 vccd1 vccd1 net1479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold504 top.cb_syn.char_path\[43\] vssd1 vssd1 vccd1 vccd1 net1457 sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 top.findLeastValue.histo_index\[1\] vssd1 vssd1 vccd1 vccd1 net1501 sky130_fd_sc_hd__dlygate4sd3_1
X_09950_ net738 net578 vssd1 vssd1 vccd1 vccd1 _00564_ sky130_fd_sc_hd__and2_1
Xhold537 top.histogram.total\[17\] vssd1 vssd1 vccd1 vccd1 net1490 sky130_fd_sc_hd__dlygate4sd3_1
Xhold559 top.path\[101\] vssd1 vssd1 vccd1 vccd1 net1512 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap289 net290 vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__clkbuf_1
X_08901_ _03325_ _05062_ _05064_ _04188_ vssd1 vssd1 vccd1 vccd1 _05071_ sky130_fd_sc_hd__o31ai_1
XANTENNA_clkbuf_4_9_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08800__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09881_ net736 net576 vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__and2_1
X_08832_ top.path\[32\] net410 _05014_ vssd1 vssd1 vccd1 vccd1 _05015_ sky130_fd_sc_hd__o21a_1
X_05975_ top.sram_interface.init_counter\[2\] top.sram_interface.init_counter\[1\]
+ top.sram_interface.init_counter\[0\] vssd1 vssd1 vccd1 vccd1 _02911_ sky130_fd_sc_hd__and3_1
XANTENNA__07643__C net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08763_ top.path\[90\] top.path\[91\] net526 vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout183_A net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07714_ top.findLeastValue.sum\[45\] top.hTree.tree_reg\[45\] net284 vssd1 vssd1
+ vccd1 vccd1 _04277_ sky130_fd_sc_hd__mux2_1
X_08694_ _04879_ _04885_ _04890_ _04875_ net1573 vssd1 vssd1 vccd1 vccd1 _01484_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_0_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout350_A net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07645_ top.findLeastValue.least1\[3\] _04199_ _04219_ vssd1 vssd1 vccd1 vccd1 _04221_
+ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_0_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10961__920 vssd1 vssd1 vccd1 vccd1 net920 _10961__920/LO sky130_fd_sc_hd__conb_1
X_07576_ net1549 _04164_ _04144_ vssd1 vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__mux2_1
XANTENNA__05720__A2 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06527_ top.dut.out\[0\] _03317_ vssd1 vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__nor2_1
XFILLER_80_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09315_ top.histogram.total\[24\] top.histogram.total\[25\] top.histogram.total\[26\]
+ top.histogram.total\[27\] net524 net523 vssd1 vssd1 vccd1 vccd1 _05250_ sky130_fd_sc_hd__mux4_1
X_09246_ top.header_synthesis.header\[4\] top.cb_syn.char_index\[4\] net518 vssd1
+ vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout615_A net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06458_ top.histogram.total\[8\] _03277_ _03278_ _03280_ vssd1 vssd1 vccd1 vccd1
+ _03281_ sky130_fd_sc_hd__and4_2
X_05409_ top.cb_syn.i\[6\] vssd1 vssd1 vccd1 vccd1 _02517_ sky130_fd_sc_hd__inv_2
X_09177_ top.cb_syn.curr_state\[5\] net475 _04862_ vssd1 vssd1 vccd1 vccd1 _05169_
+ sky130_fd_sc_hd__o21ba_1
X_06389_ net1231 _03230_ net300 vssd1 vssd1 vccd1 vccd1 _02125_ sky130_fd_sc_hd__mux2_1
X_08128_ top.cb_syn.char_path_n\[105\] net199 _04591_ vssd1 vssd1 vccd1 vccd1 _01751_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_112_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08059_ net505 net507 _04540_ net439 vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__o31a_1
Xoutput46 net46 vssd1 vssd1 vccd1 vccd1 ADR_O[11] sky130_fd_sc_hd__buf_2
Xoutput57 net57 vssd1 vssd1 vccd1 vccd1 ADR_O[22] sky130_fd_sc_hd__buf_2
X_11070_ clknet_leaf_14_clk _01618_ _00425_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[100\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 ADR_O[6] sky130_fd_sc_hd__buf_2
XANTENNA_fanout772_X net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10021_ net845 net685 vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__and2_1
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 DAT_O[15] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_8_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05539__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11972_ net453 vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09150__A2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05922__X _02892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_2_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10923_ clknet_leaf_34_clk _01478_ _00278_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.i\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10854_ clknet_leaf_77_clk _01440_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_55_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05711__A2 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10785_ clknet_leaf_47_clk _01384_ _00204_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[61\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08413__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11406_ clknet_leaf_99_clk _01954_ _00761_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[12\]
+ sky130_fd_sc_hd__dfstp_1
X_11337_ clknet_leaf_54_clk _01885_ _00692_ vssd1 vssd1 vccd1 vccd1 top.dut.out\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_74_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08177__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11268_ clknet_leaf_105_clk _01816_ _00623_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11199_ clknet_leaf_13_clk _01747_ _00554_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[101\]
+ sky130_fd_sc_hd__dfrtp_2
X_10219_ net808 net648 vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__and2_1
XANTENNA__07924__A0 top.findLeastValue.sum\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05760_ top.compVal\[34\] net173 net158 top.WB.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1
+ _02319_ sky130_fd_sc_hd__a22o_1
XANTENNA__10170__B net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05832__X _02843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05691_ net23 net415 net308 top.WB.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1 _02367_
+ sky130_fd_sc_hd__o22a_1
X_07430_ _04019_ _04026_ net404 vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_85_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05702__A2 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07361_ _03751_ net272 _03973_ net275 net1684 vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__a32o_1
X_09100_ net294 _02901_ _05118_ _05119_ vssd1 vssd1 vccd1 vccd1 _05120_ sky130_fd_sc_hd__or4_1
XANTENNA__08101__B1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06312_ top.hist_data_o\[4\] _03174_ vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__and2_1
X_09031_ net1089 top.WB.CPU_DAT_O\[26\] net292 vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__mux2_1
X_07292_ net269 _03926_ _03927_ net274 top.findLeastValue.sum\[23\] vssd1 vssd1 vccd1
+ vccd1 _01919_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_33_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06243_ _03109_ vssd1 vssd1 vccd1 vccd1 _03110_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06174_ net498 _02550_ _03005_ _03043_ vssd1 vssd1 vccd1 vccd1 _03044_ sky130_fd_sc_hd__o2bb2a_1
Xhold301 top.cb_syn.char_path\[87\] vssd1 vssd1 vccd1 vccd1 net1254 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08404__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05439__B net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold334 top.cb_syn.char_path\[32\] vssd1 vssd1 vccd1 vccd1 net1287 sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 top.cb_syn.char_path\[48\] vssd1 vssd1 vccd1 vccd1 net1276 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07000__A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold312 top.path\[51\] vssd1 vssd1 vccd1 vccd1 net1265 sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 net47 vssd1 vssd1 vccd1 vccd1 net1309 sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 top.cb_syn.char_path\[112\] vssd1 vssd1 vccd1 vccd1 net1331 sky130_fd_sc_hd__dlygate4sd3_1
Xhold345 top.path\[8\] vssd1 vssd1 vccd1 vccd1 net1298 sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 top.path\[127\] vssd1 vssd1 vccd1 vccd1 net1320 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout803 net805 vssd1 vssd1 vccd1 vccd1 net803 sky130_fd_sc_hd__clkbuf_2
XFILLER_98_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09933_ net791 net631 vssd1 vssd1 vccd1 vccd1 _00547_ sky130_fd_sc_hd__and2_1
Xhold389 top.path\[44\] vssd1 vssd1 vccd1 vccd1 net1342 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout825 net835 vssd1 vssd1 vccd1 vccd1 net825 sky130_fd_sc_hd__clkbuf_2
Xfanout814 net817 vssd1 vssd1 vccd1 vccd1 net814 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08530__S net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09864_ net770 net610 vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__and2_1
Xfanout847 net849 vssd1 vssd1 vccd1 vccd1 net847 sky130_fd_sc_hd__clkbuf_2
Xfanout858 net859 vssd1 vssd1 vccd1 vccd1 net858 sky130_fd_sc_hd__clkbuf_2
Xfanout836 net838 vssd1 vssd1 vccd1 vccd1 net836 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout869 net870 vssd1 vssd1 vccd1 vccd1 net869 sky130_fd_sc_hd__clkbuf_2
XFILLER_112_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__05455__A net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08815_ net432 _04996_ _04997_ vssd1 vssd1 vccd1 vccd1 _04998_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout186_X net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09795_ net774 net614 vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05958_ _02894_ _02895_ vssd1 vssd1 vccd1 vccd1 _02896_ sky130_fd_sc_hd__nor2_1
XFILLER_73_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08746_ top.path\[72\] net411 net329 top.path\[73\] _02523_ vssd1 vssd1 vccd1 vccd1
+ _04929_ sky130_fd_sc_hd__o221a_1
X_08677_ _02513_ _04877_ vssd1 vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout353_X net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05889_ top.cb_syn.h_element\[58\] top.cb_syn.h_element\[57\] top.cb_syn.h_element\[56\]
+ top.cb_syn.h_element\[55\] vssd1 vssd1 vccd1 vccd1 _02864_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout732_A net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05902__B _02875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07628_ top.findLeastValue.least1\[6\] _04206_ net394 vssd1 vssd1 vccd1 vccd1 _04207_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout520_X net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07559_ top.cb_syn.max_index\[6\] top.cb_syn.max_index\[5\] _04149_ vssd1 vssd1 vccd1
+ vccd1 _04150_ sky130_fd_sc_hd__or3_1
XFILLER_9_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10570_ net752 net592 vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__and2_1
X_09229_ _04485_ _05197_ vssd1 vssd1 vccd1 vccd1 _05198_ sky130_fd_sc_hd__and2b_1
XANTENNA__10255__B net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_2_Left_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_39_Left_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11122_ clknet_leaf_25_clk _01670_ _00477_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_88_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11053_ clknet_leaf_20_clk _01601_ _00408_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[83\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10004_ net818 net658 vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__and2_1
XFILLER_64_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05652__X _02732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_48_Left_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10906_ clknet_leaf_31_clk top.header_synthesis.next_zero_count\[1\] _00261_ vssd1
+ vssd1 vccd1 vccd1 top.cb_syn.zero_count\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_32_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11886_ clknet_leaf_54_clk _02402_ _01241_ vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__dfrtp_1
XANTENNA__05696__B2 top.WB.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06893__B1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10837_ clknet_leaf_76_clk _01423_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10768_ clknet_leaf_44_clk _01367_ _00187_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07842__C1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_57_Left_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10699_ clknet_leaf_111_clk _01298_ _00118_ vssd1 vssd1 vccd1 vccd1 top.path\[75\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08398__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06930_ top.compVal\[18\] top.findLeastValue.val1\[18\] net161 vssd1 vssd1 vccd1
+ vccd1 _03607_ sky130_fd_sc_hd__mux2_1
XANTENNA__10181__A net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10889__Q top.translation.index\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08600_ top.cb_syn.setup net475 _04820_ vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__and3_1
X_06861_ top.findLeastValue.histo_index\[7\] _03572_ _03568_ vssd1 vssd1 vccd1 vccd1
+ _03575_ sky130_fd_sc_hd__a21boi_1
X_05812_ net1622 _02829_ _02831_ vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_66_Left_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09580_ net793 net633 vssd1 vssd1 vccd1 vccd1 _00194_ sky130_fd_sc_hd__and2_1
X_06792_ top.findLeastValue.val1\[38\] net131 net115 top.compVal\[38\] vssd1 vssd1
+ vccd1 vccd1 _02046_ sky130_fd_sc_hd__o22a_1
X_05743_ _02548_ _02777_ vssd1 vssd1 vccd1 vccd1 _02778_ sky130_fd_sc_hd__nand2_1
XFILLER_35_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_38_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08531_ net1304 top.cb_syn.char_path_n\[45\] net224 vssd1 vssd1 vccd1 vccd1 _01563_
+ sky130_fd_sc_hd__mux2_1
X_05674_ _02748_ _02749_ vssd1 vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__or2_1
X_08462_ net1329 top.cb_syn.char_path_n\[114\] net222 vssd1 vssd1 vccd1 vccd1 _01632_
+ sky130_fd_sc_hd__mux2_1
X_07413_ top.dut.bits_in_buf\[1\] net404 _04003_ vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__and3_1
XANTENNA__07676__A2 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08393_ top.cb_syn.char_path_n\[7\] top.cb_syn.char_path_n\[8\] net513 vssd1 vssd1
+ vccd1 vccd1 _04752_ sky130_fd_sc_hd__mux2_1
X_07344_ _03769_ _03771_ vssd1 vssd1 vccd1 vccd1 _03964_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_98_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_75_Left_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07649__B net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07275_ net268 _03913_ _03914_ net273 net1680 vssd1 vssd1 vccd1 vccd1 _01923_ sky130_fd_sc_hd__a32o_1
X_06226_ _03091_ _03093_ net471 vssd1 vssd1 vccd1 vccd1 _03094_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout313_A net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09014_ top.WB.CPU_DAT_O\[11\] net1273 net319 vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__mux2_1
XFILLER_104_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06157_ top.cb_syn.max_index\[7\] _03025_ _03027_ top.hTree.nullSumIndex\[6\] vssd1
+ vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__a22o_1
Xhold120 top.hTree.nulls\[62\] vssd1 vssd1 vccd1 vccd1 net1073 sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 top.hTree.nulls\[46\] vssd1 vssd1 vccd1 vccd1 net1084 sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 net98 vssd1 vssd1 vccd1 vccd1 net1106 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09050__A1 top.WB.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold142 top.path\[76\] vssd1 vssd1 vccd1 vccd1 net1095 sky130_fd_sc_hd__dlygate4sd3_1
Xteam_05_905 vssd1 vssd1 vccd1 vccd1 team_05_905/HI gpio_out[20] sky130_fd_sc_hd__conb_1
X_06088_ top.cb_syn.char_index\[5\] top.cb_syn.char_index\[4\] _02958_ vssd1 vssd1
+ vccd1 vccd1 _02961_ sky130_fd_sc_hd__and3_1
Xteam_05_927 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] team_05_927/LO sky130_fd_sc_hd__conb_1
Xhold175 top.cb_syn.char_path\[67\] vssd1 vssd1 vccd1 vccd1 net1128 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout682_A net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_05_916 vssd1 vssd1 vccd1 vccd1 team_05_916/HI gpio_out[31] sky130_fd_sc_hd__conb_1
Xhold164 top.path\[96\] vssd1 vssd1 vccd1 vccd1 net1117 sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 top.histogram.sram_out\[11\] vssd1 vssd1 vccd1 vccd1 net1139 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout622 net626 vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__clkbuf_2
Xfanout611 net612 vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__clkbuf_2
Xteam_05_938 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] team_05_938/LO sky130_fd_sc_hd__conb_1
Xfanout633 net646 vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout600 net602 vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__clkbuf_2
X_09916_ net742 net582 vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__and2_1
Xteam_05_949 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] team_05_949/LO sky130_fd_sc_hd__conb_1
XANTENNA__05611__B2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold197 top.path\[14\] vssd1 vssd1 vccd1 vccd1 net1150 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout644 net645 vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__clkbuf_2
Xfanout655 net657 vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__buf_1
Xfanout666 net675 vssd1 vssd1 vccd1 vccd1 net666 sky130_fd_sc_hd__buf_1
XANTENNA_fanout470_X net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout688 net689 vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__buf_1
Xfanout699 net717 vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__clkbuf_2
Xfanout677 net678 vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__clkbuf_2
XFILLER_58_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_09847_ net743 net583 vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__and2_1
X_09778_ net792 net632 vssd1 vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__and2_1
XFILLER_37_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08729_ top.header_synthesis.write_num_lefts _03261_ vssd1 vssd1 vccd1 vccd1 _04913_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_107_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ clknet_leaf_66_clk _02273_ _01095_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.zero_cnt\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07667__A2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11671_ clknet_leaf_43_clk _02204_ _01026_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06875__B1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10622_ net805 net645 vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__and2_1
X_10553_ net834 net674 vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__and2_1
XFILLER_108_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_58_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10484_ net831 net671 vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_118_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08919__A2 _04188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05850__B2 top.WB.CPU_DAT_O\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09041__A1 top.WB.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09143__C_N _05088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11105_ clknet_leaf_9_clk _01653_ _00460_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11036_ clknet_leaf_17_clk _01584_ _00391_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[66\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07355__B2 top.findLeastValue.sum\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05669__B2 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11869_ clknet_leaf_7_clk _02385_ _01224_ vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05390_ net534 vssd1 vssd1 vccd1 vccd1 _02498_ sky130_fd_sc_hd__inv_2
XANTENNA__06094__A1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07060_ _03716_ _03717_ vssd1 vssd1 vccd1 vccd1 _03718_ sky130_fd_sc_hd__nor2_1
X_06011_ net1605 top.WB.CPU_DAT_O\[24\] net358 vssd1 vssd1 vccd1 vccd1 _02199_ sky130_fd_sc_hd__mux2_1
XANTENNA__09032__A1 top.WB.CPU_DAT_O\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05841__B2 top.WB.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06397__A2 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09701_ net869 net709 vssd1 vssd1 vccd1 vccd1 _00315_ sky130_fd_sc_hd__and2_1
X_07962_ net414 _02770_ vssd1 vssd1 vccd1 vccd1 _04471_ sky130_fd_sc_hd__nor2_1
XFILLER_114_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11508__Q top.findLeastValue.least1\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06913_ top.findLeastValue.val2\[27\] net147 net121 _03598_ vssd1 vssd1 vccd1 vccd1
+ _01969_ sky130_fd_sc_hd__o22a_1
X_07893_ net440 net1443 net251 top.findLeastValue.sum\[10\] _04420_ vssd1 vssd1 vccd1
+ vccd1 _01815_ sky130_fd_sc_hd__a221o_1
XANTENNA__09335__A2 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06844_ _02477_ net152 net126 _03561_ vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__a2bb2o_1
X_09632_ net759 net599 vssd1 vssd1 vccd1 vccd1 _00246_ sky130_fd_sc_hd__and2_1
X_09563_ net795 net635 vssd1 vssd1 vccd1 vccd1 _00177_ sky130_fd_sc_hd__and2_1
X_08514_ net1271 top.cb_syn.char_path_n\[62\] net235 vssd1 vssd1 vccd1 vccd1 _01580_
+ sky130_fd_sc_hd__mux2_1
X_06775_ top.findLeastValue.least1\[5\] net136 net118 net498 vssd1 vssd1 vccd1 vccd1
+ _02061_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout263_A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05726_ top.TRN_char_index\[1\] net39 net720 vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__mux2_1
XFILLER_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09494_ net755 net595 vssd1 vssd1 vccd1 vccd1 _00108_ sky130_fd_sc_hd__and2_1
X_08445_ top.cb_syn.end_check top.cb_syn.curr_state\[5\] net474 vssd1 vssd1 vccd1
+ vccd1 _04804_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_42_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05657_ top.hTree.node_reg\[36\] net310 _02735_ net480 vssd1 vssd1 vccd1 vccd1 _02736_
+ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_83_Left_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08376_ top.cb_syn.char_path_n\[110\] net330 _04734_ net510 net438 vssd1 vssd1 vccd1
+ vccd1 _04735_ sky130_fd_sc_hd__a221o_1
X_05588_ top.cb_syn.char_path\[15\] net557 net312 top.cb_syn.char_path\[111\] vssd1
+ vssd1 vccd1 vccd1 _02678_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout149_X net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout528_A top.translation.index\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07327_ net269 _03951_ _03952_ net274 net1702 vssd1 vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__a32o_1
XFILLER_99_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout316_X net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_57_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07258_ _03697_ _03700_ _03900_ _03698_ _03694_ vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__a311o_1
X_06209_ net561 _02959_ _03077_ _02557_ top.cb_syn.curr_index\[5\] vssd1 vssd1 vccd1
+ vccd1 _03078_ sky130_fd_sc_hd__a32o_1
XANTENNA_clkbuf_leaf_100_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07189_ top.findLeastValue.val1\[43\] top.findLeastValue.val2\[43\] vssd1 vssd1 vccd1
+ vccd1 _03847_ sky130_fd_sc_hd__nand2_1
XFILLER_105_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_EDGE_ROW_92_Left_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout685_X net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout430 _02535_ vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__buf_2
XANTENNA__05596__B1 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout441 net442 vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__clkbuf_4
Xfanout463 net465 vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__buf_2
Xfanout474 net477 vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__clkbuf_4
Xfanout452 net455 vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_115_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout485 net487 vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__buf_2
Xfanout496 top.findLeastValue.val1\[25\] vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__buf_2
XANTENNA__05899__A1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08837__A1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06848__B1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11723_ clknet_leaf_122_clk _02256_ _01078_ vssd1 vssd1 vccd1 vccd1 top.path\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11654_ clknet_leaf_110_clk _02187_ _01009_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10605_ net751 net591 vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_12_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07499__S1 _04071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11585_ clknet_leaf_14_clk _02133_ _00940_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_40_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10536_ net868 net708 vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_108_Right_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10467_ net729 net569 vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__and2_1
XANTENNA__07544__A_N _04134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10398_ net765 net605 vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__and2_1
XANTENNA__06413__S net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05587__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11019_ clknet_leaf_21_clk _01567_ _00374_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_52_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06560_ _02431_ top.findLeastValue.val1\[18\] vssd1 vssd1 vccd1 vccd1 _03349_ sky130_fd_sc_hd__and2_1
XFILLER_33_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05511_ _02612_ _02613_ net476 vssd1 vssd1 vccd1 vccd1 _02614_ sky130_fd_sc_hd__o21a_1
XFILLER_60_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06491_ net1567 _03285_ vssd1 vssd1 vccd1 vccd1 _03302_ sky130_fd_sc_hd__nor2_1
X_05442_ net451 net541 vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__and2_1
X_08230_ top.cb_syn.char_path_n\[54\] net205 _04642_ vssd1 vssd1 vccd1 vccd1 _01700_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__05511__B1 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08161_ top.cb_syn.char_path_n\[89\] net387 net346 top.cb_syn.char_path_n\[87\] net191
+ vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__a221o_1
X_05373_ top.findLeastValue.histo_index\[7\] vssd1 vssd1 vccd1 vccd1 _02481_ sky130_fd_sc_hd__inv_2
X_08092_ top.cb_syn.char_path_n\[123\] net206 _04573_ vssd1 vssd1 vccd1 vccd1 _01769_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__08803__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07112_ top.findLeastValue.val1\[6\] top.findLeastValue.val2\[6\] _03738_ _03737_
+ vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__a31oi_2
Xclkload51 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 clkload51/Y sky130_fd_sc_hd__clkinv_2
Xclkload62 clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 clkload62/Y sky130_fd_sc_hd__clkinv_1
Xclkload40 clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 clkload40/X sky130_fd_sc_hd__clkbuf_8
X_07043_ top.findLeastValue.val1\[28\] top.findLeastValue.val2\[28\] vssd1 vssd1 vccd1
+ vccd1 _03701_ sky130_fd_sc_hd__or2_1
Xclkload84 clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 clkload84/Y sky130_fd_sc_hd__clkinv_4
Xclkload73 clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 clkload73/Y sky130_fd_sc_hd__inv_6
Xclkload95 clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 clkload95/X sky130_fd_sc_hd__clkbuf_8
X_08994_ top.WB.CPU_DAT_O\[31\] net1182 net317 vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__mux2_1
XFILLER_102_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07945_ top.hTree.state\[6\] top.hTree.state\[3\] vssd1 vssd1 vccd1 vccd1 _04462_
+ sky130_fd_sc_hd__or2_2
XANTENNA_fanout380_A net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06790__A2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09615_ net798 net638 vssd1 vssd1 vccd1 vccd1 _00229_ sky130_fd_sc_hd__and2_1
X_07876_ net482 _04405_ vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout645_A net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout266_X net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06827_ top.findLeastValue.val1\[3\] net130 net114 top.compVal\[3\] vssd1 vssd1 vccd1
+ vccd1 _02011_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_104_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09546_ net733 net573 vssd1 vssd1 vccd1 vccd1 _00160_ sky130_fd_sc_hd__and2_1
X_06758_ _03457_ _03544_ _03445_ _03455_ vssd1 vssd1 vccd1 vccd1 _03546_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09589__B net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09477_ net728 net568 vssd1 vssd1 vccd1 vccd1 _00091_ sky130_fd_sc_hd__and2_1
X_05709_ net4 net416 net309 top.WB.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1 _02349_
+ sky130_fd_sc_hd__o22a_1
X_08428_ net515 top.cb_syn.char_path_n\[59\] vssd1 vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__or2_1
X_06689_ _02435_ top.findLeastValue.val2\[14\] _03475_ _03476_ vssd1 vssd1 vccd1 vccd1
+ _03477_ sky130_fd_sc_hd__a211o_1
XFILLER_24_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10528__B net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08359_ _02504_ _04701_ _04704_ _04717_ vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__o31a_1
Xclkload1 clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clkload1/X sky130_fd_sc_hd__clkbuf_8
X_11370_ clknet_leaf_102_clk _01918_ _00725_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10321_ net764 net604 vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__and2_1
XFILLER_118_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10252_ net862 net702 vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__and2_1
XANTENNA__08755__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10183_ net865 net705 vssd1 vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__and2_1
XANTENNA__05569__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input39_A gpio_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout282 _04198_ vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__buf_2
XANTENNA__05584__A3 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout271 net272 vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__buf_2
Xfanout260 net261 vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__buf_2
Xfanout293 net294 vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__clkbuf_4
XFILLER_75_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11706_ clknet_leaf_116_clk _02239_ _01061_ vssd1 vssd1 vccd1 vccd1 top.path\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11637_ clknet_leaf_56_clk top.dut.bit_buf_next\[9\] _00992_ vssd1 vssd1 vccd1 vccd1
+ top.dut.bit_buf\[9\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__07246__B1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11568_ clknet_leaf_102_clk _02116_ _00923_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_116_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10519_ net856 net696 vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__and2_1
Xhold708 top.findLeastValue.sum\[26\] vssd1 vssd1 vccd1 vccd1 net1661 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07797__A1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold719 top.histogram.total\[15\] vssd1 vssd1 vccd1 vccd1 net1672 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06454__D1 top.controller.state_reg\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08994__A0 top.WB.CPU_DAT_O\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11499_ clknet_leaf_91_clk _02047_ _00854_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[39\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_97_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_90_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10173__B net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08746__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05991_ _02907_ _02920_ vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__nor2_1
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06772__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07730_ top.findLeastValue.sum\[42\] _04289_ net398 vssd1 vssd1 vccd1 vccd1 _04290_
+ sky130_fd_sc_hd__mux2_1
X_07661_ top.hTree.tree_reg\[55\] net394 net286 vssd1 vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__and3_1
XFILLER_92_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07592_ net532 top.cb_syn.h_element\[47\] net539 top.cb_syn.h_element\[56\] _04135_
+ vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__a221o_1
X_09400_ top.findLeastValue.least2\[8\] net394 net248 top.hTree.tree_reg\[54\] net406
+ vssd1 vssd1 vccd1 vccd1 _05277_ sky130_fd_sc_hd__o221a_1
XFILLER_18_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06612_ _02409_ top.findLeastValue.val1\[41\] _02462_ top.compVal\[40\] vssd1 vssd1
+ vccd1 vccd1 _03401_ sky130_fd_sc_hd__a2bb2o_1
X_09331_ _02809_ net241 vssd1 vssd1 vccd1 vccd1 _05262_ sky130_fd_sc_hd__nor2_1
X_06543_ _02425_ net496 top.findLeastValue.val1\[24\] vssd1 vssd1 vccd1 vccd1 _03332_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_4_5_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09262_ _02532_ _05215_ vssd1 vssd1 vccd1 vccd1 _05217_ sky130_fd_sc_hd__or2_1
X_06474_ _03293_ _03295_ vssd1 vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__and2_1
X_05425_ top.cb_syn.zero_count\[5\] vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__inv_2
XANTENNA__09226__A1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08213_ top.cb_syn.char_path_n\[63\] net388 net347 top.cb_syn.char_path_n\[61\] net192
+ vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__a221o_1
X_09193_ top.hTree.wait_cnt top.hTree.state\[2\] net264 _05100_ top.hTree.state\[6\]
+ vssd1 vssd1 vccd1 vccd1 _00024_ sky130_fd_sc_hd__a32o_1
X_08144_ top.cb_syn.char_path_n\[97\] net209 _04599_ vssd1 vssd1 vccd1 vccd1 _01743_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__08434__C1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout226_A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05356_ top.findLeastValue.val1\[37\] vssd1 vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__inv_2
XANTENNA__08985__A0 top.WB.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08075_ _04557_ _04558_ _04561_ _04559_ vssd1 vssd1 vccd1 vccd1 _04562_ sky130_fd_sc_hd__or4b_2
X_07026_ top.findLeastValue.val1\[24\] top.findLeastValue.val2\[24\] vssd1 vssd1 vccd1
+ vccd1 _03684_ sky130_fd_sc_hd__xnor2_1
Xhold13 top.hTree.node_reg\[61\] vssd1 vssd1 vccd1 vccd1 net966 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_110_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold24 top.hTree.node_reg\[52\] vssd1 vssd1 vccd1 vccd1 net977 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 top.hTree.node_reg\[51\] vssd1 vssd1 vccd1 vccd1 net988 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05566__A3 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout762_A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold46 top.hTree.node_reg\[3\] vssd1 vssd1 vccd1 vccd1 net999 sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ top.WB.CPU_DAT_O\[15\] net1112 net321 vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_110_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold68 top.hTree.tree_reg\[51\] vssd1 vssd1 vccd1 vccd1 net1021 sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 top.hTree.node_reg\[27\] vssd1 vssd1 vccd1 vccd1 net1010 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 top.hTree.node_reg\[2\] vssd1 vssd1 vccd1 vccd1 net1032 sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ net444 net1387 net255 top.findLeastValue.sum\[3\] _04448_ vssd1 vssd1 vccd1
+ vccd1 _01808_ sky130_fd_sc_hd__a221o_1
XFILLER_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07859_ top.findLeastValue.sum\[16\] top.hTree.tree_reg\[16\] net284 vssd1 vssd1
+ vccd1 vccd1 _04393_ sky130_fd_sc_hd__mux2_1
XFILLER_44_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10870_ clknet_leaf_76_clk _01456_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_3_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09529_ net749 net589 vssd1 vssd1 vccd1 vccd1 _00143_ sky130_fd_sc_hd__and2_1
XANTENNA__06279__A1 top.cb_syn.char_index\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09112__B net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08425__C1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11422_ clknet_leaf_97_clk _01970_ _00777_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[28\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__08976__A0 top.WB.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11353_ clknet_leaf_91_clk _01901_ _00708_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_10304_ net798 net638 vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__and2_1
X_11284_ clknet_leaf_79_clk net1556 _00639_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10235_ net840 net680 vssd1 vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__and2_1
XANTENNA__06898__S net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10166_ net827 net667 vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__and2_1
XANTENNA__05962__B1 top.TRN_sram_complete vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10097_ net828 net668 vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__and2_1
XANTENNA_clkload4_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07703__B2 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05714__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10999_ clknet_leaf_28_clk _01547_ _00354_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_06190_ top.cb_syn.char_index\[3\] top.cb_syn.char_index\[2\] top.cb_syn.char_index\[1\]
+ top.cb_syn.char_index\[4\] vssd1 vssd1 vccd1 vccd1 _03060_ sky130_fd_sc_hd__a31o_1
XANTENNA__08967__A0 top.WB.CPU_DAT_O\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08431__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold505 top.hTree.node_reg\[31\] vssd1 vssd1 vccd1 vccd1 net1458 sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 top.histogram.total\[27\] vssd1 vssd1 vccd1 vccd1 net1469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold527 top.histogram.total\[10\] vssd1 vssd1 vccd1 vccd1 net1480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 top.hist_data_o\[31\] vssd1 vssd1 vccd1 vccd1 net1491 sky130_fd_sc_hd__dlygate4sd3_1
Xhold549 top.hTree.state\[7\] vssd1 vssd1 vccd1 vccd1 net1502 sky130_fd_sc_hd__dlygate4sd3_1
X_08900_ _04151_ _04187_ _05069_ vssd1 vssd1 vccd1 vccd1 _05070_ sky130_fd_sc_hd__a21o_1
X_09880_ net758 net598 vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__and2_1
X_08831_ top.path\[33\] net328 _05013_ net434 net437 vssd1 vssd1 vccd1 vccd1 _05014_
+ sky130_fd_sc_hd__o221a_1
XANTENNA__05548__A3 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05974_ top.sram_interface.init_counter\[1\] top.sram_interface.init_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02910_ sky130_fd_sc_hd__and2_1
XANTENNA__05953__A0 top.WB.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08762_ top.path\[100\] net410 net328 top.path\[101\] net522 vssd1 vssd1 vccd1 vccd1
+ _04945_ sky130_fd_sc_hd__o221a_1
X_08693_ _02513_ _04877_ vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__nand2_1
X_07713_ net445 net1520 net262 _04276_ vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout176_A _02589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07644_ top.findLeastValue.least1\[3\] top.hTree.tree_reg\[58\] net281 vssd1 vssd1
+ vccd1 vccd1 _04220_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07575_ top.cb_syn.max_index\[5\] _04136_ _04161_ _04163_ vssd1 vssd1 vccd1 vccd1
+ _04164_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout343_A net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06526_ top.dut.out\[7\] top.dut.out\[6\] top.dut.out\[5\] top.dut.out\[4\] vssd1
+ vssd1 vccd1 vccd1 _03317_ sky130_fd_sc_hd__or4b_1
XANTENNA__05460__B net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09314_ _05246_ _05247_ _05248_ net521 vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__a22o_1
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09245_ net1054 _05207_ net296 vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_header\[3\]
+ sky130_fd_sc_hd__mux2_1
X_06457_ top.histogram.total\[11\] top.histogram.total\[10\] top.histogram.total\[9\]
+ vssd1 vssd1 vccd1 vccd1 _03280_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout131_X net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05408_ top.cb_syn.zeroes\[0\] vssd1 vssd1 vccd1 vccd1 _02516_ sky130_fd_sc_hd__inv_2
X_09176_ _04867_ _05168_ vssd1 vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__or2_1
XANTENNA__08958__A0 top.WB.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06388_ _03180_ _03229_ vssd1 vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__nor2_1
X_08127_ top.cb_syn.char_path_n\[106\] net374 net334 top.cb_syn.char_path_n\[104\]
+ net179 vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__a221o_1
X_05339_ top.compVal\[2\] vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__inv_2
X_08058_ net507 net246 _04540_ vssd1 vssd1 vccd1 vccd1 _04549_ sky130_fd_sc_hd__or3_1
XANTENNA__07630__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput47 net47 vssd1 vssd1 vccd1 vccd1 ADR_O[12] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_112_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput58 net58 vssd1 vssd1 vccd1 vccd1 ADR_O[23] sky130_fd_sc_hd__buf_2
X_07009_ top.findLeastValue.val1\[37\] top.findLeastValue.val2\[37\] vssd1 vssd1 vccd1
+ vccd1 _03667_ sky130_fd_sc_hd__nor2_1
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 ADR_O[7] sky130_fd_sc_hd__buf_2
XANTENNA__05916__A _02760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10020_ net819 net659 vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_8_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07933__B2 top.findLeastValue.sum\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05944__A0 top.WB.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11971_ net453 vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__clkbuf_1
XFILLER_17_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_10922_ clknet_leaf_34_clk _01477_ _00277_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_27_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10853_ clknet_leaf_107_clk _01439_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[45\]
+ sky130_fd_sc_hd__dfxtp_1
X_10784_ clknet_leaf_76_clk _01383_ _00203_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[60\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05801__D net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08949__A0 top.WB.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11405_ clknet_leaf_96_clk _01953_ _00760_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[11\]
+ sky130_fd_sc_hd__dfstp_2
X_11336_ clknet_leaf_54_clk _01884_ _00691_ vssd1 vssd1 vccd1 vccd1 top.dut.out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_74_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11267_ clknet_leaf_105_clk _01815_ _00622_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_79_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_11198_ clknet_leaf_16_clk _01746_ _00553_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[100\]
+ sky130_fd_sc_hd__dfrtp_2
X_10218_ net814 net654 vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__and2_1
X_10149_ net814 net654 vssd1 vssd1 vccd1 vccd1 _00763_ sky130_fd_sc_hd__and2_1
XANTENNA__05935__A0 top.WB.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05959__D_N net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05690_ net25 net418 net360 top.WB.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1 _02368_
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10179__A net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07360_ top.findLeastValue.val1\[0\] top.findLeastValue.val2\[0\] vssd1 vssd1 vccd1
+ vccd1 _03973_ sky130_fd_sc_hd__or2_1
XANTENNA__09320__X _05255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06311_ top.hist_data_o\[3\] top.hist_data_o\[2\] top.hist_data_o\[1\] top.hist_data_o\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__and4_1
X_09030_ net1167 top.WB.CPU_DAT_O\[27\] net292 vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__mux2_1
X_07291_ _03803_ _03925_ _03802_ vssd1 vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__a21bo_1
X_06242_ top.findLeastValue.histo_index\[3\] net502 net503 net504 vssd1 vssd1 vccd1
+ vccd1 _03109_ sky130_fd_sc_hd__and4_1
X_06173_ top.cw2\[6\] _03003_ _02572_ vssd1 vssd1 vccd1 vccd1 _03043_ sky130_fd_sc_hd__o21ai_1
Xhold302 top.cb_syn.char_path\[57\] vssd1 vssd1 vccd1 vccd1 net1255 sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 top.cb_syn.char_path\[91\] vssd1 vssd1 vccd1 vccd1 net1288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold313 top.cb_syn.char_path\[97\] vssd1 vssd1 vccd1 vccd1 net1266 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07000__B _03657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07775__X _04326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold324 top.path\[9\] vssd1 vssd1 vccd1 vccd1 net1277 sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 top.cb_syn.char_path\[122\] vssd1 vssd1 vccd1 vccd1 net1299 sky130_fd_sc_hd__dlygate4sd3_1
X_09932_ net790 net630 vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__and2_1
Xhold357 top.hTree.tree_reg\[56\] vssd1 vssd1 vccd1 vccd1 net1310 sky130_fd_sc_hd__dlygate4sd3_1
Xhold368 top.path\[123\] vssd1 vssd1 vccd1 vccd1 net1321 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout804 net805 vssd1 vssd1 vccd1 vccd1 net804 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09365__B1 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout815 net817 vssd1 vssd1 vccd1 vccd1 net815 sky130_fd_sc_hd__buf_1
Xhold379 top.path\[121\] vssd1 vssd1 vccd1 vccd1 net1332 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09208__A net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout848 net849 vssd1 vssd1 vccd1 vccd1 net848 sky130_fd_sc_hd__buf_1
X_09863_ net770 net610 vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__and2_1
Xfanout837 net838 vssd1 vssd1 vccd1 vccd1 net837 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout293_A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout826 net835 vssd1 vssd1 vccd1 vccd1 net826 sky130_fd_sc_hd__buf_1
XANTENNA__07915__A1 top.findLeastValue.sum\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout859 net877 vssd1 vssd1 vccd1 vccd1 net859 sky130_fd_sc_hd__clkbuf_2
X_09794_ net774 net614 vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__and2_1
X_08814_ top.path\[52\] net408 net326 top.path\[53\] net521 vssd1 vssd1 vccd1 vccd1
+ _04997_ sky130_fd_sc_hd__o221a_1
XANTENNA__05926__A0 top.WB.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08745_ top.path\[74\] top.path\[75\] net527 vssd1 vssd1 vccd1 vccd1 _04928_ sky130_fd_sc_hd__mux2_1
X_05957_ net556 net465 vssd1 vssd1 vccd1 vccd1 _02895_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout558_A net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08676_ _02514_ _04876_ vssd1 vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__or2_1
X_05888_ _02554_ _02858_ _02861_ vssd1 vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__and3_1
XFILLER_26_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07627_ top.findLeastValue.least1\[6\] top.hTree.tree_reg\[61\] net285 vssd1 vssd1
+ vccd1 vccd1 _04206_ sky130_fd_sc_hd__mux2_1
X_07558_ top.cb_syn.max_index\[4\] _04148_ vssd1 vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_52_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07526__S0 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06509_ top.histogram.total\[8\] _03279_ net1647 vssd1 vssd1 vccd1 vccd1 _03310_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout513_X net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07489_ top.cb_syn.char_path_n\[4\] top.cb_syn.char_path_n\[3\] top.cb_syn.char_path_n\[2\]
+ net517 net399 net350 vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__mux4_1
X_09228_ _02514_ top.cb_syn.zero_count\[2\] _04491_ _05196_ _04487_ vssd1 vssd1 vccd1
+ vccd1 _05197_ sky130_fd_sc_hd__a311o_1
X_09159_ net962 net1515 net265 vssd1 vssd1 vccd1 vccd1 _00018_ sky130_fd_sc_hd__mux2_1
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_11121_ clknet_leaf_24_clk _01669_ _00476_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06957__A2 net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11052_ clknet_leaf_21_clk _01600_ _00407_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[82\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_103_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10003_ net818 net658 vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__and2_1
XFILLER_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input21_A DAT_I[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_13_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_103_Left_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11885_ clknet_leaf_38_clk _02401_ _01240_ vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__dfrtp_1
X_10905_ clknet_leaf_31_clk top.header_synthesis.next_zero_count\[0\] _00260_ vssd1
+ vssd1 vccd1 vccd1 top.cb_syn.zero_count\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA__08331__B2 top.cb_syn.char_path_n\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10836_ clknet_leaf_80_clk _01422_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05696__A2 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07800__S net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10767_ clknet_leaf_44_clk _01366_ _00186_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[61\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10698_ clknet_leaf_111_clk _01297_ _00117_ vssd1 vssd1 vccd1 vccd1 top.path\[74\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_112_Left_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11319_ clknet_leaf_76_clk _01867_ _00674_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10181__B net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09347__B1 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06860_ net500 _03109_ _03573_ vssd1 vssd1 vccd1 vccd1 _03574_ sky130_fd_sc_hd__and3_1
X_05811_ top.sram_interface.counter_HTREE\[3\] _02829_ _02830_ vssd1 vssd1 vccd1 vccd1
+ _02831_ sky130_fd_sc_hd__a21boi_1
XFILLER_95_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06791_ top.findLeastValue.val1\[39\] net131 net115 net1719 vssd1 vssd1 vccd1 vccd1
+ _02047_ sky130_fd_sc_hd__o22a_1
XFILLER_36_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05742_ _02776_ vssd1 vssd1 vccd1 vccd1 _02777_ sky130_fd_sc_hd__inv_2
X_08530_ net1419 top.cb_syn.char_path_n\[46\] net221 vssd1 vssd1 vccd1 vccd1 _01564_
+ sky130_fd_sc_hd__mux2_1
XFILLER_36_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05673_ top.cb_syn.char_path\[1\] net560 net315 top.cb_syn.char_path\[97\] vssd1
+ vssd1 vccd1 vccd1 _02749_ sky130_fd_sc_hd__a22o_1
X_08461_ net1389 top.cb_syn.char_path_n\[115\] net222 vssd1 vssd1 vccd1 vccd1 _01633_
+ sky130_fd_sc_hd__mux2_1
X_07412_ net354 net404 vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__nor2_1
XFILLER_50_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07508__S0 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08392_ net510 _04749_ _04750_ vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__a21o_1
XFILLER_50_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07343_ _03769_ _03771_ vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout139_A net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07649__C net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07833__B1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07274_ _03679_ _03912_ _03678_ vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__a21bo_1
X_06225_ _03040_ _03089_ _03092_ _02574_ vssd1 vssd1 vccd1 vccd1 _03093_ sky130_fd_sc_hd__a2bb2o_1
X_09013_ top.WB.CPU_DAT_O\[12\] net1095 net319 vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__mux2_1
Xhold110 _01646_ vssd1 vssd1 vccd1 vccd1 net1063 sky130_fd_sc_hd__dlygate4sd3_1
X_06156_ top.sram_interface.word_cnt\[13\] net541 _03026_ vssd1 vssd1 vccd1 vccd1
+ _03027_ sky130_fd_sc_hd__or3_2
Xhold121 net86 vssd1 vssd1 vccd1 vccd1 net1074 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08541__S net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold132 top.cb_syn.char_path\[39\] vssd1 vssd1 vccd1 vccd1 net1085 sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 top.path\[12\] vssd1 vssd1 vccd1 vccd1 net1096 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_1_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_05_906 vssd1 vssd1 vccd1 vccd1 team_05_906/HI gpio_out[21] sky130_fd_sc_hd__conb_1
X_06087_ top.cb_syn.char_index\[4\] top.cb_syn.char_index\[3\] _02957_ vssd1 vssd1
+ vccd1 vccd1 _02960_ sky130_fd_sc_hd__and3_1
Xhold165 top.path\[48\] vssd1 vssd1 vccd1 vccd1 net1118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 net103 vssd1 vssd1 vccd1 vccd1 net1129 sky130_fd_sc_hd__dlygate4sd3_1
Xteam_05_917 vssd1 vssd1 vccd1 vccd1 team_05_917/HI gpio_out[32] sky130_fd_sc_hd__conb_1
Xhold154 top.path\[92\] vssd1 vssd1 vccd1 vccd1 net1107 sky130_fd_sc_hd__dlygate4sd3_1
Xteam_05_939 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] team_05_939/LO sky130_fd_sc_hd__conb_1
Xfanout623 net626 vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__buf_1
Xfanout612 net647 vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__clkbuf_2
Xhold187 top.cb_syn.char_path\[119\] vssd1 vssd1 vccd1 vccd1 net1140 sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 top.histogram.sram_out\[23\] vssd1 vssd1 vccd1 vccd1 net1151 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout601 net602 vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__buf_1
XANTENNA__05611__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_05_928 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] team_05_928/LO sky130_fd_sc_hd__conb_1
X_09915_ net741 net581 vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__and2_1
Xfanout645 net646 vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__clkbuf_2
Xfanout634 net636 vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__clkbuf_2
X_09846_ net742 net582 vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout675_A net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout656 net657 vssd1 vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__clkbuf_2
Xfanout667 net669 vssd1 vssd1 vccd1 vccd1 net667 sky130_fd_sc_hd__clkbuf_2
Xfanout689 net718 vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__clkbuf_2
Xfanout678 net719 vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__dlymetal6s2s_1
X_09777_ net788 net628 vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout842_A net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06989_ top.findLeastValue.val1\[42\] top.findLeastValue.val1\[41\] top.findLeastValue.val1\[40\]
+ top.findLeastValue.val1\[39\] vssd1 vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__and4_1
X_08728_ top.cb_syn.num_lefts\[4\] top.cb_syn.num_lefts\[3\] top.cb_syn.num_lefts\[2\]
+ top.cb_syn.num_lefts\[1\] top.header_synthesis.count\[0\] top.header_synthesis.count\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_107_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08659_ net529 _04137_ _04529_ _04862_ _02872_ vssd1 vssd1 vccd1 vccd1 _04863_ sky130_fd_sc_hd__o2111a_1
XFILLER_54_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11670_ clknet_leaf_43_clk _02203_ _01025_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10621_ net769 net609 vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__and2_1
XANTENNA__07824__A0 top.findLeastValue.sum\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10552_ net829 net669 vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__and2_1
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10483_ net831 net671 vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_118_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08451__S net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05850__A2 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09329__B1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11104_ clknet_leaf_9_clk _01652_ _00459_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_77_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11035_ clknet_leaf_17_clk _01583_ _00390_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[65\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08687__A _04875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06759__X _03547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08599__A_N top.CB_write_complete vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05669__A2 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08855__A2 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06866__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11868_ clknet_leaf_115_clk _02384_ _01223_ vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__dfrtp_1
XFILLER_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11799_ clknet_leaf_108_clk _02316_ _01154_ vssd1 vssd1 vccd1 vccd1 top.translation.write_fin
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10819_ clknet_leaf_105_clk _01405_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_06010_ net1626 top.WB.CPU_DAT_O\[25\] net357 vssd1 vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__mux2_1
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_114_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__05841__A2 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07961_ top.findLeastValue.alternator_timer\[2\] top.findLeastValue.alternator_timer\[1\]
+ top.findLeastValue.alternator_timer\[0\] _03566_ top.findLeastValue.alternator_timer\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04470_ sky130_fd_sc_hd__a41o_1
XFILLER_101_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09700_ net867 net707 vssd1 vssd1 vccd1 vccd1 _00314_ sky130_fd_sc_hd__and2_1
X_06912_ top.compVal\[27\] top.findLeastValue.val1\[27\] net162 vssd1 vssd1 vccd1
+ vccd1 _03598_ sky130_fd_sc_hd__mux2_1
XFILLER_68_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05573__X _02666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07892_ net425 _04418_ _04419_ net258 vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__o211a_1
X_06843_ top.findLeastValue.least1\[3\] top.findLeastValue.histo_index\[3\] _03424_
+ vssd1 vssd1 vccd1 vccd1 _03561_ sky130_fd_sc_hd__mux2_1
X_09631_ net759 net599 vssd1 vssd1 vccd1 vccd1 _00245_ sky130_fd_sc_hd__and2_1
X_09562_ net795 net635 vssd1 vssd1 vccd1 vccd1 _00176_ sky130_fd_sc_hd__and2_1
X_06774_ top.findLeastValue.least1\[6\] net136 net118 net497 vssd1 vssd1 vccd1 vccd1
+ _02062_ sky130_fd_sc_hd__a22o_1
X_05725_ top.TRN_char_index\[2\] net40 net720 vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__mux2_1
XANTENNA__09099__A2 _02843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08513_ net1154 top.cb_syn.char_path_n\[63\] net233 vssd1 vssd1 vccd1 vccd1 _01581_
+ sky130_fd_sc_hd__mux2_1
X_09493_ net756 net596 vssd1 vssd1 vccd1 vccd1 _00107_ sky130_fd_sc_hd__and2_1
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08444_ top.cb_syn.cb_enable _04802_ vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__nand2_1
X_05656_ _02733_ _02734_ vssd1 vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__or2_1
XANTENNA__08059__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout423_A net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08375_ top.cb_syn.char_path_n\[111\] top.cb_syn.char_path_n\[112\] net514 vssd1
+ vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__mux2_1
X_05587_ top.cb_syn.char_path\[79\] net551 net542 top.cb_syn.char_path\[47\] vssd1
+ vssd1 vccd1 vccd1 _02677_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_102_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07326_ _03718_ _03950_ vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout211_X net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout309_X net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07257_ _03697_ _03700_ _03900_ _03698_ vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__a31o_1
X_06208_ top.cb_syn.char_index\[3\] _02957_ vssd1 vssd1 vccd1 vccd1 _03077_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout792_A net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07188_ _03842_ _03845_ vssd1 vssd1 vccd1 vccd1 _03846_ sky130_fd_sc_hd__nand2b_1
XFILLER_105_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_105_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_06139_ top.cw1\[7\] _02996_ vssd1 vssd1 vccd1 vccd1 _03010_ sky130_fd_sc_hd__xor2_1
Xfanout420 net421 vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout431 _02530_ vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06793__B1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout453 net455 vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__clkbuf_4
Xfanout475 net477 vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__buf_1
Xfanout464 net465 vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__buf_1
Xfanout442 net448 vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__buf_2
XANTENNA__08534__A1 top.cb_syn.char_path_n\[42\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout845_X net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout497 top.findLeastValue.histo_index\[6\] vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__buf_2
X_09829_ net768 net608 vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__and2_1
Xfanout486 net487 vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__buf_2
XFILLER_58_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11722_ clknet_leaf_122_clk _02255_ _01077_ vssd1 vssd1 vccd1 vccd1 top.path\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11653_ clknet_leaf_109_clk _02186_ _01008_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05520__B2 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10604_ net752 net592 vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_12_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11584_ clknet_leaf_14_clk _02132_ _00939_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_40_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10535_ net867 net707 vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__and2_1
X_10466_ net730 net570 vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__and2_1
XANTENNA__05658__X _02737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10397_ net763 net603 vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__and2_1
XANTENNA__08773__A1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06784__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11018_ clknet_leaf_7_clk _01566_ _00373_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_49_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05510_ top.cb_syn.char_path\[28\] net559 net314 top.cb_syn.char_path\[124\] vssd1
+ vssd1 vccd1 vccd1 _02613_ sky130_fd_sc_hd__a22o_1
XANTENNA__06839__A1 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06490_ net1494 _03286_ vssd1 vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__xor2_1
X_05441_ _02536_ _02548_ vssd1 vssd1 vccd1 vccd1 _02549_ sky130_fd_sc_hd__nor2_1
X_08160_ top.cb_syn.char_path_n\[89\] net208 _04607_ vssd1 vssd1 vccd1 vccd1 _01735_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__08880__A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05372_ top.findLeastValue.histo_index\[8\] vssd1 vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__inv_2
X_07111_ _03741_ _03768_ _03739_ vssd1 vssd1 vccd1 vccd1 _03769_ sky130_fd_sc_hd__o21ai_1
X_08091_ top.cb_syn.char_path_n\[124\] net385 net344 top.cb_syn.char_path_n\[122\]
+ net189 vssd1 vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__a221o_1
Xclkload52 clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 clkload52/X sky130_fd_sc_hd__clkbuf_8
Xclkload30 clknet_leaf_112_clk vssd1 vssd1 vccd1 vccd1 clkload30/X sky130_fd_sc_hd__clkbuf_4
Xclkload41 clknet_leaf_109_clk vssd1 vssd1 vccd1 vccd1 clkload41/X sky130_fd_sc_hd__clkbuf_4
X_07042_ top.findLeastValue.val1\[28\] top.findLeastValue.val2\[28\] vssd1 vssd1 vccd1
+ vccd1 _03700_ sky130_fd_sc_hd__nand2_1
Xclkload63 clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 clkload63/Y sky130_fd_sc_hd__bufinv_16
Xclkload96 clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 clkload96/Y sky130_fd_sc_hd__clkinv_4
Xclkload85 clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 clkload85/X sky130_fd_sc_hd__clkbuf_8
Xclkload74 clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 clkload74/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_87_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08993_ top.sram_interface.TRN_counter\[0\] _02889_ _02890_ vssd1 vssd1 vccd1 vccd1
+ _05088_ sky130_fd_sc_hd__or3b_4
XANTENNA__06775__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_1_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07944_ top.hTree.state\[6\] top.hTree.state\[9\] top.hTree.state\[3\] top.hTree.state\[4\]
+ net264 vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__o41a_4
X_07875_ top.hTree.tree_reg\[13\] top.findLeastValue.sum\[13\] net247 vssd1 vssd1
+ vccd1 vccd1 _04406_ sky130_fd_sc_hd__mux2_1
X_09614_ net797 net637 vssd1 vssd1 vccd1 vccd1 _00228_ sky130_fd_sc_hd__and2_1
X_06826_ top.findLeastValue.val1\[4\] net130 net114 top.compVal\[4\] vssd1 vssd1 vccd1
+ vccd1 _02012_ sky130_fd_sc_hd__o22a_1
XFILLER_71_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08819__A2 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09545_ net733 net573 vssd1 vssd1 vccd1 vccd1 _00159_ sky130_fd_sc_hd__and2_1
XANTENNA__05750__B2 top.WB.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout161_X net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06757_ _03521_ _03525_ _03539_ _03457_ vssd1 vssd1 vccd1 vccd1 _03545_ sky130_fd_sc_hd__a211o_1
XFILLER_36_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout259_X net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06688_ top.compVal\[15\] _02493_ vssd1 vssd1 vccd1 vccd1 _03476_ sky130_fd_sc_hd__nor2_1
X_05708_ net5 net416 net309 top.WB.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1 _02350_
+ sky130_fd_sc_hd__o22a_1
X_09476_ net732 net572 vssd1 vssd1 vccd1 vccd1 _00090_ sky130_fd_sc_hd__and2_1
X_08427_ top.cb_syn.char_path_n\[61\] top.cb_syn.char_path_n\[62\] top.cb_syn.char_path_n\[63\]
+ top.cb_syn.char_path_n\[64\] net516 net512 vssd1 vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__mux4_1
X_05639_ top.hTree.node_reg\[39\] net310 _02720_ net480 vssd1 vssd1 vccd1 vccd1 _02721_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__05502__B2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout805_A net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09886__A net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09101__D _02763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08358_ net506 _04714_ _04716_ top.cb_syn.end_cnt\[4\] vssd1 vssd1 vccd1 vccd1 _04717_
+ sky130_fd_sc_hd__o31a_1
Xclkload2 clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clkload2/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__06058__A2 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08289_ top.cb_syn.char_path_n\[25\] net383 net344 top.cb_syn.char_path_n\[23\] net187
+ vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__a221o_1
X_07309_ net1648 net273 net268 _03939_ vssd1 vssd1 vccd1 vccd1 _01914_ sky130_fd_sc_hd__a22o_1
XFILLER_109_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10320_ net764 net604 vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_115_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10251_ net866 net706 vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__and2_1
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10182_ net865 net705 vssd1 vssd1 vccd1 vccd1 _00796_ sky130_fd_sc_hd__and2_1
XANTENNA__07963__C1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout250 _04199_ vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__clkbuf_4
XFILLER_115_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout272 _03864_ vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__buf_2
Xfanout261 net267 vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__buf_2
Xfanout283 net284 vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__clkbuf_4
Xfanout294 _02896_ vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_66_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08684__B _04134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07494__A1 _04084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11705_ clknet_leaf_116_clk _02238_ _01060_ vssd1 vssd1 vccd1 vccd1 top.path\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11636_ clknet_leaf_55_clk top.dut.bit_buf_next\[8\] _00991_ vssd1 vssd1 vccd1 vccd1
+ top.dut.bit_buf\[8\] sky130_fd_sc_hd__dfrtp_1
X_11567_ clknet_leaf_106_clk _02115_ _00922_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10518_ net855 net695 vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__and2_1
Xhold709 top.findLeastValue.sum\[30\] vssd1 vssd1 vccd1 vccd1 net1662 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_77_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11498_ clknet_leaf_92_clk _02046_ _00853_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[38\]
+ sky130_fd_sc_hd__dfstp_2
X_10449_ net753 net593 vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__and2_1
XFILLER_111_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05990_ top.sram_interface.init_counter\[5\] _02906_ vssd1 vssd1 vccd1 vccd1 _02920_
+ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_41_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09171__A1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_56_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07660_ net263 _04232_ _04233_ net1310 net446 vssd1 vssd1 vccd1 vccd1 _01861_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_88_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07591_ top.cb_syn.h_element\[56\] top.cb_syn.h_element\[47\] _04145_ vssd1 vssd1
+ vccd1 vccd1 _04177_ sky130_fd_sc_hd__mux2_1
XFILLER_80_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06611_ top.compVal\[42\] _02461_ _03397_ _03398_ vssd1 vssd1 vccd1 vccd1 _03400_
+ sky130_fd_sc_hd__o211a_1
X_09330_ net486 _02809_ net262 _00053_ vssd1 vssd1 vccd1 vccd1 _05261_ sky130_fd_sc_hd__o211ai_2
X_06542_ top.compVal\[28\] _02470_ _02471_ net494 vssd1 vssd1 vccd1 vccd1 _03331_
+ sky130_fd_sc_hd__a22o_1
X_09261_ _05213_ _05215_ _05216_ _05214_ top.cb_syn.zero_count\[1\] vssd1 vssd1 vccd1
+ vccd1 top.header_synthesis.next_zero_count\[1\] sky130_fd_sc_hd__a32o_1
XFILLER_33_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05496__B1 _02601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08212_ top.cb_syn.char_path_n\[63\] net209 _04633_ vssd1 vssd1 vccd1 vccd1 _01709_
+ sky130_fd_sc_hd__o21a_1
X_06473_ top.histogram.total\[30\] _03292_ vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__or2_1
X_05424_ top.cb_syn.zero_count\[2\] vssd1 vssd1 vccd1 vccd1 _02532_ sky130_fd_sc_hd__inv_2
X_09192_ top.controller.fin_reg\[6\] net1589 _05176_ vssd1 vssd1 vccd1 vccd1 _00013_
+ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_114_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08143_ top.cb_syn.char_path_n\[98\] net388 net346 top.cb_syn.char_path_n\[96\] net191
+ vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout121_A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05355_ top.findLeastValue.val1\[38\] vssd1 vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__inv_2
X_08074_ _02497_ _04480_ _04560_ vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__a21o_1
XANTENNA__05739__A net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07025_ net496 top.findLeastValue.val2\[25\] vssd1 vssd1 vccd1 vccd1 _03683_ sky130_fd_sc_hd__xnor2_1
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold14 top.hTree.node_reg\[62\] vssd1 vssd1 vccd1 vccd1 net967 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout588_A net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold36 top.sram_interface.init_counter\[21\] vssd1 vssd1 vccd1 vccd1 net989 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_110_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xhold25 top.hTree.node_reg\[58\] vssd1 vssd1 vccd1 vccd1 net978 sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ top.WB.CPU_DAT_O\[16\] net1386 net323 vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__mux2_1
Xhold47 top.hTree.node_reg\[1\] vssd1 vssd1 vccd1 vccd1 net1000 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_110_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09162__A1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold69 top.hTree.tree_reg\[52\] vssd1 vssd1 vccd1 vccd1 net1022 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 top.hTree.node_reg\[19\] vssd1 vssd1 vccd1 vccd1 net1011 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout755_A net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07927_ net429 _04446_ _04447_ net260 vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__o211a_1
X_07858_ net441 net1450 net253 top.findLeastValue.sum\[17\] _04392_ vssd1 vssd1 vccd1
+ vccd1 _01822_ sky130_fd_sc_hd__a221o_1
XANTENNA__08370__C1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout543_X net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07789_ top.findLeastValue.sum\[30\] top.hTree.tree_reg\[30\] net285 vssd1 vssd1
+ vccd1 vccd1 _04337_ sky130_fd_sc_hd__mux2_1
XFILLER_44_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06809_ top.findLeastValue.val1\[21\] net128 net112 top.compVal\[21\] vssd1 vssd1
+ vccd1 vccd1 _02029_ sky130_fd_sc_hd__o22a_1
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09528_ net755 net595 vssd1 vssd1 vccd1 vccd1 _00142_ sky130_fd_sc_hd__and2_1
XFILLER_12_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09459_ net869 net709 vssd1 vssd1 vccd1 vccd1 _00073_ sky130_fd_sc_hd__and2_1
XFILLER_101_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07688__X _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11421_ clknet_leaf_98_clk _01969_ _00776_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[27\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11352_ clknet_leaf_91_clk _01900_ _00707_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_10303_ net798 net638 vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__and2_1
X_11283_ clknet_leaf_79_clk net1460 _00638_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10234_ net840 net680 vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__and2_1
X_10165_ net821 net661 vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_72_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10096_ net828 net668 vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__and2_1
XFILLER_74_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08361__C1 _02504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05714__B2 top.WB.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06911__B1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10998_ clknet_leaf_29_clk _01546_ _00353_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11619_ clknet_leaf_67_clk _02167_ _00974_ vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__dfrtp_1
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold517 top.hTree.nullSumIndex\[0\] vssd1 vssd1 vccd1 vccd1 net1470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold506 top.hTree.tree_reg\[26\] vssd1 vssd1 vccd1 vccd1 net1459 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xhold539 top.histogram.total\[11\] vssd1 vssd1 vccd1 vccd1 net1492 sky130_fd_sc_hd__dlygate4sd3_1
Xhold528 top.hist_data_o\[11\] vssd1 vssd1 vccd1 vccd1 net1481 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08830_ top.path\[34\] top.path\[35\] net528 vssd1 vssd1 vccd1 vccd1 _05013_ sky130_fd_sc_hd__mux2_1
X_05973_ top.sram_interface.init_counter\[9\] top.sram_interface.init_counter\[8\]
+ _02908_ vssd1 vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__and3_1
XANTENNA__09144__A1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08761_ net435 _04943_ vssd1 vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__or2_1
X_08692_ _04880_ _04885_ _04889_ _04875_ top.cb_syn.zeroes\[4\] vssd1 vssd1 vccd1
+ vccd1 _01485_ sky130_fd_sc_hd__a32o_1
X_07712_ _04274_ _04275_ net487 vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__mux2_1
X_07643_ top.hTree.tree_reg\[58\] net398 net286 vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__and3_1
XANTENNA__08352__C1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05705__B2 top.WB.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout169_A _02845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07574_ net537 _04160_ _04162_ net531 vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__a22o_1
X_09313_ top.histogram.total\[20\] top.histogram.total\[21\] top.histogram.total\[22\]
+ top.histogram.total\[23\] net524 net523 vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__mux4_1
X_06525_ top.histogram.eof_n top.histogram.state\[0\] vssd1 vssd1 vccd1 vccd1 _03316_
+ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout336_A net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_60_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_clk sky130_fd_sc_hd__clkbuf_8
X_09244_ top.header_synthesis.header\[3\] top.cb_syn.char_index\[3\] net518 vssd1
+ vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__mux2_1
XANTENNA__08544__S net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06456_ _03277_ _03278_ vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__and2_1
X_05407_ top.cb_syn.zeroes\[1\] vssd1 vssd1 vccd1 vccd1 _02515_ sky130_fd_sc_hd__inv_2
X_09175_ net536 _05096_ _05167_ _02930_ vssd1 vssd1 vccd1 vccd1 _05168_ sky130_fd_sc_hd__a22o_1
X_08126_ top.cb_syn.char_path_n\[106\] net196 _04590_ vssd1 vssd1 vccd1 vccd1 _01752_
+ sky130_fd_sc_hd__o21a_1
X_06387_ top.hist_data_o\[9\] _03179_ top.hist_data_o\[10\] vssd1 vssd1 vccd1 vccd1
+ _03229_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout124_X net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05338_ top.compVal\[3\] vssd1 vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__inv_2
X_08057_ top.cb_syn.end_cnt\[4\] _04548_ _04545_ vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput48 net48 vssd1 vssd1 vccd1 vccd1 ADR_O[13] sky130_fd_sc_hd__buf_2
X_07008_ _03665_ vssd1 vssd1 vccd1 vccd1 _03666_ sky130_fd_sc_hd__inv_2
Xoutput59 net59 vssd1 vssd1 vccd1 vccd1 ADR_O[24] sky130_fd_sc_hd__buf_2
XANTENNA__05475__Y _02583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout493_X net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08186__A2 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08959_ top.WB.CPU_DAT_O\[14\] top.cb_syn.h_element\[46\] net369 vssd1 vssd1 vccd1
+ vccd1 _01351_ sky130_fd_sc_hd__mux2_1
X_11970_ net453 vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__clkbuf_1
X_10921_ clknet_leaf_34_clk _01476_ _00276_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07697__B2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10852_ clknet_leaf_108_clk _01438_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[44\]
+ sky130_fd_sc_hd__dfxtp_1
X_10783_ clknet_leaf_77_clk _01382_ _00202_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[59\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_51_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08454__S net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06763__A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11404_ clknet_leaf_96_clk _01952_ _00759_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[10\]
+ sky130_fd_sc_hd__dfstp_1
X_11335_ clknet_leaf_54_clk _01883_ _00690_ vssd1 vssd1 vccd1 vccd1 top.dut.out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_74_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11266_ clknet_leaf_105_clk _01814_ _00621_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_79_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08177__A2 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10217_ net810 net650 vssd1 vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__and2_1
XFILLER_79_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11197_ clknet_leaf_16_clk _01745_ _00552_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[99\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09374__B2 _04290_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06003__A net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10148_ net814 net654 vssd1 vssd1 vccd1 vccd1 _00762_ sky130_fd_sc_hd__and2_1
XFILLER_39_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10079_ net852 net692 vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__and2_1
XANTENNA__09126__A1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05699__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11352__Q top.findLeastValue.sum\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xclkbuf_leaf_42_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_clk sky130_fd_sc_hd__clkbuf_8
X_07290_ _03802_ _03803_ _03925_ vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__nand3b_1
X_06310_ top.hist_data_o\[1\] top.hist_data_o\[0\] vssd1 vssd1 vccd1 vccd1 _03173_
+ sky130_fd_sc_hd__nand2_1
X_06241_ net1413 net141 _03108_ net160 vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__a22o_1
X_06172_ _03040_ _03041_ _03039_ vssd1 vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__or3b_1
Xhold314 top.cb_syn.char_path\[117\] vssd1 vssd1 vccd1 vccd1 net1267 sky130_fd_sc_hd__dlygate4sd3_1
Xhold325 top.hTree.closing vssd1 vssd1 vccd1 vccd1 net1278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold303 top.cb_syn.char_path\[37\] vssd1 vssd1 vccd1 vccd1 net1256 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09931_ net776 net616 vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__and2_1
Xhold347 top.cb_syn.char_path\[54\] vssd1 vssd1 vccd1 vccd1 net1300 sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 top.cb_syn.char_path\[34\] vssd1 vssd1 vccd1 vccd1 net1322 sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 top.path\[50\] vssd1 vssd1 vccd1 vccd1 net1311 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05623__B1 _02707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold336 top.path\[98\] vssd1 vssd1 vccd1 vccd1 net1289 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout805 net806 vssd1 vssd1 vccd1 vccd1 net805 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08168__A2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout816 net817 vssd1 vssd1 vccd1 vccd1 net816 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07376__B1 _03553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout849 net878 vssd1 vssd1 vccd1 vccd1 net849 sky130_fd_sc_hd__clkbuf_2
X_09862_ net770 net610 vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__and2_1
Xfanout838 net879 vssd1 vssd1 vccd1 vccd1 net838 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09365__B2 _04326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout827 net829 vssd1 vssd1 vccd1 vccd1 net827 sky130_fd_sc_hd__clkbuf_2
X_09793_ net774 net614 vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__and2_1
X_08813_ top.path\[54\] top.path\[55\] net525 vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__mux2_1
XFILLER_85_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_05956_ net452 _02891_ vssd1 vssd1 vccd1 vccd1 _02894_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout286_A _04197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08744_ top.path\[76\] top.path\[77\] top.path\[78\] top.path\[79\] net527 net523
+ vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout453_A net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08675_ top.cb_syn.zeroes\[1\] top.cb_syn.zeroes\[0\] vssd1 vssd1 vccd1 vccd1 _04876_
+ sky130_fd_sc_hd__nand2_1
X_05887_ _02858_ _02861_ vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__and2_1
XANTENNA__07679__B2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07626_ net458 net1453 net257 _04205_ vssd1 vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__o22a_1
XFILLER_14_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout620_A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07557_ top.cb_syn.max_index\[3\] top.cb_syn.max_index\[2\] top.cb_syn.max_index\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__or3_1
XFILLER_81_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_33_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout718_A net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09212__D_N top.controller.fin_reg\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07526__S1 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06508_ net1480 _03308_ vssd1 vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__xor2_1
X_07488_ _04075_ _04076_ _04077_ _04078_ _04072_ _04071_ vssd1 vssd1 vccd1 vccd1 _04079_
+ sky130_fd_sc_hd__mux4_1
X_06439_ top.header_synthesis.count\[2\] _03256_ _03263_ vssd1 vssd1 vccd1 vccd1 _03265_
+ sky130_fd_sc_hd__o21ai_1
X_09227_ _04486_ _04490_ _04492_ vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_32_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09158_ top.hTree.wait_cnt net1535 net264 _05100_ top.hTree.state\[9\] vssd1 vssd1
+ vccd1 vccd1 _00027_ sky130_fd_sc_hd__a32o_1
X_09089_ net1545 _05108_ _05109_ _02581_ vssd1 vssd1 vccd1 vccd1 _00037_ sky130_fd_sc_hd__a211o_1
X_08109_ top.cb_syn.char_path_n\[115\] net375 net335 top.cb_syn.char_path_n\[113\]
+ net180 vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__a221o_1
X_11120_ clknet_leaf_25_clk _01668_ _00475_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[22\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__05614__B1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07367__B1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09118__B net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11051_ clknet_leaf_21_clk _01599_ _00406_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[81\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10002_ net818 net658 vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__and2_1
XFILLER_57_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11814__D net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input14_A DAT_I[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11884_ clknet_leaf_39_clk _02400_ _01239_ vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__dfrtp_1
X_10904_ clknet_leaf_38_clk top.header_synthesis.next_write_char_path _00259_ vssd1
+ vssd1 vccd1 vccd1 top.header_synthesis.write_char_path sky130_fd_sc_hd__dfrtp_1
X_10835_ clknet_leaf_79_clk _01421_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06893__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_24_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_8
X_10766_ clknet_leaf_44_clk _01365_ _00185_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[60\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10697_ clknet_leaf_119_clk _01296_ _00116_ vssd1 vssd1 vccd1 vccd1 top.path\[73\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05853__B1 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08398__A2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05605__B1 _02692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11318_ clknet_leaf_77_clk _01866_ _00673_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[61\]
+ sky130_fd_sc_hd__dfrtp_1
X_11249_ clknet_leaf_75_clk _01797_ _00604_ vssd1 vssd1 vccd1 vccd1 top.hTree.wait_cnt
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05810_ _02821_ _02826_ vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__nand2b_1
X_06790_ top.findLeastValue.val1\[40\] net131 net115 net1700 vssd1 vssd1 vccd1 vccd1
+ _02048_ sky130_fd_sc_hd__o22a_1
X_05741_ top.sram_interface.write_counter_FLV\[1\] top.sram_interface.write_counter_FLV\[0\]
+ top.sram_interface.write_counter_FLV\[2\] vssd1 vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__or3b_1
X_05672_ top.cb_syn.char_path\[65\] net554 net544 top.cb_syn.char_path\[33\] vssd1
+ vssd1 vccd1 vccd1 _02748_ sky130_fd_sc_hd__a22o_1
X_08460_ net1366 top.cb_syn.char_path_n\[116\] net222 vssd1 vssd1 vccd1 vccd1 _01634_
+ sky130_fd_sc_hd__mux2_1
X_07411_ _03988_ _04004_ top.dut.bits_in_buf_next\[0\] vssd1 vssd1 vccd1 vccd1 _04010_
+ sky130_fd_sc_hd__mux2_1
X_08391_ top.cb_syn.char_path_n\[13\] net391 net330 top.cb_syn.char_path_n\[14\] _02504_
+ vssd1 vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__a221o_1
XANTENNA__07508__S1 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_15_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_18_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07342_ _03775_ net270 _03962_ net275 net1678 vssd1 vssd1 vccd1 vccd1 _01904_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_98_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07833__A1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07273_ _03678_ _03679_ _03912_ vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__nand3b_1
X_06224_ top.cw1\[4\] _02993_ vssd1 vssd1 vccd1 vccd1 _03092_ sky130_fd_sc_hd__xor2_1
XANTENNA__05844__B1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09012_ top.WB.CPU_DAT_O\[13\] net1175 net319 vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__mux2_1
X_06155_ top.hTree.write_HT_fin top.WorR net548 vssd1 vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__o21a_1
Xhold100 top.hTree.node_reg\[10\] vssd1 vssd1 vccd1 vccd1 net1053 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 top.cb_syn.char_path\[92\] vssd1 vssd1 vccd1 vccd1 net1075 sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 top.hTree.tree_reg\[53\] vssd1 vssd1 vccd1 vccd1 net1064 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout201_A net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold133 top.cb_syn.char_path\[5\] vssd1 vssd1 vccd1 vccd1 net1086 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 top.path\[82\] vssd1 vssd1 vccd1 vccd1 net1097 sky130_fd_sc_hd__dlygate4sd3_1
X_06086_ _02958_ vssd1 vssd1 vccd1 vccd1 _02959_ sky130_fd_sc_hd__inv_2
Xhold155 top.cb_syn.char_path\[27\] vssd1 vssd1 vccd1 vccd1 net1108 sky130_fd_sc_hd__dlygate4sd3_1
Xteam_05_907 vssd1 vssd1 vccd1 vccd1 team_05_907/HI gpio_out[22] sky130_fd_sc_hd__conb_1
Xteam_05_918 vssd1 vssd1 vccd1 vccd1 team_05_918/HI gpio_out[33] sky130_fd_sc_hd__conb_1
Xhold177 top.path\[64\] vssd1 vssd1 vccd1 vccd1 net1130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 top.path\[79\] vssd1 vssd1 vccd1 vccd1 net1119 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout624 net625 vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__clkbuf_2
Xfanout613 net614 vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__clkbuf_2
Xfanout602 net607 vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__clkbuf_2
Xhold188 top.path\[122\] vssd1 vssd1 vccd1 vccd1 net1141 sky130_fd_sc_hd__dlygate4sd3_1
Xteam_05_929 vssd1 vssd1 vccd1 vccd1 gpio_oeb[9] team_05_929/LO sky130_fd_sc_hd__conb_1
Xhold199 top.path\[110\] vssd1 vssd1 vccd1 vccd1 net1152 sky130_fd_sc_hd__dlygate4sd3_1
X_09914_ net740 net580 vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__and2_1
Xfanout646 net647 vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__buf_2
XANTENNA__07962__A net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout635 net636 vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__clkbuf_2
X_09845_ net760 net600 vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__and2_1
XANTENNA_input6_A DAT_I[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout657 net664 vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__07364__A3 _03547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout191_X net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout679 net681 vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__clkbuf_2
Xfanout668 net669 vssd1 vssd1 vccd1 vccd1 net668 sky130_fd_sc_hd__clkbuf_2
XFILLER_85_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09776_ net788 net628 vssd1 vssd1 vccd1 vccd1 _00390_ sky130_fd_sc_hd__and2_1
X_06988_ _03642_ _03643_ _03644_ _03645_ vssd1 vssd1 vccd1 vccd1 _03646_ sky130_fd_sc_hd__and4_1
X_08727_ net447 _04188_ net1116 vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__o21a_1
X_05939_ top.WB.CPU_DAT_O\[16\] net1118 net304 vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout835_A net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ top.cb_syn.setup top.cb_syn.curr_state\[0\] net431 vssd1 vssd1 vccd1 vccd1
+ _04862_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09889__A net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07609_ top.hTree.state\[3\] top.hTree.state\[4\] net264 vssd1 vssd1 vccd1 vccd1
+ _04192_ sky130_fd_sc_hd__o21a_1
X_08589_ _04813_ top.cb_syn.char_index\[2\] _04807_ vssd1 vssd1 vccd1 vccd1 _01512_
+ sky130_fd_sc_hd__mux2_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__06875__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10620_ net862 net702 vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__and2_1
X_10551_ net829 net669 vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__and2_1
X_10482_ net870 net710 vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__and2_1
XANTENNA__08017__B net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11103_ clknet_leaf_13_clk _01651_ _00458_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_11034_ clknet_leaf_18_clk _01582_ _00389_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[64\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_49_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11867_ clknet_leaf_100_clk _02383_ _01222_ vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__dfrtp_1
X_11798_ clknet_leaf_58_clk _00016_ _01153_ vssd1 vssd1 vccd1 vccd1 top.controller.state_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10818_ clknet_leaf_105_clk _01404_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10749_ clknet_leaf_2_clk _01348_ _00168_ vssd1 vssd1 vccd1 vccd1 top.path\[125\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09017__A0 top.WB.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06251__B1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07960_ _02496_ _04192_ _04193_ vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__o21bai_1
XFILLER_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09326__X top.controller.fin_TRN vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06911_ top.findLeastValue.val2\[28\] net147 net121 _03597_ vssd1 vssd1 vccd1 vccd1
+ _01970_ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_4_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_8
X_07891_ net482 _04417_ vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__or2_1
X_06842_ _02476_ net152 net126 _03560_ vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__a2bb2o_1
X_09630_ net750 net590 vssd1 vssd1 vccd1 vccd1 _00244_ sky130_fd_sc_hd__and2_1
X_09561_ net795 net635 vssd1 vssd1 vccd1 vccd1 _00175_ sky130_fd_sc_hd__and2_1
X_06773_ top.findLeastValue.least1\[7\] net288 net117 vssd1 vssd1 vccd1 vccd1 _02063_
+ sky130_fd_sc_hd__o21a_1
X_05724_ top.TRN_char_index\[3\] net41 net720 vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__mux2_1
X_08512_ net1136 top.cb_syn.char_path_n\[64\] net233 vssd1 vssd1 vccd1 vccd1 _01582_
+ sky130_fd_sc_hd__mux2_1
X_09492_ net731 net571 vssd1 vssd1 vccd1 vccd1 _00106_ sky130_fd_sc_hd__and2_1
X_08443_ _02929_ _04801_ _04543_ vssd1 vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout249_A _04199_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05655_ top.cb_syn.char_path\[4\] top.sram_interface.word_cnt\[0\] net316 top.cb_syn.char_path\[100\]
+ vssd1 vssd1 vccd1 vccd1 _02734_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout151_A net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08059__A1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08374_ _02503_ _04731_ _04732_ vssd1 vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__nor3_1
X_05586_ net1208 net138 _02676_ net174 vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_102_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07325_ _03718_ _03950_ vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout416_A _02759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09008__A0 top.WB.CPU_DAT_O\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07256_ _03708_ _03899_ _03702_ vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__a21o_1
X_06207_ net495 _03073_ _03075_ _02943_ net467 vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__o221a_1
X_07187_ _03843_ _03844_ vssd1 vssd1 vccd1 vccd1 _03845_ sky130_fd_sc_hd__and2b_1
X_06138_ net1307 net143 _03009_ net159 vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout785_A net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06069_ top.sram_interface.init_counter\[3\] _02911_ vssd1 vssd1 vccd1 vccd1 _02944_
+ sky130_fd_sc_hd__or2_1
XFILLER_105_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout421 net422 vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__clkbuf_2
Xfanout432 net435 vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__buf_2
Xfanout410 _02788_ vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__clkbuf_4
Xfanout454 net455 vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__buf_2
XFILLER_98_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout465 top.controller.state_reg\[5\] vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__clkbuf_2
Xfanout443 net444 vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__buf_2
Xfanout476 net477 vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__clkbuf_4
XFILLER_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout487 net493 vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__clkbuf_2
Xfanout498 top.findLeastValue.histo_index\[5\] vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__buf_2
X_09828_ net768 net608 vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__and2_1
XFILLER_104_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09759_ net742 net582 vssd1 vssd1 vccd1 vccd1 _00373_ sky130_fd_sc_hd__and2_1
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout838_X net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09412__A net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11721_ clknet_leaf_122_clk _02254_ _01076_ vssd1 vssd1 vccd1 vccd1 top.path\[52\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05520__A2 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11652_ clknet_leaf_112_clk _02185_ _01007_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11450__Q top.findLeastValue.least2\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10603_ net751 net591 vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_12_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11583_ clknet_leaf_14_clk _02131_ _00938_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_40_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10534_ net859 net699 vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__and2_1
X_10465_ net728 net568 vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_79_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10396_ net763 net603 vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__and2_1
XFILLER_2_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__05587__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11017_ clknet_leaf_8_clk _01565_ _00372_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07733__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_0_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05440_ _02480_ _02547_ vssd1 vssd1 vccd1 vccd1 _02548_ sky130_fd_sc_hd__nor2_2
X_05371_ top.findLeastValue.least2\[1\] vssd1 vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__inv_2
XANTENNA__11360__Q top.findLeastValue.sum\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07110_ _03764_ _03767_ vssd1 vssd1 vccd1 vccd1 _03768_ sky130_fd_sc_hd__nor2_1
X_08090_ top.cb_syn.char_path_n\[124\] net206 _04572_ vssd1 vssd1 vccd1 vccd1 _01770_
+ sky130_fd_sc_hd__o21a_1
Xclkload20 clknet_leaf_121_clk vssd1 vssd1 vccd1 vccd1 clkload20/Y sky130_fd_sc_hd__clkinv_2
Xclkload53 clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 clkload53/Y sky130_fd_sc_hd__inv_6
X_07041_ _03696_ _03698_ vssd1 vssd1 vccd1 vccd1 _03699_ sky130_fd_sc_hd__nor2_1
Xclkload31 clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 clkload31/X sky130_fd_sc_hd__clkbuf_4
Xclkload42 clknet_leaf_110_clk vssd1 vssd1 vccd1 vccd1 clkload42/Y sky130_fd_sc_hd__bufinv_16
Xclkload64 clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 clkload64/Y sky130_fd_sc_hd__inv_6
Xclkload75 clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 clkload75/Y sky130_fd_sc_hd__inv_6
Xclkload86 clknet_leaf_95_clk vssd1 vssd1 vccd1 vccd1 clkload86/Y sky130_fd_sc_hd__clkinv_2
Xclkload97 clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 clkload97/Y sky130_fd_sc_hd__inv_8
XANTENNA__08764__A2 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06775__B2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08992_ top.WB.CPU_DAT_O\[0\] net1117 net324 vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__mux2_1
X_07943_ net444 net1583 net255 top.findLeastValue.sum\[0\] _04460_ vssd1 vssd1 vccd1
+ vccd1 _01805_ sky130_fd_sc_hd__a221o_1
XFILLER_95_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07874_ top.findLeastValue.sum\[13\] top.hTree.tree_reg\[13\] net283 vssd1 vssd1
+ vccd1 vccd1 _04405_ sky130_fd_sc_hd__mux2_1
XFILLER_110_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_09613_ net802 net642 vssd1 vssd1 vccd1 vccd1 _00227_ sky130_fd_sc_hd__and2_1
XFILLER_56_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06825_ top.findLeastValue.val1\[5\] net131 net115 top.compVal\[5\] vssd1 vssd1 vccd1
+ vccd1 _02013_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout366_A net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09544_ net748 net588 vssd1 vssd1 vccd1 vccd1 _00158_ sky130_fd_sc_hd__and2_1
X_06756_ _02410_ top.findLeastValue.val2\[39\] _03533_ _03543_ vssd1 vssd1 vccd1 vccd1
+ _03544_ sky130_fd_sc_hd__a22o_1
X_06687_ top.findLeastValue.val2\[14\] _02435_ top.compVal\[15\] _02493_ vssd1 vssd1
+ vccd1 vccd1 _03475_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout154_X net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05707_ net6 net415 net308 top.WB.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 _02351_
+ sky130_fd_sc_hd__o22a_1
X_09475_ net732 net572 vssd1 vssd1 vccd1 vccd1 _00089_ sky130_fd_sc_hd__and2_1
X_08426_ top.cb_syn.char_path_n\[53\] net392 net331 top.cb_syn.char_path_n\[54\] _02505_
+ vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__a221o_1
X_05638_ _02718_ _02719_ vssd1 vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__or2_1
XANTENNA__05502__A2 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout700_A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08357_ top.cb_syn.char_path_n\[82\] net332 _04715_ vssd1 vssd1 vccd1 vccd1 _04716_
+ sky130_fd_sc_hd__a21oi_1
X_05569_ top.cb_syn.char_path\[82\] net551 net543 top.cb_syn.char_path\[50\] vssd1
+ vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__a22o_1
XANTENNA__09886__B net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09378__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload3 clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clkload3/X sky130_fd_sc_hd__clkbuf_8
X_08288_ top.cb_syn.char_path_n\[25\] net206 _04671_ vssd1 vssd1 vccd1 vccd1 _01671_
+ sky130_fd_sc_hd__o21a_1
X_07308_ _03788_ _03935_ vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__xnor2_1
XANTENNA__05919__B net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07239_ _03817_ _03820_ _03829_ vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__a21oi_1
X_10250_ net862 net702 vssd1 vssd1 vccd1 vccd1 _00864_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_115_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05494__X _02600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05569__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10181_ net842 net682 vssd1 vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__and2_1
XFILLER_105_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout240 net243 vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__buf_2
Xfanout262 net267 vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__clkbuf_4
Xfanout273 _03658_ vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__clkbuf_4
Xfanout251 net252 vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__buf_2
XFILLER_115_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xfanout295 _05102_ vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__buf_2
Xfanout284 _04197_ vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_45_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ clknet_leaf_115_clk _02237_ _01059_ vssd1 vssd1 vccd1 vccd1 top.path\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09315__S0 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11635_ clknet_leaf_56_clk top.dut.bit_buf_next\[7\] _00990_ vssd1 vssd1 vccd1 vccd1
+ top.dut.bit_buf\[7\] sky130_fd_sc_hd__dfrtp_1
X_11566_ clknet_leaf_38_clk _02114_ _00921_ vssd1 vssd1 vccd1 vccd1 top.header_synthesis.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07246__A2 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10517_ net868 net708 vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__and2_1
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11497_ clknet_leaf_92_clk _02045_ _00852_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[37\]
+ sky130_fd_sc_hd__dfstp_1
X_10448_ net753 net593 vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__and2_1
X_10379_ net856 net696 vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__and2_1
XFILLER_97_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07954__A0 top.findLeastValue.least1\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06757__A1 _03521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11355__Q top.findLeastValue.sum\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07590_ net1521 _04176_ _04144_ vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__mux2_1
XFILLER_80_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06610_ _02409_ top.findLeastValue.val1\[41\] vssd1 vssd1 vccd1 vccd1 _03399_ sky130_fd_sc_hd__nand2_1
XANTENNA__07124__X _03782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06541_ _02421_ top.findLeastValue.val1\[29\] vssd1 vssd1 vccd1 vccd1 _03330_ sky130_fd_sc_hd__nor2_1
X_09260_ top.cb_syn.zero_count\[0\] top.cb_syn.zero_count\[1\] vssd1 vssd1 vccd1 vccd1
+ _05216_ sky130_fd_sc_hd__or2_1
XANTENNA__08131__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06472_ net1388 _03293_ _03294_ vssd1 vssd1 vccd1 vccd1 _02106_ sky130_fd_sc_hd__a21o_1
X_05423_ top.cb_syn.zero_count\[0\] vssd1 vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__inv_2
X_08211_ top.cb_syn.char_path_n\[64\] net388 net347 top.cb_syn.char_path_n\[62\] net192
+ vssd1 vssd1 vccd1 vccd1 _04633_ sky130_fd_sc_hd__a221o_1
XANTENNA__08891__A net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05496__B2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09191_ top.controller.fin_reg\[1\] top.controller.fin_reg\[2\] top.controller.fin_reg\[3\]
+ top.controller.fin_reg\[5\] vssd1 vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__nor4_1
XFILLER_21_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08142_ top.cb_syn.char_path_n\[98\] net203 _04598_ vssd1 vssd1 vccd1 vccd1 _01744_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__05579__X _02671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05354_ top.findLeastValue.val1\[40\] vssd1 vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__inv_2
Xclkload120 clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 clkload120/Y sky130_fd_sc_hd__clkinv_4
X_08073_ _02553_ _02867_ _02870_ vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__and3_1
XANTENNA__05739__B net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout114_A net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07024_ _03678_ _03681_ vssd1 vssd1 vccd1 vccd1 _03682_ sky130_fd_sc_hd__nand2_1
XANTENNA__08830__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_08975_ top.WB.CPU_DAT_O\[17\] net1377 net323 vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__mux2_1
Xhold15 top.sram_interface.init_counter\[20\] vssd1 vssd1 vccd1 vccd1 net968 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 top.hTree.node_reg\[55\] vssd1 vssd1 vccd1 vccd1 net979 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 top.hTree.node_reg\[59\] vssd1 vssd1 vccd1 vccd1 net990 sky130_fd_sc_hd__dlygate4sd3_1
X_07926_ net488 _04445_ vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_110_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold48 top.hTree.node_reg\[57\] vssd1 vssd1 vccd1 vccd1 net1001 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold59 top.hTree.node_reg\[15\] vssd1 vssd1 vccd1 vccd1 net1012 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08370__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07857_ net426 _04390_ _04391_ net259 vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout748_A net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07788_ net443 net1408 net254 top.findLeastValue.sum\[31\] _04336_ vssd1 vssd1 vccd1
+ vccd1 _01836_ sky130_fd_sc_hd__a221o_1
XFILLER_44_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06808_ top.findLeastValue.val1\[22\] net128 net112 top.compVal\[22\] vssd1 vssd1
+ vccd1 vccd1 _02030_ sky130_fd_sc_hd__o22a_1
X_09527_ net755 net595 vssd1 vssd1 vccd1 vccd1 _00141_ sky130_fd_sc_hd__and2_1
X_06739_ _02412_ top.findLeastValue.val2\[36\] top.findLeastValue.val2\[35\] _02413_
+ vssd1 vssd1 vccd1 vccd1 _03527_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout536_X net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09458_ net869 net709 vssd1 vssd1 vccd1 vccd1 _00072_ sky130_fd_sc_hd__and2_1
XFILLER_101_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08409_ top.cb_syn.char_path_n\[29\] net392 _04767_ net511 _02504_ vssd1 vssd1 vccd1
+ vccd1 _04768_ sky130_fd_sc_hd__a221o_1
X_09389_ net405 _04256_ vssd1 vssd1 vccd1 vccd1 _05270_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_22_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08425__A1 _02506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11420_ clknet_leaf_103_clk _01968_ _00775_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[26\]
+ sky130_fd_sc_hd__dfstp_1
X_11351_ clknet_leaf_93_clk _01899_ _00706_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10302_ net799 net639 vssd1 vssd1 vccd1 vccd1 _00916_ sky130_fd_sc_hd__and2_1
XFILLER_106_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11282_ clknet_leaf_80_clk net1540 _00637_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_105_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10233_ net840 net680 vssd1 vssd1 vccd1 vccd1 _00847_ sky130_fd_sc_hd__and2_1
XANTENNA_input44_A nrst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10164_ net827 net667 vssd1 vssd1 vccd1 vccd1 _00778_ sky130_fd_sc_hd__and2_1
XANTENNA__05962__A2 _02899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10095_ net812 net652 vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__and2_1
XANTENNA__08900__A2 _04187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05714__A2 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10997_ clknet_leaf_29_clk _01545_ _00352_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07872__C1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11618_ clknet_leaf_62_clk _02166_ _00973_ vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__dfrtp_1
XFILLER_7_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xhold507 _01831_ vssd1 vssd1 vccd1 vccd1 net1460 sky130_fd_sc_hd__dlygate4sd3_1
X_11549_ clknet_leaf_123_clk _02097_ _00904_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[22\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold518 top.path\[69\] vssd1 vssd1 vccd1 vccd1 net1471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold529 top.hist_data_o\[18\] vssd1 vssd1 vccd1 vccd1 net1482 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05972_ top.sram_interface.init_counter\[7\] top.sram_interface.init_counter\[6\]
+ _02907_ vssd1 vssd1 vccd1 vccd1 _02908_ sky130_fd_sc_hd__and3_1
X_08760_ top.path\[102\] top.path\[103\] net528 vssd1 vssd1 vccd1 vccd1 _04943_ sky130_fd_sc_hd__mux2_1
X_08691_ top.cb_syn.zeroes\[4\] _04878_ vssd1 vssd1 vccd1 vccd1 _04889_ sky130_fd_sc_hd__or2_1
X_07711_ top.hTree.tree_reg\[46\] top.findLeastValue.least2\[0\] net248 vssd1 vssd1
+ vccd1 vccd1 _04275_ sky130_fd_sc_hd__mux2_1
X_07642_ net262 _04217_ _04218_ net1367 net445 vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_0_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07573_ top.cb_syn.max_index\[5\] _04149_ vssd1 vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__xnor2_1
X_09312_ top.histogram.total\[16\] net408 net326 top.histogram.total\[17\] net436
+ vssd1 vssd1 vccd1 vccd1 _05247_ sky130_fd_sc_hd__o221a_1
X_06524_ _03272_ _03315_ vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__nor2_1
X_09243_ net1098 _05206_ net296 vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_header\[2\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout231_A net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06455_ top.histogram.total\[7\] top.histogram.total\[6\] vssd1 vssd1 vccd1 vccd1
+ _03278_ sky130_fd_sc_hd__and2_1
XFILLER_119_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05406_ top.cb_syn.zeroes\[2\] vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__inv_2
X_09174_ top.cb_syn.char_path_n\[2\] net517 net474 net530 vssd1 vssd1 vccd1 vccd1
+ _05167_ sky130_fd_sc_hd__and4b_1
XANTENNA__06345__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06853__B _03325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06386_ net1139 _03228_ net300 vssd1 vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__mux2_1
X_08125_ top.cb_syn.char_path_n\[107\] net374 net334 top.cb_syn.char_path_n\[105\]
+ net179 vssd1 vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__a221o_1
X_05337_ top.compVal\[4\] vssd1 vssd1 vccd1 vccd1 _02445_ sky130_fd_sc_hd__inv_2
XANTENNA__07030__A top.findLeastValue.val1\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__05469__B net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout117_X net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08056_ net505 net507 net246 _04540_ vssd1 vssd1 vccd1 vccd1 _04548_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_112_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput49 net49 vssd1 vssd1 vccd1 vccd1 ADR_O[14] sky130_fd_sc_hd__buf_2
X_07007_ top.findLeastValue.val1\[37\] top.findLeastValue.val2\[37\] vssd1 vssd1 vccd1
+ vccd1 _03665_ sky130_fd_sc_hd__nand2_1
XANTENNA__05641__B2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout865_A net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout486_X net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08958_ top.WB.CPU_DAT_O\[15\] top.cb_syn.h_element\[47\] net369 vssd1 vssd1 vccd1
+ vccd1 _01352_ sky130_fd_sc_hd__mux2_1
X_08889_ _02459_ _02795_ net397 vssd1 vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__o21a_1
X_07909_ top.findLeastValue.sum\[6\] top.hTree.tree_reg\[6\] net284 vssd1 vssd1 vccd1
+ vccd1 _04433_ sky130_fd_sc_hd__mux2_1
X_10920_ clknet_leaf_34_clk _01475_ _00275_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.i\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_71_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10851_ clknet_leaf_109_clk _01437_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[43\]
+ sky130_fd_sc_hd__dfxtp_1
X_10782_ clknet_leaf_47_clk _01381_ _00201_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_40_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11403_ clknet_leaf_96_clk _01951_ _00758_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[9\]
+ sky130_fd_sc_hd__dfstp_1
X_11334_ clknet_leaf_54_clk _01882_ _00689_ vssd1 vssd1 vccd1 vccd1 top.dut.out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_55_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08470__S net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11265_ clknet_leaf_104_clk _01813_ _00620_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05395__A top.cb_syn.end_cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10216_ net814 net654 vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__and2_1
X_11196_ clknet_leaf_16_clk _01744_ _00551_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[98\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_94_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06003__B net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10147_ net825 net665 vssd1 vssd1 vccd1 vccd1 _00761_ sky130_fd_sc_hd__and2_1
X_10078_ net852 net692 vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_113_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08993__X _05088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05699__B2 top.WB.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_06240_ _03094_ _03100_ _03106_ _03107_ vssd1 vssd1 vccd1 vccd1 _03108_ sky130_fd_sc_hd__or4_1
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06171_ top.findLeastValue.histo_index\[6\] net499 net412 _03013_ vssd1 vssd1 vccd1
+ vccd1 _03041_ sky130_fd_sc_hd__and4_1
Xhold326 top.histogram.sram_out\[28\] vssd1 vssd1 vccd1 vccd1 net1279 sky130_fd_sc_hd__dlygate4sd3_1
Xwire290 _02837_ vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__buf_1
Xhold315 top.cb_syn.char_path\[50\] vssd1 vssd1 vccd1 vccd1 net1268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold304 top.path\[55\] vssd1 vssd1 vccd1 vccd1 net1257 sky130_fd_sc_hd__dlygate4sd3_1
X_09930_ net783 net623 vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__and2_1
Xhold348 top.histogram.sram_out\[26\] vssd1 vssd1 vccd1 vccd1 net1301 sky130_fd_sc_hd__dlygate4sd3_1
Xhold359 top.cb_syn.char_path\[18\] vssd1 vssd1 vccd1 vccd1 net1312 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05623__B2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold337 top.path\[78\] vssd1 vssd1 vccd1 vccd1 net1290 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout806 net807 vssd1 vssd1 vccd1 vccd1 net806 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09861_ net771 net611 vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__and2_1
Xfanout839 net841 vssd1 vssd1 vccd1 vccd1 net839 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout817 net824 vssd1 vssd1 vccd1 vccd1 net817 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout828 net829 vssd1 vssd1 vccd1 vccd1 net828 sky130_fd_sc_hd__clkbuf_2
X_09792_ net773 net613 vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__and2_1
X_08812_ _04993_ _04994_ _04991_ vssd1 vssd1 vccd1 vccd1 _04995_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_5_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08743_ net432 net524 vssd1 vssd1 vccd1 vccd1 _04926_ sky130_fd_sc_hd__nand2_1
X_05955_ top.WB.CPU_DAT_O\[0\] net1334 net307 vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout181_A net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout279_A _04198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08674_ _04870_ _04874_ vssd1 vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__or2_4
X_05886_ _02859_ _02860_ top.cb_syn.h_element\[54\] vssd1 vssd1 vccd1 vccd1 _02861_
+ sky130_fd_sc_hd__o21a_2
XFILLER_26_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08876__A1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07625_ _04203_ _04204_ net487 vssd1 vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout446_A net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07556_ net532 top.cb_syn.h_element\[52\] net539 top.cb_syn.h_element\[61\] vssd1
+ vssd1 vccd1 vccd1 _04147_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06507_ _03281_ net1493 vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__nor2_1
X_09226_ net519 net1654 _04919_ _05192_ vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_write_char_path
+ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout234_X net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07487_ top.cb_syn.char_path_n\[32\] top.cb_syn.char_path_n\[31\] top.cb_syn.char_path_n\[30\]
+ top.cb_syn.char_path_n\[29\] net401 net352 vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__mux4_1
XFILLER_42_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_06438_ net1676 _03257_ _03264_ vssd1 vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_32_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout401_X net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09157_ top.hTree.wait_cnt net264 vssd1 vssd1 vccd1 vccd1 _05162_ sky130_fd_sc_hd__nand2_1
X_06369_ _03186_ _03217_ net301 vssd1 vssd1 vccd1 vccd1 _03218_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09053__A1 top.WB.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05862__B2 top.WB.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09088_ _03172_ _05101_ vssd1 vssd1 vccd1 vccd1 _05109_ sky130_fd_sc_hd__nor2_1
X_08108_ top.cb_syn.char_path_n\[115\] net197 _04581_ vssd1 vssd1 vccd1 vccd1 _01761_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__05767__X _02788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08039_ top.cb_syn.h_element\[54\] _02553_ vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__nor2_1
XANTENNA__06811__B1 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11050_ clknet_leaf_8_clk _01598_ _00405_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[80\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_76_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10001_ net836 net676 vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__and2_1
XFILLER_103_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07206__Y _03864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11883_ clknet_leaf_39_clk _02399_ _01238_ vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__dfrtp_1
X_10903_ clknet_leaf_39_clk top.header_synthesis.next_header\[8\] _00258_ vssd1 vssd1
+ vccd1 vccd1 top.header_synthesis.header\[8\] sky130_fd_sc_hd__dfrtp_1
X_10834_ clknet_leaf_79_clk _01420_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08465__S net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05550__B1 _02646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07827__C1 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_17_Left_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10765_ clknet_leaf_44_clk _01364_ _00184_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10696_ clknet_leaf_111_clk _01295_ _00115_ vssd1 vssd1 vccd1 vccd1 top.path\[72\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__05853__B2 top.WB.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09044__A1 top.WB.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07809__S net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11317_ clknet_leaf_76_clk _01865_ _00672_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[60\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05396__Y _02504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05605__B2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06802__B1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_26_Left_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11248_ clknet_leaf_68_clk _01796_ _00603_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.alternator_timer\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11179_ clknet_leaf_21_clk _01727_ _00534_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[81\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_95_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06030__A1 top.WB.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09325__A net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05740_ net452 _02763_ _02773_ vssd1 vssd1 vccd1 vccd1 _02775_ sky130_fd_sc_hd__a21o_1
XFILLER_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05671_ net1079 net145 _02747_ net177 vssd1 vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__a22o_1
XANTENNA__11363__Q top.findLeastValue.sum\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07410_ net354 _04001_ _04005_ _04009_ vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__a31o_1
XFILLER_90_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__05541__B1 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08375__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08390_ top.cb_syn.char_path_n\[15\] top.cb_syn.char_path_n\[16\] net514 vssd1 vssd1
+ vccd1 vccd1 _04749_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_35_Left_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07341_ _03770_ _03772_ _03774_ vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_18_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07272_ top.findLeastValue.val1\[25\] top.findLeastValue.val2\[25\] _03705_ _03910_
+ _03681_ vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__o221ai_2
XTAP_TAPCELL_ROW_98_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06223_ _02572_ _03002_ _03090_ net368 top.findLeastValue.histo_index\[3\] vssd1
+ vssd1 vccd1 vccd1 _03091_ sky130_fd_sc_hd__a32o_1
XANTENNA__09035__A1 top.WB.CPU_DAT_O\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05844__B2 top.WB.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09011_ top.WB.CPU_DAT_O\[14\] net1290 net319 vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__mux2_1
Xhold101 top.header_synthesis.header\[2\] vssd1 vssd1 vccd1 vccd1 net1054 sky130_fd_sc_hd__dlygate4sd3_1
X_06154_ _02454_ net362 net550 vssd1 vssd1 vccd1 vccd1 _03025_ sky130_fd_sc_hd__a21o_2
XPHY_EDGE_ROW_103_Right_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold123 top.cb_syn.char_path\[29\] vssd1 vssd1 vccd1 vccd1 net1076 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_44_Left_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold134 top.path\[7\] vssd1 vssd1 vccd1 vccd1 net1087 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 top.path\[30\] vssd1 vssd1 vccd1 vccd1 net1065 sky130_fd_sc_hd__dlygate4sd3_1
Xteam_05_908 vssd1 vssd1 vccd1 vccd1 team_05_908/HI gpio_out[23] sky130_fd_sc_hd__conb_1
Xhold145 top.header_synthesis.header\[1\] vssd1 vssd1 vccd1 vccd1 net1098 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06085_ top.cb_syn.char_index\[3\] _02957_ vssd1 vssd1 vccd1 vccd1 _02958_ sky130_fd_sc_hd__and2_1
Xhold167 top.cb_syn.char_path\[26\] vssd1 vssd1 vccd1 vccd1 net1120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 top.cb_syn.char_path\[65\] vssd1 vssd1 vccd1 vccd1 net1109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 top.cb_syn.char_path\[96\] vssd1 vssd1 vccd1 vccd1 net1131 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout614 net616 vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__clkbuf_2
Xhold189 top.histogram.sram_out\[14\] vssd1 vssd1 vccd1 vccd1 net1142 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout603 net607 vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__clkbuf_2
X_09913_ net740 net580 vssd1 vssd1 vccd1 vccd1 _00527_ sky130_fd_sc_hd__and2_1
Xfanout647 net44 vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__buf_4
Xfanout625 net626 vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__clkbuf_2
Xfanout636 net646 vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout396_A net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09844_ net761 net601 vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__and2_1
Xfanout658 net659 vssd1 vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__clkbuf_2
XANTENNA__05763__A top.controller.state_reg\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout669 net675 vssd1 vssd1 vccd1 vccd1 net669 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__06021__A1 top.WB.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09775_ net789 net629 vssd1 vssd1 vccd1 vccd1 _00389_ sky130_fd_sc_hd__and2_1
X_06987_ top.findLeastValue.val1\[2\] top.findLeastValue.val1\[1\] top.findLeastValue.val1\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03645_ sky130_fd_sc_hd__and3_1
X_08726_ _04905_ _04898_ top.cb_syn.i\[0\] vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__mux2_1
XFILLER_100_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05938_ top.WB.CPU_DAT_O\[17\] net1234 net304 vssd1 vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__mux2_1
X_05869_ top.sram_interface.init_counter\[17\] top.sram_interface.init_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_107_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08657_ net1634 net190 vssd1 vssd1 vccd1 vccd1 _01492_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09889__B net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout351_X net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_53_Left_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout449_X net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07608_ net461 net954 _04190_ vssd1 vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__o21a_1
XFILLER_26_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08588_ top.cb_syn.h_element\[57\] top.cb_syn.h_element\[48\] net532 vssd1 vssd1
+ vccd1 vccd1 _04813_ sky130_fd_sc_hd__mux2_1
XANTENNA__05532__B1 _02631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07539_ _04129_ vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout616_X net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_10_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10550_ net828 net668 vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__and2_1
X_09209_ top.cb_syn.char_path_n\[2\] top.cb_syn.char_path_n\[1\] _02930_ net431 vssd1
+ vssd1 vccd1 vccd1 _05185_ sky130_fd_sc_hd__a31o_1
X_10481_ net861 net701 vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__and2_1
XANTENNA__09026__A1 top.WB.CPU_DAT_O\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_62_Left_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05599__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11102_ clknet_leaf_13_clk _01650_ _00457_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold690 top.findLeastValue.sum\[24\] vssd1 vssd1 vccd1 vccd1 net1643 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11033_ clknet_leaf_43_clk _01581_ _00388_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06012__A1 top.WB.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_71_Left_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05523__B1 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11866_ clknet_leaf_121_clk _02382_ _01221_ vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__dfrtp_1
X_11797_ clknet_leaf_58_clk _00015_ _01152_ vssd1 vssd1 vccd1 vccd1 top.controller.state_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_15_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10817_ clknet_leaf_109_clk _01403_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08923__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10748_ clknet_leaf_119_clk _01347_ _00167_ vssd1 vssd1 vccd1 vccd1 top.path\[124\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10679_ clknet_leaf_123_clk _01278_ _00098_ vssd1 vssd1 vccd1 vccd1 top.path\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_93_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11358__Q top.findLeastValue.sum\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06910_ top.compVal\[28\] top.findLeastValue.val1\[28\] net162 vssd1 vssd1 vccd1
+ vccd1 _03597_ sky130_fd_sc_hd__mux2_1
XFILLER_95_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07890_ top.findLeastValue.sum\[10\] _04417_ net395 vssd1 vssd1 vccd1 vccd1 _04418_
+ sky130_fd_sc_hd__mux2_1
X_06841_ top.findLeastValue.least1\[4\] net500 _03424_ vssd1 vssd1 vccd1 vccd1 _03560_
+ sky130_fd_sc_hd__mux2_1
X_09560_ net843 net683 vssd1 vssd1 vccd1 vccd1 _00174_ sky130_fd_sc_hd__and2_1
X_06772_ top.findLeastValue.least1\[8\] net133 net117 _02767_ vssd1 vssd1 vccd1 vccd1
+ _02064_ sky130_fd_sc_hd__o22a_1
X_05723_ top.TRN_char_index\[4\] net42 net720 vssd1 vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__mux2_1
X_08511_ net1109 top.cb_syn.char_path_n\[65\] net234 vssd1 vssd1 vccd1 vccd1 _01583_
+ sky130_fd_sc_hd__mux2_1
X_09491_ net728 net568 vssd1 vssd1 vccd1 vccd1 _00105_ sky130_fd_sc_hd__and2_1
X_08442_ top.cb_syn.cb_length\[1\] top.cb_syn.cb_length\[0\] vssd1 vssd1 vccd1 vccd1
+ _04801_ sky130_fd_sc_hd__nand2b_1
X_05654_ top.cb_syn.char_path\[68\] net552 net543 top.cb_syn.char_path\[36\] vssd1
+ vssd1 vccd1 vccd1 _02733_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout144_A net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08059__A2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08373_ _04728_ _04729_ _04730_ net507 _02504_ vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__o221a_1
X_05585_ top.histogram.sram_out\[16\] net364 _02674_ _02675_ vssd1 vssd1 vccd1 vccd1
+ _02676_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_102_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08833__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07324_ _03719_ _03944_ vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__nand2b_1
X_07255_ _03809_ _03816_ _03685_ vssd1 vssd1 vccd1 vccd1 _03899_ sky130_fd_sc_hd__a21o_1
X_06206_ _02945_ _03074_ vssd1 vssd1 vccd1 vccd1 _03075_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout311_A _02690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout409_A _02788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06353__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07186_ top.findLeastValue.val1\[41\] top.findLeastValue.val2\[41\] vssd1 vssd1 vccd1
+ vccd1 _03844_ sky130_fd_sc_hd__nand2_1
X_06137_ _02983_ _02986_ _03008_ vssd1 vssd1 vccd1 vccd1 _03009_ sky130_fd_sc_hd__or3_1
X_06068_ _02942_ vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__inv_2
Xfanout422 _02599_ vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__clkbuf_4
Xfanout400 net402 vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__buf_4
XANTENNA__05596__A3 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout411 _02788_ vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__06793__A2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout455 net72 vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__buf_2
Xfanout466 top.controller.state_reg\[4\] vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__clkbuf_4
XANTENNA__05493__A net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout444 net448 vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__clkbuf_2
Xfanout433 net435 vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__clkbuf_2
Xfanout477 net481 vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__clkbuf_4
Xfanout499 top.findLeastValue.histo_index\[5\] vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__dlymetal6s2s_1
X_09827_ net768 net608 vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__and2_1
Xfanout488 net493 vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__clkbuf_2
XFILLER_104_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09758_ net739 net579 vssd1 vssd1 vccd1 vccd1 _00372_ sky130_fd_sc_hd__and2_1
X_08709_ _04900_ vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_68_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09689_ net785 net625 vssd1 vssd1 vccd1 vccd1 _00303_ sky130_fd_sc_hd__and2_1
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11720_ clknet_leaf_122_clk _02253_ _01075_ vssd1 vssd1 vccd1 vccd1 top.path\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09412__B _04221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11651_ clknet_leaf_112_clk _02184_ _01006_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11582_ clknet_leaf_108_clk _02130_ _00937_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10602_ net810 net650 vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_12_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10533_ net860 net700 vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__and2_1
XFILLER_22_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08207__C1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10464_ net728 net568 vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_79_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10395_ net763 net603 vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__and2_1
XFILLER_111_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08930__A0 top.WB.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11016_ clknet_leaf_6_clk _01564_ _00371_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07733__A1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_48_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09238__A1 top.cb_syn.char_index\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11849_ clknet_leaf_116_clk _02365_ _01204_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[27\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08653__S net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05370_ top.findLeastValue.least2\[2\] vssd1 vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__inv_2
XANTENNA__08997__A0 top.WB.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload10 clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clkload10/X sky130_fd_sc_hd__clkbuf_8
Xclkload43 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 clkload43/Y sky130_fd_sc_hd__inv_8
Xclkload21 clknet_leaf_123_clk vssd1 vssd1 vccd1 vccd1 clkload21/X sky130_fd_sc_hd__clkbuf_8
Xclkload32 clknet_leaf_114_clk vssd1 vssd1 vccd1 vccd1 clkload32/X sky130_fd_sc_hd__clkbuf_8
X_07040_ top.findLeastValue.val1\[29\] top.findLeastValue.val2\[29\] vssd1 vssd1 vccd1
+ vccd1 _03698_ sky130_fd_sc_hd__nor2_1
Xclkload54 clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 clkload54/Y sky130_fd_sc_hd__bufinv_16
Xclkload65 clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 clkload65/Y sky130_fd_sc_hd__inv_6
Xclkload76 clknet_leaf_79_clk vssd1 vssd1 vccd1 vccd1 clkload76/X sky130_fd_sc_hd__clkbuf_4
Xclkload87 clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 clkload87/Y sky130_fd_sc_hd__inv_6
Xclkload98 clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 clkload98/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__06775__A2 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05578__A3 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08991_ top.WB.CPU_DAT_O\[1\] net1121 net324 vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__mux2_1
X_07942_ net429 _04458_ _04459_ net260 vssd1 vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__o211a_1
XFILLER_110_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07873_ net441 net1582 net252 top.findLeastValue.sum\[14\] _04404_ vssd1 vssd1 vccd1
+ vccd1 _01819_ sky130_fd_sc_hd__a221o_1
X_09612_ net851 net691 vssd1 vssd1 vccd1 vccd1 _00226_ sky130_fd_sc_hd__and2_1
XFILLER_55_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06824_ top.findLeastValue.val1\[6\] net130 net114 net1689 vssd1 vssd1 vccd1 vccd1
+ _02014_ sky130_fd_sc_hd__o22a_1
X_09543_ net746 net586 vssd1 vssd1 vccd1 vccd1 _00157_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_104_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout261_A net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout359_A net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06755_ _02411_ top.findLeastValue.val2\[38\] _03531_ _03542_ vssd1 vssd1 vccd1 vccd1
+ _03543_ sky130_fd_sc_hd__a22o_1
X_05706_ net7 net417 net359 top.WB.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1 _02352_
+ sky130_fd_sc_hd__a22o_1
X_06686_ _03471_ _03472_ _03473_ vssd1 vssd1 vccd1 vccd1 _03474_ sky130_fd_sc_hd__a21o_1
X_09474_ net750 net590 vssd1 vssd1 vccd1 vccd1 _00088_ sky130_fd_sc_hd__and2_1
X_08425_ _02506_ top.cb_syn.char_path_n\[56\] _04783_ net511 vssd1 vssd1 vccd1 vccd1
+ _04784_ sky130_fd_sc_hd__o211a_1
X_05637_ top.cb_syn.char_path\[7\] net558 net313 top.cb_syn.char_path\[103\] vssd1
+ vssd1 vccd1 vccd1 _02719_ sky130_fd_sc_hd__a22o_1
X_08356_ top.cb_syn.char_path_n\[81\] net391 _04698_ net510 net508 vssd1 vssd1 vccd1
+ vccd1 _04715_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout526_A top.translation.index\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload4 clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clkload4/X sky130_fd_sc_hd__clkbuf_8
X_05568_ net1328 net139 _02661_ net175 vssd1 vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_63_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07307_ net269 _03937_ _03938_ net274 top.findLeastValue.sum\[19\] vssd1 vssd1 vccd1
+ vccd1 _01915_ sky130_fd_sc_hd__a32o_1
XANTENNA__08988__A0 top.WB.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout314_X net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08287_ top.cb_syn.char_path_n\[26\] net384 net344 top.cb_syn.char_path_n\[24\] net189
+ vssd1 vssd1 vccd1 vccd1 _04671_ sky130_fd_sc_hd__a221o_1
X_05499_ _02602_ _02603_ net477 vssd1 vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__o21a_1
X_07238_ net271 _03877_ _03886_ net276 net1631 vssd1 vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__a32o_1
X_07169_ _03825_ _03826_ vssd1 vssd1 vccd1 vccd1 _03827_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_115_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07963__A1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07621__C_N net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10180_ net842 net682 vssd1 vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__and2_1
Xfanout230 net235 vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__clkbuf_2
Xfanout241 net243 vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__buf_2
XFILLER_115_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06112__A top.cb_syn.char_index\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout263 net266 vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__buf_2
XFILLER_59_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout252 net256 vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__clkbuf_2
Xfanout274 _03658_ vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__buf_2
Xfanout296 _04918_ vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__clkbuf_4
Xfanout285 net286 vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__clkbuf_4
XFILLER_74_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08039__A top.cb_syn.h_element\[54\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11703_ clknet_leaf_115_clk _02236_ _01058_ vssd1 vssd1 vccd1 vccd1 top.path\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11634_ clknet_leaf_56_clk top.dut.bit_buf_next\[6\] _00989_ vssd1 vssd1 vccd1 vccd1
+ top.dut.bit_buf\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_91_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08979__A0 top.WB.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09315__S1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11565_ clknet_leaf_38_clk _02113_ _00920_ vssd1 vssd1 vccd1 vccd1 top.header_synthesis.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10516_ net868 net708 vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__and2_1
XANTENNA__05398__A net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11496_ clknet_leaf_92_clk _02044_ _00851_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[36\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__06454__A1 _03269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10447_ net748 net588 vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__and2_1
X_10378_ net854 net694 vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__and2_1
XFILLER_97_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_90_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05717__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_9_Left_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06540_ _02420_ top.findLeastValue.val1\[30\] top.findLeastValue.val1\[29\] _02421_
+ vssd1 vssd1 vccd1 vccd1 _03329_ sky130_fd_sc_hd__a22o_1
X_06471_ top.histogram.total\[31\] top.histogram.total\[30\] _03292_ vssd1 vssd1 vccd1
+ vccd1 _03294_ sky130_fd_sc_hd__and3b_1
XANTENNA__11371__Q top.findLeastValue.sum\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05496__A2 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06142__B1 _02767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08210_ top.cb_syn.char_path_n\[64\] net209 _04632_ vssd1 vssd1 vccd1 vccd1 _01710_
+ sky130_fd_sc_hd__o21a_1
X_05422_ net480 vssd1 vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__inv_2
XANTENNA__07890__A0 top.findLeastValue.sum\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09190_ top.hTree.state\[6\] _05099_ _05175_ net1502 vssd1 vssd1 vccd1 vccd1 _00025_
+ sky130_fd_sc_hd__a22o_1
XFILLER_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08141_ top.cb_syn.char_path_n\[99\] net381 net339 top.cb_syn.char_path_n\[97\] net185
+ vssd1 vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__a221o_1
XANTENNA__08434__A2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05353_ top.findLeastValue.val1\[42\] vssd1 vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__inv_2
XFILLER_119_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_08072_ top.cb_syn.left_check top.cb_syn.h_element\[54\] _02553_ _02858_ vssd1 vssd1
+ vccd1 vccd1 _04559_ sky130_fd_sc_hd__or4b_1
Xclkload121 clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 clkload121/Y sky130_fd_sc_hd__clkinv_8
Xclkload110 clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 clkload110/Y sky130_fd_sc_hd__clkinv_2
XFILLER_106_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07023_ _03679_ _03680_ vssd1 vssd1 vccd1 vccd1 _03681_ sky130_fd_sc_hd__and2_1
XANTENNA__05595__X _02684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08974_ top.WB.CPU_DAT_O\[18\] net1132 net323 vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold16 top.hTree.node_reg\[53\] vssd1 vssd1 vccd1 vccd1 net969 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 top.hTree.node_reg\[50\] vssd1 vssd1 vccd1 vccd1 net980 sky130_fd_sc_hd__dlygate4sd3_1
X_07925_ top.findLeastValue.sum\[3\] _04445_ net398 vssd1 vssd1 vccd1 vccd1 _04446_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07028__A top.findLeastValue.val1\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold38 top.hTree.node_reg\[12\] vssd1 vssd1 vccd1 vccd1 net991 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_110_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout476_A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold49 top.hTree.node_reg\[56\] vssd1 vssd1 vccd1 vccd1 net1002 sky130_fd_sc_hd__dlygate4sd3_1
X_07856_ net483 _04389_ vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__or2_1
XANTENNA__05708__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07787_ net430 _04334_ _04335_ net261 vssd1 vssd1 vccd1 vccd1 _04336_ sky130_fd_sc_hd__o211a_1
X_06807_ top.findLeastValue.val1\[23\] net128 net112 net1673 vssd1 vssd1 vccd1 vccd1
+ _02031_ sky130_fd_sc_hd__o22a_1
XANTENNA__10389__A net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09526_ net755 net595 vssd1 vssd1 vccd1 vccd1 _00140_ sky130_fd_sc_hd__and2_1
XFILLER_37_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06738_ top.findLeastValue.val2\[36\] _02412_ top.compVal\[37\] _02485_ vssd1 vssd1
+ vccd1 vccd1 _03526_ sky130_fd_sc_hd__o2bb2a_1
X_09457_ net869 net709 vssd1 vssd1 vccd1 vccd1 _00071_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_42_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08673__A2 top.cb_syn.char_path_n\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09070__D_N top.cb_syn.h_element\[54\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08408_ top.cb_syn.char_path_n\[31\] top.cb_syn.char_path_n\[32\] net515 vssd1 vssd1
+ vccd1 vccd1 _04767_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout431_X net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06669_ _03446_ _03448_ _03452_ _03456_ vssd1 vssd1 vccd1 vccd1 _03457_ sky130_fd_sc_hd__or4b_1
X_09388_ net986 net240 _05268_ _05269_ vssd1 vssd1 vccd1 vccd1 _01443_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_22_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08339_ top.cb_syn.char_path_n\[83\] top.cb_syn.char_path_n\[84\] top.cb_syn.end_cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__mux2_1
X_11350_ clknet_leaf_97_clk _01898_ _00705_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10301_ net798 net638 vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_76_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11281_ clknet_leaf_80_clk net1466 _00636_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_106_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09418__A net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10232_ net829 net669 vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__and2_1
XFILLER_105_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05947__A0 top.WB.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10163_ net827 net667 vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__and2_1
XANTENNA_input37_A gpio_in[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10094_ net834 net674 vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__and2_1
XFILLER_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08361__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10996_ clknet_leaf_29_clk _01544_ _00351_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05478__A2 _02581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11617_ clknet_leaf_64_clk _02165_ _00972_ vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__dfrtp_1
XFILLER_30_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11548_ clknet_leaf_123_clk _02096_ _00903_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[21\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold508 top.sram_interface.word_cnt\[7\] vssd1 vssd1 vccd1 vccd1 net1461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold519 top.histogram.state\[7\] vssd1 vssd1 vccd1 vccd1 net1472 sky130_fd_sc_hd__dlygate4sd3_1
X_11479_ clknet_leaf_101_clk _02027_ _00834_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[19\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_112_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05938__A0 top.WB.CPU_DAT_O\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05971_ top.sram_interface.init_counter\[5\] _02906_ vssd1 vssd1 vccd1 vccd1 _02907_
+ sky130_fd_sc_hd__and2_1
XFILLER_111_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07710_ top.findLeastValue.least2\[0\] top.hTree.tree_reg\[46\] net279 vssd1 vssd1
+ vccd1 vccd1 _04274_ sky130_fd_sc_hd__mux2_1
X_08690_ _04882_ _04885_ _04888_ _04875_ net1675 vssd1 vssd1 vccd1 vccd1 _01486_ sky130_fd_sc_hd__a32o_1
XFILLER_66_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08352__A1 _02506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08378__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07641_ net486 _04215_ vssd1 vssd1 vccd1 vccd1 _04218_ sky130_fd_sc_hd__or2_1
X_07572_ net532 top.cb_syn.h_element\[50\] net539 top.cb_syn.h_element\[59\] _04135_
+ vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_0_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09311_ net432 _05245_ vssd1 vssd1 vccd1 vccd1 _05246_ sky130_fd_sc_hd__or2_1
X_06523_ net1621 _03271_ vssd1 vssd1 vccd1 vccd1 _03315_ sky130_fd_sc_hd__nor2_1
XFILLER_34_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09242_ top.header_synthesis.header\[2\] top.cb_syn.char_index\[2\] net518 vssd1
+ vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__mux2_1
X_06454_ _03269_ _03270_ _03274_ _03276_ top.controller.state_reg\[4\] vssd1 vssd1
+ vccd1 vccd1 _03277_ sky130_fd_sc_hd__o2111a_1
X_05405_ top.cb_syn.zeroes\[3\] vssd1 vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__inv_2
X_09173_ net1696 _05166_ _04821_ vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__a21o_1
XANTENNA__08407__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06385_ _03178_ _03181_ _03227_ vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout224_A _04805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08124_ top.cb_syn.char_path_n\[107\] net196 _04589_ vssd1 vssd1 vccd1 vccd1 _01753_
+ sky130_fd_sc_hd__o21a_1
X_05336_ top.compVal\[5\] vssd1 vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__inv_2
XANTENNA__07030__B top.findLeastValue.val2\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08055_ _04545_ _04547_ top.cb_syn.end_cnt\[5\] vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_112_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09368__B1 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07006_ _03660_ _03661_ _03662_ vssd1 vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__nand3_1
XANTENNA__05641__A2 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05929__A0 top.WB.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07918__B2 top.findLeastValue.sum\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08957_ top.WB.CPU_DAT_O\[16\] top.cb_syn.h_element\[48\] net370 vssd1 vssd1 vccd1
+ vccd1 _01353_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08888_ _02799_ net492 top.findLeastValue.least2\[8\] top.hTree.write_HT_fin vssd1
+ vssd1 vccd1 vccd1 _05058_ sky130_fd_sc_hd__and4b_1
X_07908_ net440 net1579 net251 top.findLeastValue.sum\[7\] _04432_ vssd1 vssd1 vccd1
+ vccd1 _01812_ sky130_fd_sc_hd__a221o_1
X_07839_ top.findLeastValue.sum\[20\] top.hTree.tree_reg\[20\] net285 vssd1 vssd1
+ vccd1 vccd1 _04377_ sky130_fd_sc_hd__mux2_1
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout646_X net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_27_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10850_ clknet_leaf_109_clk _01436_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_55_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07920__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10781_ clknet_leaf_47_clk _01380_ _00200_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09509_ net725 net565 vssd1 vssd1 vccd1 vccd1 _00123_ sky130_fd_sc_hd__and2_1
XFILLER_31_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07854__A0 top.findLeastValue.sum\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_117_Right_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11402_ clknet_leaf_95_clk _01950_ _00757_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[8\]
+ sky130_fd_sc_hd__dfstp_2
X_11333_ clknet_leaf_54_clk _01881_ _00688_ vssd1 vssd1 vccd1 vccd1 top.dut.out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11264_ clknet_leaf_105_clk _01812_ _00619_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10215_ net815 net655 vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__and2_1
X_11195_ clknet_leaf_17_clk _01743_ _00550_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[97\]
+ sky130_fd_sc_hd__dfrtp_2
X_10146_ net825 net665 vssd1 vssd1 vccd1 vccd1 _00760_ sky130_fd_sc_hd__and2_1
X_10077_ net852 net692 vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__and2_1
XANTENNA__08334__A1 top.cb_syn.char_path_n\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05699__A2 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload2_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08926__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07830__S net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10979_ clknet_leaf_10_clk _01527_ _00334_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_99_Left_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07845__A0 top.findLeastValue.sum\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06170_ net549 _02573_ vssd1 vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__nand2_1
Xhold305 top.histogram.sram_out\[15\] vssd1 vssd1 vccd1 vccd1 net1258 sky130_fd_sc_hd__dlygate4sd3_1
Xhold316 top.cb_syn.char_path\[14\] vssd1 vssd1 vccd1 vccd1 net1269 sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 net65 vssd1 vssd1 vccd1 vccd1 net1302 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09058__A net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold338 top.path\[35\] vssd1 vssd1 vccd1 vccd1 net1291 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05623__A2 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold327 top.path\[108\] vssd1 vssd1 vccd1 vccd1 net1280 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout807 net34 vssd1 vssd1 vccd1 vccd1 net807 sky130_fd_sc_hd__buf_4
X_09860_ net771 net611 vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__and2_1
XFILLER_98_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07376__A2 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout818 net819 vssd1 vssd1 vccd1 vccd1 net818 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout829 net835 vssd1 vssd1 vccd1 vccd1 net829 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09791_ net742 net582 vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__and2_1
X_08811_ top.path\[56\] net408 net326 top.path\[57\] net436 vssd1 vssd1 vccd1 vccd1
+ _04994_ sky130_fd_sc_hd__o221a_1
X_05954_ top.WB.CPU_DAT_O\[1\] net1421 net307 vssd1 vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__mux2_1
X_08742_ top.translation.write_fin top.TRN_sram_complete vssd1 vssd1 vccd1 vccd1 _04925_
+ sky130_fd_sc_hd__and2b_1
X_08673_ _02457_ top.cb_syn.char_path_n\[2\] _02935_ _04529_ _04873_ vssd1 vssd1 vccd1
+ vccd1 _04874_ sky130_fd_sc_hd__o2111ai_1
XFILLER_38_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05885_ top.cb_syn.h_element\[52\] top.cb_syn.h_element\[51\] top.cb_syn.h_element\[50\]
+ top.cb_syn.h_element\[53\] vssd1 vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__or4b_1
X_07624_ top.hTree.tree_reg\[62\] top.findLeastValue.least1\[7\] net248 vssd1 vssd1
+ vccd1 vccd1 _04204_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout174_A net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11824__Q top.WB.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07740__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07555_ top.cb_syn.h_element\[61\] top.cb_syn.h_element\[52\] _04145_ vssd1 vssd1
+ vccd1 vccd1 _04146_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout341_A net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07486_ top.cb_syn.char_path_n\[28\] top.cb_syn.char_path_n\[27\] top.cb_syn.char_path_n\[26\]
+ top.cb_syn.char_path_n\[25\] net401 net352 vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__mux4_1
XANTENNA__06356__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06506_ top.histogram.total\[10\] _03308_ net1492 vssd1 vssd1 vccd1 vccd1 _03309_
+ sky130_fd_sc_hd__a21oi_1
X_06437_ _03258_ _03263_ vssd1 vssd1 vccd1 vccd1 _03264_ sky130_fd_sc_hd__and2b_1
X_09225_ net1507 _02540_ _05193_ _05195_ _04913_ vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_write_num_lefts
+ sky130_fd_sc_hd__a41o_1
XANTENNA_fanout606_A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09156_ _05159_ _05160_ _05161_ vssd1 vssd1 vccd1 vccd1 _00043_ sky130_fd_sc_hd__or3_1
X_06368_ top.hist_data_o\[17\] _03185_ vssd1 vssd1 vccd1 vccd1 _03217_ sky130_fd_sc_hd__nor2_1
X_09087_ net295 _05106_ _05107_ _05103_ vssd1 vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__a211o_1
X_06299_ _02494_ _02572_ _02574_ _02458_ net368 vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__a221o_1
XANTENNA__07695__B _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08107_ top.cb_syn.char_path_n\[116\] net375 net335 top.cb_syn.char_path_n\[114\]
+ net180 vssd1 vssd1 vccd1 vccd1 _04581_ sky130_fd_sc_hd__a221o_1
X_05319_ top.compVal\[22\] vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_110_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_110_clk
+ sky130_fd_sc_hd__clkbuf_8
X_08038_ net1507 _02527_ _04532_ vssd1 vssd1 vccd1 vccd1 _01782_ sky130_fd_sc_hd__mux2_1
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10000_ net837 net677 vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__and2_1
X_09989_ net862 net702 vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__and2_1
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11882_ clknet_leaf_39_clk _02398_ _01237_ vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__dfrtp_1
X_10902_ clknet_leaf_39_clk top.header_synthesis.next_header\[7\] _00257_ vssd1 vssd1
+ vccd1 vccd1 top.header_synthesis.header\[7\] sky130_fd_sc_hd__dfrtp_1
X_10833_ clknet_leaf_80_clk _01419_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_10764_ clknet_leaf_47_clk _01363_ _00183_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05550__B2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08047__A top.cb_syn.end_cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10695_ clknet_leaf_113_clk _01294_ _00114_ vssd1 vssd1 vccd1 vccd1 top.path\[71\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08481__S net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05853__A2 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_101_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_101_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11316_ clknet_leaf_76_clk _01864_ _00671_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_10_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05605__A2 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11247_ clknet_leaf_68_clk _01795_ _00602_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.alternator_timer\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_95_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07825__S net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11178_ clknet_leaf_9_clk _01726_ _00533_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[80\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10129_ net838 net678 vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__and2_1
XFILLER_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08656__S net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05670_ top.histogram.sram_out\[2\] net367 net422 top.hTree.node_reg\[2\] _02746_
+ vssd1 vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__a221o_1
XFILLER_35_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_18_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07340_ net270 _03960_ _03961_ net275 net1681 vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_18_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09010_ top.WB.CPU_DAT_O\[15\] net1119 net319 vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__mux2_1
X_07271_ net496 top.findLeastValue.val2\[25\] _03705_ _03910_ vssd1 vssd1 vccd1 vccd1
+ _03911_ sky130_fd_sc_hd__o22a_1
X_06222_ top.cw2\[4\] _03001_ vssd1 vssd1 vccd1 vccd1 _03090_ sky130_fd_sc_hd__or2_1
XANTENNA__05844__A2 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06904__S net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06153_ _02942_ _03019_ _03023_ _02417_ net449 vssd1 vssd1 vccd1 vccd1 _03024_ sky130_fd_sc_hd__a221o_1
Xhold124 top.header_synthesis.header\[6\] vssd1 vssd1 vccd1 vccd1 net1077 sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 top.hTree.tree_reg\[61\] vssd1 vssd1 vccd1 vccd1 net1055 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 top.hTree.node_reg\[30\] vssd1 vssd1 vccd1 vccd1 net1088 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 net73 vssd1 vssd1 vccd1 vccd1 net1066 sky130_fd_sc_hd__dlygate4sd3_1
X_06084_ top.cb_syn.char_index\[1\] top.cb_syn.char_index\[0\] top.cb_syn.char_index\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02957_ sky130_fd_sc_hd__o21a_1
Xhold146 top.hTree.tree_reg\[58\] vssd1 vssd1 vccd1 vccd1 net1099 sky130_fd_sc_hd__dlygate4sd3_1
Xteam_05_909 vssd1 vssd1 vccd1 vccd1 team_05_909/HI gpio_out[24] sky130_fd_sc_hd__conb_1
Xhold168 top.path\[97\] vssd1 vssd1 vccd1 vccd1 net1121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 top.cb_syn.char_path\[74\] vssd1 vssd1 vccd1 vccd1 net1110 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout615 net616 vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__clkbuf_2
Xhold179 top.path\[114\] vssd1 vssd1 vccd1 vccd1 net1132 sky130_fd_sc_hd__dlygate4sd3_1
X_09912_ net759 net599 vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__and2_1
Xfanout604 net607 vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__buf_1
Xfanout626 net647 vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__clkbuf_2
Xfanout637 net640 vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__clkbuf_2
XFILLER_98_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09843_ net761 net601 vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__and2_1
XANTENNA__07735__S net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout648 net651 vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__clkbuf_2
XFILLER_112_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout389_A net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06859__B net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout659 net664 vssd1 vssd1 vccd1 vccd1 net659 sky130_fd_sc_hd__clkbuf_2
XANTENNA__05763__B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09774_ net789 net629 vssd1 vssd1 vccd1 vccd1 _00388_ sky130_fd_sc_hd__and2_1
X_06986_ top.findLeastValue.val1\[6\] top.findLeastValue.val1\[5\] top.findLeastValue.val1\[4\]
+ top.findLeastValue.val1\[3\] vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout177_X net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08725_ _04899_ _04905_ _04911_ _04898_ top.cb_syn.i\[1\] vssd1 vssd1 vccd1 vccd1
+ _01474_ sky130_fd_sc_hd__a32o_1
X_05937_ top.WB.CPU_DAT_O\[18\] net1311 net304 vssd1 vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__mux2_1
X_05868_ top.sram_interface.init_counter\[15\] top.sram_interface.init_counter\[14\]
+ top.sram_interface.init_counter\[13\] top.sram_interface.init_counter\[12\] vssd1
+ vssd1 vccd1 vccd1 _02847_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_107_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ top.cb_syn.cb_length\[1\] _04861_ net210 vssd1 vssd1 vccd1 vccd1 _01493_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08566__S net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_54_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08587_ _04812_ top.cb_syn.char_index\[3\] _04807_ vssd1 vssd1 vccd1 vccd1 _01513_
+ sky130_fd_sc_hd__mux2_1
XFILLER_81_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07607_ net445 _04188_ vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__nor2_1
X_07538_ top.cb_syn.pulse_first _02872_ vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__or2_1
XANTENNA__05532__B2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05799_ top.WorR _02529_ _02807_ _02815_ vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__or4_1
X_07469_ _04050_ _04059_ _04051_ vssd1 vssd1 vccd1 vccd1 _04060_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout511_X net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_69_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09208_ net517 _02930_ vssd1 vssd1 vccd1 vccd1 _05184_ sky130_fd_sc_hd__nor2_1
X_10480_ net861 net701 vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__and2_1
XFILLER_10_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09139_ net548 net468 _02548_ _05149_ vssd1 vssd1 vccd1 vccd1 _05150_ sky130_fd_sc_hd__a31o_1
XANTENNA_clkbuf_leaf_112_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06245__C1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06115__A top.cb_syn.char_index\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11101_ clknet_leaf_13_clk _01649_ _00456_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__06796__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold680 top.translation.write_fin vssd1 vssd1 vccd1 vccd1 net1633 sky130_fd_sc_hd__dlygate4sd3_1
Xhold691 top.header_synthesis.count\[6\] vssd1 vssd1 vccd1 vccd1 net1644 sky130_fd_sc_hd__dlygate4sd3_1
X_11032_ clknet_leaf_42_clk _01580_ _00387_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_92_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11865_ clknet_leaf_115_clk _02381_ _01220_ vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__dfrtp_1
X_11796_ clknet_leaf_58_clk _00014_ _01151_ vssd1 vssd1 vccd1 vccd1 top.controller.state_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_15_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10816_ clknet_leaf_109_clk _01402_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_10747_ clknet_leaf_120_clk _01346_ _00166_ vssd1 vssd1 vccd1 vccd1 top.path\[123\]
+ sky130_fd_sc_hd__dfrtp_1
X_10678_ clknet_leaf_123_clk _01277_ _00097_ vssd1 vssd1 vccd1 vccd1 top.path\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08776__A1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__06787__B1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06840_ _02475_ net152 net126 _03559_ vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__a2bb2o_1
X_06771_ net504 net412 net119 net134 top.cw1\[0\] vssd1 vssd1 vccd1 vccd1 _02065_
+ sky130_fd_sc_hd__a32o_1
XANTENNA__05762__B2 top.WB.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05722_ top.TRN_char_index\[5\] net43 net720 vssd1 vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__mux2_1
X_08510_ net1083 top.cb_syn.char_path_n\[66\] net227 vssd1 vssd1 vccd1 vccd1 _01584_
+ sky130_fd_sc_hd__mux2_1
X_09490_ net733 net573 vssd1 vssd1 vccd1 vccd1 _00104_ sky130_fd_sc_hd__and2_1
XANTENNA__08161__C1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08441_ top.cb_syn.end_cnt\[6\] _04722_ _04748_ _04775_ _04799_ vssd1 vssd1 vccd1
+ vccd1 _04800_ sky130_fd_sc_hd__a32oi_4
X_05653_ net1283 net145 _02732_ net177 vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_34_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05514__B2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08372_ _02505_ _04723_ _04726_ net506 vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__o211a_1
X_05584_ net457 top.hTree.node_reg\[48\] net361 net420 top.hTree.node_reg\[16\] vssd1
+ vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_102_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07323_ top.findLeastValue.sum\[14\] net274 net269 _03949_ vssd1 vssd1 vccd1 vccd1
+ _01910_ sky130_fd_sc_hd__a22o_1
X_07254_ _03809_ _03816_ vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__and2_1
X_06205_ top.sram_interface.init_counter\[4\] _02944_ top.sram_interface.init_counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03074_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_57_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07185_ top.findLeastValue.val1\[41\] top.findLeastValue.val2\[41\] vssd1 vssd1 vccd1
+ vccd1 _03843_ sky130_fd_sc_hd__nor2_1
X_06136_ _02579_ _02984_ _03007_ net469 _02990_ vssd1 vssd1 vccd1 vccd1 _03008_ sky130_fd_sc_hd__a221o_1
XANTENNA__06778__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06067_ net495 _02851_ vssd1 vssd1 vccd1 vccd1 _02942_ sky130_fd_sc_hd__and2_2
XFILLER_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06196__A2_N _02767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout401 net402 vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__buf_4
Xfanout412 net413 vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__buf_2
Xfanout423 net424 vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__clkbuf_4
XANTENNA__05774__A top.findLeastValue.least1\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout294_X net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout456 net458 vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__buf_2
Xfanout445 net448 vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__clkbuf_4
Xfanout434 net435 vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__buf_2
XANTENNA__07727__C1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout467 top.controller.state_reg\[4\] vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__buf_1
Xfanout478 net479 vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__buf_2
Xfanout489 net492 vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__buf_2
X_09826_ net768 net608 vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__and2_1
XFILLER_104_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07742__A2 _04298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09757_ net739 net579 vssd1 vssd1 vccd1 vccd1 _00371_ sky130_fd_sc_hd__and2_1
X_06969_ top.findLeastValue.val2\[14\] top.findLeastValue.val2\[13\] top.findLeastValue.val2\[12\]
+ top.findLeastValue.val2\[11\] vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__and4_1
X_08708_ top.cb_syn.i\[3\] top.cb_syn.i\[2\] top.cb_syn.i\[1\] top.cb_syn.i\[0\] vssd1
+ vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout559_X net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05753__B2 top.WB.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09688_ net785 net625 vssd1 vssd1 vccd1 vccd1 _00302_ sky130_fd_sc_hd__and2_1
X_08639_ net210 _04849_ vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__nand2_1
XANTENNA__09131__D net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11650_ clknet_leaf_112_clk _02183_ _01005_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11581_ clknet_leaf_108_clk _02129_ _00936_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10601_ net752 net592 vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_12_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10532_ net858 net698 vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__and2_1
XFILLER_6_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10463_ net723 net563 vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_79_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10394_ net763 net603 vssd1 vssd1 vccd1 vccd1 _01008_ sky130_fd_sc_hd__and2_1
X_11015_ clknet_leaf_4_clk _01563_ _00370_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_64_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08391__C1 _02504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06941__B1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08143__C1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08694__B1 _04875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11848_ clknet_leaf_116_clk _02364_ _01203_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[26\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_33_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11779_ clknet_leaf_73_clk _02312_ _01134_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.counter_HTREE\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload11 clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clkload11/X sky130_fd_sc_hd__clkbuf_8
Xclkload44 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 clkload44/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload33 clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 clkload33/X sky130_fd_sc_hd__clkbuf_4
Xclkload22 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 clkload22/Y sky130_fd_sc_hd__clkinv_2
Xclkload66 clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 clkload66/Y sky130_fd_sc_hd__inv_6
Xclkload55 clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 clkload55/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__09410__A2 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload77 clknet_leaf_80_clk vssd1 vssd1 vccd1 vccd1 clkload77/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__11369__Q top.findLeastValue.sum\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload99 clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 clkload99/Y sky130_fd_sc_hd__inv_6
Xclkload88 clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 clkload88/X sky130_fd_sc_hd__clkbuf_4
X_08990_ top.WB.CPU_DAT_O\[2\] net1289 net324 vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__mux2_1
X_07941_ net488 _04457_ vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__or2_1
X_07872_ net426 _04402_ _04403_ net261 vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__o211a_1
X_09611_ net851 net691 vssd1 vssd1 vccd1 vccd1 _00225_ sky130_fd_sc_hd__and2_1
XANTENNA__08382__C1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06823_ top.findLeastValue.val1\[7\] net130 net114 top.compVal\[7\] vssd1 vssd1 vccd1
+ vccd1 _02015_ sky130_fd_sc_hd__o22a_1
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_09542_ net746 net586 vssd1 vssd1 vccd1 vccd1 _00156_ sky130_fd_sc_hd__and2_1
X_06754_ _03527_ _03541_ _03526_ vssd1 vssd1 vccd1 vccd1 _03542_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_104_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05705_ net8 net415 net308 top.WB.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 _02353_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07314__A _03782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout254_A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11832__Q top.WB.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06685_ _02439_ top.findLeastValue.val2\[10\] top.findLeastValue.val2\[9\] _02440_
+ vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__a22o_1
X_09473_ net750 net590 vssd1 vssd1 vccd1 vccd1 _00087_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_90_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_90_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__06160__A1 top.cb_syn.char_index\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05499__B1 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08424_ net515 top.cb_syn.char_path_n\[55\] vssd1 vssd1 vccd1 vccd1 _04783_ sky130_fd_sc_hd__or2_1
X_05636_ top.cb_syn.char_path\[71\] net552 net542 top.cb_syn.char_path\[39\] vssd1
+ vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__a22o_1
X_08355_ net512 _04696_ _04713_ vssd1 vssd1 vccd1 vccd1 _04714_ sky130_fd_sc_hd__a21oi_1
X_05567_ top.histogram.sram_out\[19\] net364 _02659_ _02660_ vssd1 vssd1 vccd1 vccd1
+ _02661_ sky130_fd_sc_hd__a211o_1
Xclkload5 clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clkload5/X sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout421_A net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07306_ _03792_ _03936_ vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__nand2_1
X_05498_ top.cb_syn.char_path\[30\] net559 net314 top.cb_syn.char_path\[126\] vssd1
+ vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__a22o_1
X_08286_ top.cb_syn.char_path_n\[26\] net206 _04670_ vssd1 vssd1 vccd1 vccd1 _01672_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__06364__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07660__B2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07237_ _03671_ _03832_ _03836_ vssd1 vssd1 vccd1 vccd1 _03886_ sky130_fd_sc_hd__nand3_1
XANTENNA_fanout790_A net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07168_ _02466_ _02486_ vssd1 vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_115_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06119_ top.cw1\[1\] top.cw1\[0\] vssd1 vssd1 vccd1 vccd1 _02991_ sky130_fd_sc_hd__nand2_1
XFILLER_3_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06766__A3 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07099_ _03754_ _03755_ _03748_ vssd1 vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__a21o_1
XANTENNA__09165__A1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout231 net235 vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__clkbuf_4
Xfanout220 net221 vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__clkbuf_4
XFILLER_115_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout264 net266 vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__buf_2
Xfanout253 net256 vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__clkbuf_4
Xfanout242 net243 vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__buf_2
XFILLER_115_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout297 _03998_ vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__buf_2
XFILLER_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08373__C1 _02504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09809_ net787 net627 vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__and2_1
Xfanout286 _04197_ vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__clkbuf_4
Xfanout275 net277 vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__buf_2
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ clknet_leaf_115_clk _02235_ _01057_ vssd1 vssd1 vccd1 vccd1 top.path\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08754__S net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_81_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_clk sky130_fd_sc_hd__clkbuf_8
X_11633_ clknet_leaf_55_clk top.dut.bit_buf_next\[5\] _00988_ vssd1 vssd1 vccd1 vccd1
+ top.dut.bit_buf\[5\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__08607__X _04826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11564_ clknet_leaf_37_clk _02112_ _00919_ vssd1 vssd1 vccd1 vccd1 top.header_synthesis.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10515_ net868 net708 vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__and2_1
XANTENNA__07651__A1 top.findLeastValue.least1\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06454__A2 _03270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11495_ clknet_leaf_87_clk _02043_ _00850_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[35\]
+ sky130_fd_sc_hd__dfstp_1
X_10446_ net748 net588 vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__and2_1
XANTENNA__05685__Y _02759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10377_ net855 net695 vssd1 vssd1 vccd1 vccd1 _00991_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_90_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08929__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05717__B2 top.WB.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_72_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_clk sky130_fd_sc_hd__clkbuf_8
X_06470_ top.histogram.total\[30\] _03292_ vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__nand2_1
X_05421_ net556 vssd1 vssd1 vccd1 vccd1 _02529_ sky130_fd_sc_hd__inv_2
X_08140_ top.cb_syn.char_path_n\[99\] net201 _04597_ vssd1 vssd1 vccd1 vccd1 _01745_
+ sky130_fd_sc_hd__o21a_1
XFILLER_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05352_ top.findLeastValue.val1\[44\] vssd1 vssd1 vccd1 vccd1 _02460_ sky130_fd_sc_hd__inv_2
X_08071_ top.cb_syn.wait_cycle net540 _02553_ _02862_ vssd1 vssd1 vccd1 vccd1 _04558_
+ sky130_fd_sc_hd__a22o_1
Xclkload122 clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 clkload122/Y sky130_fd_sc_hd__inv_6
Xclkload111 clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 clkload111/Y sky130_fd_sc_hd__clkinv_4
Xclkload100 clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 clkload100/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__07642__A1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07642__B2 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__05653__B1 _02732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06912__S net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07022_ top.findLeastValue.val1\[26\] top.findLeastValue.val2\[26\] vssd1 vssd1 vccd1
+ vccd1 _03680_ sky130_fd_sc_hd__or2_1
XANTENNA__11827__Q top.WB.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08973_ top.WB.CPU_DAT_O\[19\] net1275 net324 vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__mux2_1
Xhold17 top.sram_interface.init_counter\[14\] vssd1 vssd1 vccd1 vccd1 net970 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 top.hTree.node_reg\[54\] vssd1 vssd1 vccd1 vccd1 net981 sky130_fd_sc_hd__dlygate4sd3_1
X_07924_ top.findLeastValue.sum\[3\] top.hTree.tree_reg\[3\] net282 vssd1 vssd1 vccd1
+ vccd1 _04445_ sky130_fd_sc_hd__mux2_1
XANTENNA__07028__B top.findLeastValue.val2\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold39 top.hTree.node_reg\[47\] vssd1 vssd1 vccd1 vccd1 net992 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout371_A net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08370__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07855_ top.findLeastValue.sum\[17\] _04389_ net395 vssd1 vssd1 vccd1 vccd1 _04390_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__05708__B2 top.WB.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06905__B1 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_119_Left_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06359__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07786_ net489 _04333_ vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__or2_1
XFILLER_43_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06806_ top.findLeastValue.val1\[24\] net132 net116 top.compVal\[24\] vssd1 vssd1
+ vccd1 vccd1 _02032_ sky130_fd_sc_hd__o22a_1
XANTENNA__08658__B1 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09525_ net755 net595 vssd1 vssd1 vccd1 vccd1 _00139_ sky130_fd_sc_hd__and2_1
X_06737_ _03505_ _03524_ _03514_ vssd1 vssd1 vccd1 vccd1 _03525_ sky130_fd_sc_hd__o21ba_1
XFILLER_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09456_ net869 net709 vssd1 vssd1 vccd1 vccd1 _00070_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_63_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout636_A net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout257_X net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08574__S net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06668_ top.compVal\[40\] _02484_ _03445_ _03447_ vssd1 vssd1 vccd1 vccd1 _03456_
+ sky130_fd_sc_hd__o211a_1
XFILLER_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08407_ top.cb_syn.char_path_n\[25\] net392 _04765_ vssd1 vssd1 vccd1 vccd1 _04766_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05619_ top.cb_syn.char_path\[10\] net557 net312 top.cb_syn.char_path\[106\] vssd1
+ vssd1 vccd1 vccd1 _02704_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout424_X net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09387_ top.hTree.nulls\[49\] net405 net244 vssd1 vssd1 vccd1 vccd1 _05269_ sky130_fd_sc_hd__o21a_1
X_06599_ _03327_ _03338_ _03382_ _03387_ vssd1 vssd1 vccd1 vccd1 _03388_ sky130_fd_sc_hd__a2bb2o_2
X_08338_ net512 _02506_ vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_22_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08269_ top.cb_syn.char_path_n\[35\] net381 net339 top.cb_syn.char_path_n\[33\] net185
+ vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__a221o_1
X_10300_ net799 net639 vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__and2_1
X_11280_ clknet_leaf_77_clk _01828_ _00635_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_106_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10231_ net821 net661 vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__and2_1
XANTENNA__11737__Q top.CB_write_complete vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07492__S0 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10162_ net817 net657 vssd1 vssd1 vccd1 vccd1 _00776_ sky130_fd_sc_hd__and2_1
X_10093_ net834 net674 vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__and2_1
XFILLER_101_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_54_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_87_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10995_ clknet_leaf_24_clk _01543_ _00350_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08744__S0 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08484__S net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07321__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11616_ clknet_leaf_63_clk _02164_ _00971_ vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07624__A1 top.findLeastValue.least1\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11547_ clknet_leaf_123_clk _02095_ _00902_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[20\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold509 top.histogram.total\[24\] vssd1 vssd1 vccd1 vccd1 net1462 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05635__B1 _02717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11478_ clknet_leaf_101_clk _02026_ _00833_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[18\]
+ sky130_fd_sc_hd__dfstp_1
X_10429_ net875 net715 vssd1 vssd1 vccd1 vccd1 _01043_ sky130_fd_sc_hd__and2_1
XANTENNA__09377__B2 _04278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05970_ top.sram_interface.init_counter\[4\] top.sram_interface.init_counter\[3\]
+ _02905_ vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__and3_1
XANTENNA__06060__B1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07640_ net486 _04216_ vssd1 vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__nand2_1
X_07571_ top.cb_syn.h_element\[59\] top.cb_syn.h_element\[50\] _04145_ vssd1 vssd1
+ vccd1 vccd1 _04160_ sky130_fd_sc_hd__mux2_1
XFILLER_80_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_45_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_clk sky130_fd_sc_hd__clkbuf_8
X_09310_ top.histogram.total\[18\] top.histogram.total\[19\] net524 vssd1 vssd1 vccd1
+ vccd1 _05245_ sky130_fd_sc_hd__mux2_1
X_06522_ net1560 _03272_ vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__xor2_1
X_09241_ net1057 _05205_ net296 vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_header\[1\]
+ sky130_fd_sc_hd__mux2_1
X_06453_ top.histogram.total\[5\] top.histogram.total\[4\] vssd1 vssd1 vccd1 vccd1
+ _03276_ sky130_fd_sc_hd__and2_1
XANTENNA__07863__A1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05404_ top.cb_syn.zeroes\[4\] vssd1 vssd1 vccd1 vccd1 _02512_ sky130_fd_sc_hd__inv_2
X_09172_ top.cb_syn.setup net475 _02932_ vssd1 vssd1 vccd1 vccd1 _05166_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_60_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06384_ top.hist_data_o\[11\] _03180_ vssd1 vssd1 vccd1 vccd1 _03227_ sky130_fd_sc_hd__nor2_1
XFILLER_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05335_ top.compVal\[6\] vssd1 vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__inv_2
X_08123_ top.cb_syn.char_path_n\[108\] net377 net334 top.cb_syn.char_path_n\[106\]
+ net179 vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__a221o_1
X_08054_ net535 net246 _04541_ vssd1 vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout217_A net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07005_ _03661_ _03662_ vssd1 vssd1 vccd1 vccd1 _03663_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_112_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09368__B2 _04314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08040__A1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08956_ top.WB.CPU_DAT_O\[17\] top.cb_syn.h_element\[49\] net369 vssd1 vssd1 vccd1
+ vccd1 _01354_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07907_ net425 _04430_ _04431_ net258 vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__o211a_1
X_08887_ _02519_ _02785_ net1650 vssd1 vssd1 vccd1 vccd1 _01458_ sky130_fd_sc_hd__o21a_1
X_07838_ net445 net1440 net253 top.findLeastValue.sum\[21\] _04376_ vssd1 vssd1 vccd1
+ vccd1 _01826_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_27_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_36_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout541_X net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07769_ top.findLeastValue.sum\[34\] top.hTree.tree_reg\[34\] net280 vssd1 vssd1
+ vccd1 vccd1 _04321_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09508_ net758 net598 vssd1 vssd1 vccd1 vccd1 _00122_ sky130_fd_sc_hd__and2_1
X_10780_ clknet_leaf_79_clk _01379_ _00199_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout806_X net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09439_ net973 vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__clkbuf_1
XFILLER_52_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11401_ clknet_leaf_95_clk _01949_ _00756_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[7\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__05617__B1 _02702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11332_ clknet_leaf_54_clk _01880_ _00687_ vssd1 vssd1 vccd1 vccd1 top.dut.out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11263_ clknet_leaf_106_clk _01811_ _00618_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11194_ clknet_leaf_18_clk _01742_ _00549_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[96\]
+ sky130_fd_sc_hd__dfrtp_2
X_10214_ net815 net655 vssd1 vssd1 vccd1 vccd1 _00828_ sky130_fd_sc_hd__and2_1
XANTENNA__06042__B1 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10145_ net825 net665 vssd1 vssd1 vccd1 vccd1 _00759_ sky130_fd_sc_hd__and2_1
XFILLER_79_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08479__S net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10076_ net853 net693 vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_89_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08334__A2 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_27_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_90_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10978_ clknet_leaf_11_clk _01526_ _00333_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold306 top.histogram.sram_out\[27\] vssd1 vssd1 vccd1 vccd1 net1259 sky130_fd_sc_hd__dlygate4sd3_1
Xhold317 net78 vssd1 vssd1 vccd1 vccd1 net1270 sky130_fd_sc_hd__dlygate4sd3_1
Xhold339 top.hTree.nulls\[57\] vssd1 vssd1 vccd1 vccd1 net1292 sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 top.cb_syn.char_path\[81\] vssd1 vssd1 vccd1 vccd1 net1281 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout819 net824 vssd1 vssd1 vccd1 vccd1 net819 sky130_fd_sc_hd__clkbuf_2
X_08810_ net432 _04992_ vssd1 vssd1 vccd1 vccd1 _04993_ sky130_fd_sc_hd__or2_1
Xfanout808 net811 vssd1 vssd1 vccd1 vccd1 net808 sky130_fd_sc_hd__clkbuf_2
X_09790_ net742 net582 vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__and2_1
X_08741_ _04924_ _04916_ top.header_synthesis.bit1 _04923_ vssd1 vssd1 vccd1 vccd1
+ _01471_ sky130_fd_sc_hd__o2bb2a_1
X_05953_ top.WB.CPU_DAT_O\[2\] net1415 net307 vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__mux2_1
X_08672_ net530 net536 net529 net538 vssd1 vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__or4_1
X_05884_ top.cb_syn.h_element\[49\] top.cb_syn.h_element\[48\] top.cb_syn.h_element\[47\]
+ top.cb_syn.h_element\[46\] vssd1 vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__or4_1
XANTENNA__10013__A net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07623_ top.findLeastValue.least1\[7\] top.hTree.tree_reg\[62\] net279 vssd1 vssd1
+ vccd1 vccd1 _04203_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_18_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout167_A _03423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06887__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07554_ _04121_ top.cb_syn.h_element\[63\] vssd1 vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__nand2b_4
X_07485_ top.cb_syn.char_path_n\[24\] top.cb_syn.char_path_n\[23\] top.cb_syn.char_path_n\[22\]
+ top.cb_syn.char_path_n\[21\] net401 net352 vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_52_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11840__Q top.WB.CPU_DAT_O\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06505_ top.histogram.total\[9\] top.histogram.total\[8\] _03279_ vssd1 vssd1 vccd1
+ vccd1 _03308_ sky130_fd_sc_hd__and3_1
X_06436_ _03261_ _03262_ _03246_ vssd1 vssd1 vccd1 vccd1 _03263_ sky130_fd_sc_hd__a21bo_1
X_09224_ top.cb_syn.num_lefts\[7\] top.cb_syn.num_lefts\[6\] _04843_ _05194_ vssd1
+ vssd1 vccd1 vccd1 _05195_ sky130_fd_sc_hd__or4_1
XANTENNA__05847__B1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09155_ net451 net459 net562 _02556_ vssd1 vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__a31o_1
X_06367_ net1272 net301 _03216_ vssd1 vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout122_X net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06298_ net1302 net143 _03162_ net159 vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__a22o_1
X_09086_ top.histogram.out_of_init top.histogram.eof_n _02534_ net295 vssd1 vssd1
+ vccd1 vccd1 _05107_ sky130_fd_sc_hd__and4b_1
X_08106_ top.cb_syn.char_path_n\[116\] net204 _04580_ vssd1 vssd1 vccd1 vccd1 _01762_
+ sky130_fd_sc_hd__o21a_1
X_05318_ top.compVal\[23\] vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__inv_2
XFILLER_107_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08037_ net540 net529 _02871_ _04478_ _04531_ vssd1 vssd1 vccd1 vccd1 _04532_ sky130_fd_sc_hd__o221a_1
XANTENNA__06272__B1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06811__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout870_A net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07367__A3 _03547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09210__B1 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09988_ net864 net704 vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__and2_1
X_08939_ top.WB.CPU_DAT_O\[15\] net1356 net371 vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__mux2_1
XANTENNA__06401__A net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout756_X net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08316__A2 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10901_ clknet_leaf_39_clk top.header_synthesis.next_header\[6\] _00256_ vssd1 vssd1
+ vccd1 vccd1 top.header_synthesis.header\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_44_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11881_ clknet_leaf_39_clk _02397_ _01236_ vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__dfrtp_1
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05774__D_N top.findLeastValue.least1\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10832_ clknet_leaf_79_clk _01418_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05550__A2 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10763_ clknet_leaf_47_clk _01362_ _00182_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08047__B net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05838__B1 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10694_ clknet_leaf_113_clk _01293_ _00113_ vssd1 vssd1 vccd1 vccd1 top.path\[70\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05687__A net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08788__C1 top.translation.index\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11315_ clknet_leaf_71_clk _01863_ _00670_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_10_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06802__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11246_ clknet_leaf_68_clk _01794_ _00601_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.alternator_timer\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11177_ clknet_leaf_8_clk _01725_ _00532_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[79\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07763__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10128_ net842 net682 vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__and2_1
X_10059_ net845 net685 vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__and2_1
XFILLER_63_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07818__A1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_07270_ _03684_ _03898_ vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__nor2_1
X_06221_ top.findLeastValue.histo_index\[3\] _02767_ _03013_ _03088_ vssd1 vssd1 vccd1
+ vccd1 _03089_ sky130_fd_sc_hd__o2bb2a_1
X_06152_ top.hist_addr\[6\] _03022_ vssd1 vssd1 vccd1 vccd1 _03023_ sky130_fd_sc_hd__nand2_1
XFILLER_8_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_06083_ top.cb_syn.char_index\[2\] top.cb_syn.char_index\[1\] vssd1 vssd1 vccd1 vccd1
+ _02956_ sky130_fd_sc_hd__nand2_1
Xhold125 top.cb_syn.char_path\[59\] vssd1 vssd1 vccd1 vccd1 net1078 sky130_fd_sc_hd__dlygate4sd3_1
Xhold103 top.hTree.node_reg\[28\] vssd1 vssd1 vccd1 vccd1 net1056 sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 top.path\[15\] vssd1 vssd1 vccd1 vccd1 net1067 sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 top.sram_interface.init_counter\[11\] vssd1 vssd1 vccd1 vccd1 net1100 sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 top.cb_syn.char_path\[95\] vssd1 vssd1 vccd1 vccd1 net1111 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_8
X_09911_ net759 net599 vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__and2_1
Xhold136 top.path\[26\] vssd1 vssd1 vccd1 vccd1 net1089 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08701__A top.cb_syn.h_element\[63\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold169 net90 vssd1 vssd1 vccd1 vccd1 net1122 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout605 net606 vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06920__S net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout638 net639 vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__clkbuf_2
XFILLER_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout616 net647 vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__clkbuf_2
Xfanout627 net631 vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__clkbuf_2
X_09842_ net760 net600 vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__and2_1
Xfanout649 net651 vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__buf_1
X_09773_ net789 net629 vssd1 vssd1 vccd1 vccd1 _00387_ sky130_fd_sc_hd__and2_1
XANTENNA__06859__C net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08724_ top.cb_syn.i\[1\] top.cb_syn.i\[0\] vssd1 vssd1 vccd1 vccd1 _04911_ sky130_fd_sc_hd__or2_1
XANTENNA__11835__Q top.WB.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06985_ top.findLeastValue.val1\[14\] top.findLeastValue.val1\[13\] top.findLeastValue.val1\[12\]
+ top.findLeastValue.val1\[11\] vssd1 vssd1 vccd1 vccd1 _03643_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout284_A _04197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_7_0_clk_X clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05936_ top.WB.CPU_DAT_O\[19\] net1265 net304 vssd1 vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__mux2_1
XFILLER_26_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08655_ _04858_ _04860_ vssd1 vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__nor2_1
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05867_ net1731 net170 net156 top.WB.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 _02275_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09532__A net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08586_ top.cb_syn.h_element\[58\] top.cb_syn.h_element\[49\] net532 vssd1 vssd1
+ vccd1 vccd1 _04812_ sky130_fd_sc_hd__mux2_1
X_07606_ net458 _04188_ vssd1 vssd1 vccd1 vccd1 _04190_ sky130_fd_sc_hd__nand2_1
XFILLER_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07537_ top.cb_syn.h_element\[63\] _04122_ _04127_ vssd1 vssd1 vccd1 vccd1 _04128_
+ sky130_fd_sc_hd__and3_1
XANTENNA__05532__A2 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05798_ _02803_ _02812_ _02814_ _02817_ vssd1 vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__or4_1
XANTENNA__11570__Q top.histogram.sram_out\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout716_A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07468_ _04054_ _04058_ _04052_ vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__a21oi_4
X_06419_ top.header_synthesis.count\[6\] _03249_ _03246_ vssd1 vssd1 vccd1 vccd1 _03250_
+ sky130_fd_sc_hd__a21oi_1
X_07399_ top.dut.bits_in_buf_next\[2\] net297 vssd1 vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__nor2_1
X_09207_ net529 net474 _05182_ _05183_ vssd1 vssd1 vccd1 vccd1 _00011_ sky130_fd_sc_hd__o22a_1
XFILLER_108_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09138_ top.WorR net548 top.hTree.write_HT_fin net461 vssd1 vssd1 vccd1 vccd1 _05149_
+ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_118_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10914__Q top.header_synthesis.enable vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09069_ net517 net474 _02931_ _05092_ vssd1 vssd1 vccd1 vccd1 _05093_ sky130_fd_sc_hd__a31o_1
X_11100_ clknet_leaf_17_clk _01648_ _00455_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__05599__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold670 top.dut.out\[1\] vssd1 vssd1 vccd1 vccd1 net1623 sky130_fd_sc_hd__dlygate4sd3_1
Xhold681 top.cb_syn.cb_length\[0\] vssd1 vssd1 vccd1 vccd1 net1634 sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 top.cb_syn.cb_length\[6\] vssd1 vssd1 vccd1 vccd1 net1645 sky130_fd_sc_hd__dlygate4sd3_1
X_11031_ clknet_leaf_42_clk _01579_ _00386_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[61\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11972__A net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input12_A DAT_I[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11864_ clknet_leaf_116_clk _02380_ _01219_ vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__dfrtp_1
XANTENNA__06181__C1 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08058__A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10815_ clknet_leaf_105_clk _01401_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_11795_ clknet_leaf_58_clk net1590 _01150_ vssd1 vssd1 vccd1 vccd1 top.controller.state_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08492__S net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10746_ clknet_leaf_120_clk _01345_ _00165_ vssd1 vssd1 vccd1 vccd1 top.path\[122\]
+ sky130_fd_sc_hd__dfrtp_1
X_10677_ clknet_leaf_0_clk _01276_ _00096_ vssd1 vssd1 vccd1 vccd1 top.path\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11229_ clknet_leaf_27_clk _01777_ _00584_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.end_cnt\[2\]
+ sky130_fd_sc_hd__dfstp_1
X_06770_ net1501 net412 net119 net134 top.cw1\[1\] vssd1 vssd1 vccd1 vccd1 _02066_
+ sky130_fd_sc_hd__a32o_1
X_05721_ top.TRN_char_index\[6\] net35 net720 vssd1 vssd1 vccd1 vccd1 _02337_ sky130_fd_sc_hd__mux2_1
X_08440_ top.cb_syn.end_cnt\[5\] _04798_ top.cb_syn.end_cnt\[6\] vssd1 vssd1 vccd1
+ vccd1 _04799_ sky130_fd_sc_hd__a21oi_1
X_05652_ top.histogram.sram_out\[5\] net364 net419 top.hTree.node_reg\[5\] _02731_
+ vssd1 vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_34_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05514__A2 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08371_ top.cb_syn.char_path_n\[113\] top.cb_syn.char_path_n\[114\] top.cb_syn.char_path_n\[115\]
+ top.cb_syn.char_path_n\[116\] net514 net510 vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__mux4_1
X_05583_ _02672_ _02673_ net472 vssd1 vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_102_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07322_ _03714_ _03945_ vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07253_ net1710 net277 net272 _03897_ vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__a22o_1
X_06204_ _03022_ _03072_ vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__nor2_1
X_07184_ _03840_ _03841_ vssd1 vssd1 vccd1 vccd1 _03842_ sky130_fd_sc_hd__nand2_1
X_06135_ top.cw2\[7\] _02572_ _03005_ _03006_ vssd1 vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_57_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06778__A1 top.findLeastValue.least1\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06066_ net1029 net141 net137 vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__a21o_1
Xfanout402 _04074_ vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__clkbuf_4
Xfanout413 net414 vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__clkbuf_2
Xfanout424 _02537_ vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__buf_2
XFILLER_86_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xfanout457 net458 vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__clkbuf_4
X_09825_ net768 net608 vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__and2_1
Xfanout446 net447 vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__buf_2
Xfanout435 _02524_ vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__buf_2
XANTENNA_input4_A DAT_I[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout479 net481 vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__buf_2
Xfanout468 net469 vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__buf_2
XANTENNA_fanout287_X net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout666_A net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06968_ top.findLeastValue.val2\[10\] top.findLeastValue.val2\[9\] top.findLeastValue.val2\[8\]
+ top.findLeastValue.val2\[7\] vssd1 vssd1 vccd1 vccd1 _03626_ sky130_fd_sc_hd__and4_1
X_09756_ net736 net576 vssd1 vssd1 vccd1 vccd1 _00370_ sky130_fd_sc_hd__and2_1
X_09687_ net784 net624 vssd1 vssd1 vccd1 vccd1 _00301_ sky130_fd_sc_hd__and2_1
X_08707_ top.cb_syn.i\[1\] top.cb_syn.i\[0\] vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__nand2_1
XFILLER_100_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05919_ net550 net465 vssd1 vssd1 vccd1 vccd1 _02889_ sky130_fd_sc_hd__nand2_1
XFILLER_67_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout454_X net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08638_ _04848_ _04846_ top.cb_syn.cb_length\[4\] vssd1 vssd1 vccd1 vccd1 _04849_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06899_ top.findLeastValue.val2\[34\] net150 net125 _03591_ vssd1 vssd1 vccd1 vccd1
+ _01976_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout719_X net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08569_ net1165 top.cb_syn.char_path_n\[7\] net225 vssd1 vssd1 vccd1 vccd1 _01525_
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10600_ net808 net648 vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_12_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11580_ clknet_leaf_108_clk _02128_ _00935_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10531_ net859 net699 vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__and2_1
X_10462_ net723 net563 vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_79_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10393_ net763 net603 vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__and2_1
XFILLER_108_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_92_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11014_ clknet_leaf_4_clk _01562_ _00369_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07718__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08391__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_11847_ clknet_leaf_116_clk _02363_ _01202_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[25\]
+ sky130_fd_sc_hd__dfrtp_4
X_11778_ clknet_leaf_50_clk net961 _01133_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.CB_read_counter
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10729_ clknet_leaf_118_clk _01328_ _00148_ vssd1 vssd1 vccd1 vccd1 top.path\[105\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload12 clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clkload12/X sky130_fd_sc_hd__clkbuf_8
XFILLER_70_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload34 clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 clkload34/Y sky130_fd_sc_hd__inv_6
Xclkload23 clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 clkload23/Y sky130_fd_sc_hd__clkinv_2
Xclkload67 clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 clkload67/Y sky130_fd_sc_hd__bufinv_16
Xclkload56 clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 clkload56/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload45 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 clkload45/Y sky130_fd_sc_hd__inv_6
Xclkload78 clknet_leaf_81_clk vssd1 vssd1 vccd1 vccd1 clkload78/Y sky130_fd_sc_hd__inv_8
XANTENNA_clkbuf_leaf_53_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload89 clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 clkload89/Y sky130_fd_sc_hd__clkinv_4
X_07940_ top.hTree.tree_reg\[0\] top.findLeastValue.sum\[0\] net250 vssd1 vssd1 vccd1
+ vccd1 _04458_ sky130_fd_sc_hd__mux2_1
XANTENNA__08906__C1 _05072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08382__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07871_ net483 _04401_ vssd1 vssd1 vccd1 vccd1 _04403_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_68_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09610_ net851 net691 vssd1 vssd1 vccd1 vccd1 _00224_ sky130_fd_sc_hd__and2_1
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06822_ top.findLeastValue.val1\[8\] net130 net114 top.compVal\[8\] vssd1 vssd1 vccd1
+ vccd1 _02016_ sky130_fd_sc_hd__o22a_1
XFILLER_110_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_09541_ net746 net586 vssd1 vssd1 vccd1 vccd1 _00155_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_111_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06753_ _02413_ top.findLeastValue.val2\[35\] _03532_ _03540_ vssd1 vssd1 vccd1 vccd1
+ _03541_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_104_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05704_ net9 net415 net308 top.WB.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1 _02354_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10021__A net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06684_ _02440_ top.findLeastValue.val2\[9\] top.findLeastValue.val2\[8\] _02441_
+ vssd1 vssd1 vccd1 vccd1 _03472_ sky130_fd_sc_hd__o22a_1
X_09472_ net747 net587 vssd1 vssd1 vccd1 vccd1 _00086_ sky130_fd_sc_hd__and2_1
X_08423_ top.cb_syn.char_path_n\[49\] top.cb_syn.char_path_n\[50\] top.cb_syn.char_path_n\[51\]
+ top.cb_syn.char_path_n\[52\] net514 net510 vssd1 vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__mux4_1
X_05635_ net1129 net138 _02717_ net174 vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__a22o_1
X_08354_ top.cb_syn.char_path_n\[85\] net392 net331 top.cb_syn.char_path_n\[86\] net438
+ vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__a221o_1
X_05566_ net457 top.hTree.node_reg\[51\] net361 net420 top.hTree.node_reg\[19\] vssd1
+ vssd1 vccd1 vccd1 _02660_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout247_A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09021__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07305_ _03792_ _03936_ vssd1 vssd1 vccd1 vccd1 _03937_ sky130_fd_sc_hd__or2_1
XANTENNA__06448__B1 top.controller.state_reg\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_08285_ top.cb_syn.char_path_n\[27\] net385 net344 top.cb_syn.char_path_n\[25\] net189
+ vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__a221o_1
X_05497_ top.cb_syn.char_path\[94\] net554 net545 top.cb_syn.char_path\[62\] vssd1
+ vssd1 vccd1 vccd1 _02602_ sky130_fd_sc_hd__a22o_1
Xclkload6 clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clkload6/X sky130_fd_sc_hd__clkbuf_8
X_07236_ net271 _03884_ _03885_ net276 net1580 vssd1 vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout202_X net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05671__B2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07167_ top.findLeastValue.val1\[35\] top.findLeastValue.val2\[35\] vssd1 vssd1 vccd1
+ vccd1 _03825_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_115_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06118_ _02578_ _02964_ _02987_ _02989_ vssd1 vssd1 vccd1 vccd1 _02990_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout783_A net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07098_ _03748_ _03755_ vssd1 vssd1 vccd1 vccd1 _03756_ sky130_fd_sc_hd__nand2b_1
XFILLER_105_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout210 net211 vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__clkbuf_4
Xfanout232 net235 vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__clkbuf_4
X_06049_ net1042 net144 vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__and2_1
Xfanout221 net224 vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__clkbuf_4
XFILLER_101_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout265 net266 vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__clkbuf_2
Xfanout243 _05261_ vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__clkbuf_2
Xfanout254 net255 vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__clkbuf_4
Xfanout298 _03998_ vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__clkbuf_2
Xfanout287 _03325_ vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__buf_2
X_09808_ net787 net627 vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__and2_1
Xfanout276 net277 vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__buf_2
X_09739_ net777 net617 vssd1 vssd1 vccd1 vccd1 _00353_ sky130_fd_sc_hd__and2_1
XANTENNA__08125__B1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11701_ clknet_leaf_116_clk _02234_ _01056_ vssd1 vssd1 vccd1 vccd1 top.path\[32\]
+ sky130_fd_sc_hd__dfrtp_1
X_11632_ clknet_leaf_55_clk top.dut.bit_buf_next\[4\] _00987_ vssd1 vssd1 vccd1 vccd1
+ top.dut.bit_buf\[4\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11563_ clknet_leaf_37_clk _02111_ _00918_ vssd1 vssd1 vccd1 vccd1 top.header_synthesis.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__07651__A2 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11494_ clknet_leaf_86_clk _02042_ _00849_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[34\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__08770__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10514_ net816 net656 vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__and2_1
X_10445_ net751 net591 vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__and2_1
XANTENNA__07939__A0 top.findLeastValue.sum\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10376_ net855 net695 vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__and2_1
XFILLER_97_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_15_0_clk_X clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05717__A2 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05420_ top.cb_syn.curr_state\[2\] vssd1 vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__inv_2
XFILLER_81_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05351_ top.findLeastValue.least1\[8\] vssd1 vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__inv_2
X_08070_ _04534_ _04556_ vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__or2_1
Xclkload112 clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 clkload112/Y sky130_fd_sc_hd__inv_4
Xclkload101 clknet_leaf_76_clk vssd1 vssd1 vccd1 vccd1 clkload101/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__06850__B1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05653__B2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07021_ top.findLeastValue.val1\[26\] top.findLeastValue.val2\[26\] vssd1 vssd1 vccd1
+ vccd1 _03679_ sky130_fd_sc_hd__nand2_1
X_08972_ top.WB.CPU_DAT_O\[20\] net1357 net321 vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__mux2_1
Xhold18 top.sram_interface.init_counter\[15\] vssd1 vssd1 vccd1 vccd1 net971 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09805__A net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold29 top.hTree.node_reg\[32\] vssd1 vssd1 vccd1 vccd1 net982 sky130_fd_sc_hd__dlygate4sd3_1
X_07923_ net440 net1452 net251 top.findLeastValue.sum\[4\] _04444_ vssd1 vssd1 vccd1
+ vccd1 _01809_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_110_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout197_A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07854_ top.findLeastValue.sum\[17\] top.hTree.tree_reg\[17\] net278 vssd1 vssd1
+ vccd1 vccd1 _04389_ sky130_fd_sc_hd__mux2_1
XFILLER_96_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05708__A2 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06905__A1 top.findLeastValue.val2\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06805_ net496 net129 net113 top.compVal\[25\] vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout364_A net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07785_ top.findLeastValue.sum\[31\] _04333_ net397 vssd1 vssd1 vccd1 vccd1 _04334_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__11843__Q top.WB.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06736_ _03508_ _03523_ _03507_ vssd1 vssd1 vccd1 vccd1 _03524_ sky130_fd_sc_hd__o21a_1
X_09524_ net741 net581 vssd1 vssd1 vccd1 vccd1 _00138_ sky130_fd_sc_hd__and2_1
X_09455_ net869 net709 vssd1 vssd1 vccd1 vccd1 _00069_ sky130_fd_sc_hd__and2_1
XFILLER_52_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06667_ _03447_ _03454_ _03446_ vssd1 vssd1 vccd1 vccd1 _03455_ sky130_fd_sc_hd__a21o_1
X_08406_ top.cb_syn.char_path_n\[26\] net331 _04764_ net511 _02504_ vssd1 vssd1 vccd1
+ vccd1 _04765_ sky130_fd_sc_hd__a221o_1
XFILLER_12_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_05618_ top.cb_syn.char_path\[74\] net551 net542 top.cb_syn.char_path\[42\] vssd1
+ vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__a22o_1
X_09386_ net406 _04261_ vssd1 vssd1 vccd1 vccd1 _05268_ sky130_fd_sc_hd__nand2_1
XFILLER_61_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06598_ _03329_ _03331_ _03383_ _03386_ vssd1 vssd1 vccd1 vccd1 _03387_ sky130_fd_sc_hd__nor4_1
X_08337_ top.cb_syn.char_path_n\[87\] top.cb_syn.char_path_n\[88\] net516 vssd1 vssd1
+ vccd1 vccd1 _04696_ sky130_fd_sc_hd__mux2_1
X_05549_ top.histogram.sram_out\[22\] net365 _02644_ _02645_ vssd1 vssd1 vccd1 vccd1
+ _02646_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout417_X net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07633__A2 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08268_ top.cb_syn.char_path_n\[35\] net201 _04661_ vssd1 vssd1 vccd1 vccd1 _01681_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__06841__A0 top.findLeastValue.least1\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07219_ _03845_ _03872_ vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__or2_1
XFILLER_105_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08199_ top.cb_syn.char_path_n\[70\] net380 net339 top.cb_syn.char_path_n\[68\] net184
+ vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__a221o_1
X_10230_ net829 net669 vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout786_X net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07492__S1 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10161_ net816 net656 vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__and2_1
X_10092_ net834 net674 vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__and2_1
XANTENNA__07934__S net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10994_ clknet_leaf_26_clk _01542_ _00349_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05580__B1 _02671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07857__C1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08744__S1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07321__A1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11615_ clknet_leaf_62_clk _02163_ _00970_ vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__dfrtp_1
XFILLER_51_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_11546_ clknet_leaf_0_clk _02094_ _00901_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06832__B1 _03553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05635__B2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_11477_ clknet_leaf_99_clk _02025_ _00832_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[17\]
+ sky130_fd_sc_hd__dfstp_1
X_10428_ net874 net714 vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__and2_1
X_10359_ net874 net714 vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__and2_1
XANTENNA__07844__S net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_05_890 vssd1 vssd1 vccd1 vccd1 team_05_890/HI gpio_out[5] sky130_fd_sc_hd__conb_1
XFILLER_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06899__B1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07570_ net1474 _04159_ _04144_ vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__mux2_1
XANTENNA__05571__B1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06521_ _03273_ _03314_ vssd1 vssd1 vccd1 vccd1 _02077_ sky130_fd_sc_hd__nor2_1
X_09240_ top.header_synthesis.header\[1\] top.cb_syn.char_index\[1\] net518 vssd1
+ vssd1 vccd1 vccd1 _05205_ sky130_fd_sc_hd__mux2_1
XFILLER_80_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06452_ _03271_ _03274_ vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__and2_1
X_05403_ top.cb_syn.zeroes\[5\] vssd1 vssd1 vccd1 vccd1 _02511_ sky130_fd_sc_hd__inv_2
XANTENNA__05874__A1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09171_ net366 _05101_ _05108_ net1558 vssd1 vssd1 vccd1 vccd1 _00036_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_60_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06383_ net299 _03182_ _03225_ _03226_ vssd1 vssd1 vccd1 vccd1 _02127_ sky130_fd_sc_hd__o31ai_1
XANTENNA__08273__C1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05334_ top.compVal\[7\] vssd1 vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__inv_2
X_08122_ top.cb_syn.char_path_n\[108\] net195 _04588_ vssd1 vssd1 vccd1 vccd1 _01754_
+ sky130_fd_sc_hd__o21a_1
X_08053_ net535 _04538_ vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__nor2_1
X_07004_ top.findLeastValue.val1\[38\] top.findLeastValue.val2\[38\] vssd1 vssd1 vccd1
+ vccd1 _03662_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout112_A net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11838__Q top.WB.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08955_ top.WB.CPU_DAT_O\[18\] top.cb_syn.h_element\[50\] net370 vssd1 vssd1 vccd1
+ vccd1 _01355_ sky130_fd_sc_hd__mux2_1
XANTENNA__07754__S net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05782__B net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout579_A net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07906_ net482 _04429_ vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__or2_1
X_08886_ top.sram_interface.TRN_counter\[0\] _05053_ _05057_ vssd1 vssd1 vccd1 vccd1
+ _01459_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_71_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08423__S0 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07837_ net428 _04374_ _04375_ net262 vssd1 vssd1 vccd1 vccd1 _04376_ sky130_fd_sc_hd__o211a_1
XFILLER_56_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_fanout367_X net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05562__B1 _02656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07768_ net443 net1427 net254 top.findLeastValue.sum\[35\] _04320_ vssd1 vssd1 vccd1
+ vccd1 _01840_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_27_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09507_ net740 net580 vssd1 vssd1 vccd1 vccd1 _00121_ sky130_fd_sc_hd__and2_1
X_06719_ _02420_ top.findLeastValue.val2\[30\] top.findLeastValue.val2\[29\] _02421_
+ vssd1 vssd1 vccd1 vccd1 _03507_ sky130_fd_sc_hd__o22a_1
X_07699_ net397 _04264_ vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_55_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09438_ net965 vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__clkbuf_1
X_09369_ net985 net238 net216 _04310_ vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__a22o_1
XANTENNA__09056__A1 top.WB.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05865__B2 top.WB.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07929__S net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11400_ clknet_leaf_95_clk _01948_ _00755_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[6\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_40_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11331_ clknet_leaf_69_clk _01879_ _00686_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.startup
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__06814__B1 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05617__B2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05957__B net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11262_ clknet_leaf_105_clk _01810_ _00617_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11193_ clknet_leaf_42_clk _01741_ _00548_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[95\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10213_ net825 net665 vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__and2_1
XANTENNA_input42_A gpio_in[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06042__A1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10144_ net826 net666 vssd1 vssd1 vccd1 vccd1 _00758_ sky130_fd_sc_hd__and2_1
XFILLER_48_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10075_ net852 net692 vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_89_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05553__B1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10977_ clknet_leaf_9_clk _01525_ _00332_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05856__B2 top.WB.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09047__A1 top.WB.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__07839__S net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__05500__X _02605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06805__B1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08270__A2 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold307 net82 vssd1 vssd1 vccd1 vccd1 net1260 sky130_fd_sc_hd__dlygate4sd3_1
X_11529_ clknet_leaf_5_clk _02077_ _00884_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold318 top.cb_syn.char_path\[62\] vssd1 vssd1 vccd1 vccd1 net1271 sky130_fd_sc_hd__dlygate4sd3_1
Xhold329 top.path\[93\] vssd1 vssd1 vccd1 vccd1 net1282 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout809 net811 vssd1 vssd1 vccd1 vccd1 net809 sky130_fd_sc_hd__buf_1
XANTENNA__06033__A1 top.WB.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08740_ top.header_synthesis.write_num_lefts _02542_ net296 _04919_ _04923_ vssd1
+ vssd1 vccd1 vccd1 _04924_ sky130_fd_sc_hd__o311a_1
X_05952_ top.WB.CPU_DAT_O\[3\] net1291 net307 vssd1 vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__mux2_1
X_05883_ _02498_ top.cb_syn.wait_cycle vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__nor2_1
X_08671_ _04546_ _04800_ _04803_ net246 net1529 vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__a32o_1
XFILLER_78_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07622_ net262 _04201_ _04202_ net1315 net448 vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__a32o_1
XANTENNA__10013__B net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05544__B1 _02641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07553_ _04128_ _04129_ _04143_ vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__o21a_2
X_07484_ top.cb_syn.char_path_n\[20\] top.cb_syn.char_path_n\[19\] top.cb_syn.char_path_n\[18\]
+ top.cb_syn.char_path_n\[17\] net400 net352 vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_52_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06504_ net1601 _03281_ vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__xor2_1
X_09223_ top.cb_syn.num_lefts\[5\] top.cb_syn.num_lefts\[4\] top.cb_syn.num_lefts\[3\]
+ top.cb_syn.num_lefts\[2\] vssd1 vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__or4_1
X_06435_ top.header_synthesis.enable top.header_synthesis.char_added top.header_synthesis.write_num_lefts
+ vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__a21o_1
XANTENNA__09038__A1 top.WB.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05847__B2 top.WB.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09154_ net549 net470 _02547_ _02767_ vssd1 vssd1 vccd1 vccd1 _05160_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_32_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout327_A net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07749__S net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08105_ top.cb_syn.char_path_n\[117\] net383 net342 top.cb_syn.char_path_n\[115\]
+ net187 vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__a221o_1
X_06366_ _03187_ _03215_ net301 vssd1 vssd1 vccd1 vccd1 _03216_ sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_4_3_0_clk_X clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06297_ net467 _03156_ _03158_ _03161_ vssd1 vssd1 vccd1 vccd1 _03162_ sky130_fd_sc_hd__a31o_1
X_09085_ _05104_ _05105_ vssd1 vssd1 vccd1 vccd1 _05106_ sky130_fd_sc_hd__nor2_1
X_05317_ top.compVal\[25\] vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout115_X net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08036_ _04530_ vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout696_A net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06024__A1 top.WB.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09987_ net864 net704 vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout863_A net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07772__A1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08938_ top.WB.CPU_DAT_O\[16\] net1303 net371 vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08869_ net437 _05047_ vssd1 vssd1 vccd1 vccd1 _05048_ sky130_fd_sc_hd__nand2_1
X_10900_ clknet_leaf_39_clk top.header_synthesis.next_header\[5\] _00255_ vssd1 vssd1
+ vccd1 vccd1 top.header_synthesis.header\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_84_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05535__B1 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11880_ clknet_leaf_23_clk _02396_ _01235_ vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_84_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10831_ clknet_leaf_46_clk _01417_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_10762_ clknet_leaf_47_clk _01361_ _00181_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08047__C net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09029__A1 top.WB.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05838__B2 top.WB.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10693_ clknet_leaf_112_clk _01292_ _00112_ vssd1 vssd1 vccd1 vccd1 top.path\[69\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11314_ clknet_leaf_77_clk _01862_ _00669_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_10_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11245_ clknet_leaf_68_clk _01793_ _00600_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.alternator_timer\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__06015__A1 top.WB.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11176_ clknet_leaf_8_clk _01724_ _00531_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[78\]
+ sky130_fd_sc_hd__dfrtp_1
X_10127_ net839 net679 vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__and2_1
X_10058_ net859 net699 vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__and2_1
XANTENNA__05526__B1 _02626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06220_ net500 _03012_ vssd1 vssd1 vccd1 vccd1 _03088_ sky130_fd_sc_hd__nor2_1
X_06151_ top.hist_addr\[5\] top.hist_addr\[4\] _03021_ vssd1 vssd1 vccd1 vccd1 _03022_
+ sky130_fd_sc_hd__and3_1
X_06082_ _02851_ _02954_ _02582_ vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__a21oi_1
Xhold104 top.header_synthesis.header\[0\] vssd1 vssd1 vccd1 vccd1 net1057 sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 net95 vssd1 vssd1 vccd1 vccd1 net1079 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold115 top.path\[13\] vssd1 vssd1 vccd1 vccd1 net1068 sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 top.cb_syn.char_path\[68\] vssd1 vssd1 vccd1 vccd1 net1090 sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 top.path\[126\] vssd1 vssd1 vccd1 vccd1 net1101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold159 top.path\[111\] vssd1 vssd1 vccd1 vccd1 net1112 sky130_fd_sc_hd__dlygate4sd3_1
X_09910_ net758 net598 vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__and2_1
XANTENNA__06006__A1 top.WB.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout606 net607 vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__clkbuf_2
Xfanout639 net640 vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__clkbuf_2
Xfanout617 net619 vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkload14_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08951__A0 top.WB.CPU_DAT_O\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout628 net631 vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__clkbuf_2
X_09841_ net787 net627 vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__and2_1
XANTENNA__08400__C1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09772_ net790 net630 vssd1 vssd1 vccd1 vccd1 _00386_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_13_Left_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06984_ top.findLeastValue.val1\[10\] top.findLeastValue.val1\[9\] top.findLeastValue.val1\[8\]
+ top.findLeastValue.val1\[7\] vssd1 vssd1 vccd1 vccd1 _03642_ sky130_fd_sc_hd__and4_1
XANTENNA__10024__A net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08723_ top.cb_syn.i\[2\] _04898_ _04905_ _04910_ vssd1 vssd1 vccd1 vccd1 _01475_
+ sky130_fd_sc_hd__a22o_1
X_05935_ top.WB.CPU_DAT_O\[20\] net1416 net304 vssd1 vssd1 vccd1 vccd1 _02254_ sky130_fd_sc_hd__mux2_1
XANTENNA__08703__A0 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout277_A _03658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05517__B1 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08654_ _04801_ _04857_ _04563_ vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07604__Y _04188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05866_ top.compVal\[1\] net170 net156 top.WB.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1
+ _02276_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06190__B1 top.cb_syn.char_index\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08585_ _04811_ top.cb_syn.char_index\[4\] _04807_ vssd1 vssd1 vccd1 vccd1 _01514_
+ sky130_fd_sc_hd__mux2_1
X_05797_ _02815_ _02816_ vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__nand2_1
X_07605_ net445 _04187_ vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout444_A net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11851__Q top.WB.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09024__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07536_ _04126_ _04125_ vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__and2b_1
XFILLER_41_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_22_Left_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07467_ _04056_ _04057_ _04055_ vssd1 vssd1 vccd1 vccd1 _04058_ sky130_fd_sc_hd__a21o_2
X_09206_ _02530_ _02873_ vssd1 vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout611_A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06418_ top.header_synthesis.count\[5\] _03245_ _03248_ vssd1 vssd1 vccd1 vccd1 _03249_
+ sky130_fd_sc_hd__and3_1
X_07398_ net297 vssd1 vssd1 vccd1 vccd1 top.dut.out_valid_next sky130_fd_sc_hd__inv_2
X_09137_ net465 _05132_ top.sram_interface.word_cnt\[9\] vssd1 vssd1 vccd1 vccd1 _05148_
+ sky130_fd_sc_hd__o21a_1
X_06349_ net1468 _03205_ net302 vssd1 vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__mux2_1
X_09068_ top.CB_write_complete top.cb_syn.end_cond net529 net474 top.cb_syn.curr_state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05092_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_118_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08019_ _04516_ _04520_ top.cb_syn.count\[6\] vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__a21o_1
XANTENNA__06796__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold671 top.cb_syn.curr_index\[7\] vssd1 vssd1 vccd1 vccd1 net1624 sky130_fd_sc_hd__dlygate4sd3_1
Xhold660 top.findLeastValue.sum\[33\] vssd1 vssd1 vccd1 vccd1 net1613 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_31_Left_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11030_ clknet_leaf_27_clk _01578_ _00385_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[60\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold682 top.sram_interface.write_counter_FLV\[1\] vssd1 vssd1 vccd1 vccd1 net1635
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold693 top.hist_data_o\[23\] vssd1 vssd1 vccd1 vccd1 net1646 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout866_X net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08942__A0 top.WB.CPU_DAT_O\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11863_ clknet_leaf_115_clk _02379_ _01218_ vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__dfrtp_1
X_10814_ clknet_leaf_106_clk _01400_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_40_Left_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11794_ clknet_leaf_58_clk _00012_ _01149_ vssd1 vssd1 vccd1 vccd1 top.controller.state_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10745_ clknet_leaf_120_clk _01344_ _00164_ vssd1 vssd1 vccd1 vccd1 top.path\[121\]
+ sky130_fd_sc_hd__dfrtp_1
X_10676_ clknet_leaf_2_clk _01275_ _00095_ vssd1 vssd1 vccd1 vccd1 top.path\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10109__A net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06787__A2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11228_ clknet_leaf_35_clk _01776_ _00583_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.end_cnt\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_4_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11159_ clknet_leaf_18_clk _01707_ _00514_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[61\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08933__A0 top.WB.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06539__A2 top.findLeastValue.val1\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06041__B net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05720_ net2 net416 net309 top.WB.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 _02338_
+ sky130_fd_sc_hd__o22a_1
X_05651_ top.hTree.node_reg\[37\] net310 _02730_ net480 vssd1 vssd1 vccd1 vccd1 _02731_
+ sky130_fd_sc_hd__a22o_1
X_08370_ top.cb_syn.char_path_n\[117\] net392 net331 top.cb_syn.char_path_n\[118\]
+ net438 vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_34_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05582_ top.cb_syn.char_path\[16\] net557 net312 top.cb_syn.char_path\[112\] vssd1
+ vssd1 vccd1 vccd1 _02673_ sky130_fd_sc_hd__a22o_1
X_07321_ net269 _03947_ _03948_ net274 net1697 vssd1 vssd1 vccd1 vccd1 _01911_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_102_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07252_ _03887_ _03896_ vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__nor2_1
X_06203_ top.hist_addr\[4\] _03021_ top.hist_addr\[5\] vssd1 vssd1 vccd1 vccd1 _03072_
+ sky130_fd_sc_hd__a21oi_1
X_07183_ top.findLeastValue.val1\[40\] top.findLeastValue.val2\[40\] vssd1 vssd1 vccd1
+ vccd1 _03841_ sky130_fd_sc_hd__nand2_1
X_06134_ _02481_ net368 _02997_ _02998_ vssd1 vssd1 vccd1 vccd1 _03006_ sky130_fd_sc_hd__a22o_1
XANTENNA__10019__A net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08847__S0 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06778__A2 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06065_ net1026 net141 _02941_ vssd1 vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__a21o_1
Xfanout414 _02766_ vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__buf_2
XANTENNA__05774__C top.findLeastValue.least1\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11846__Q top.WB.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09019__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_86_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_fanout394_A net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08924__A0 top.WB.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout447 net448 vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__clkbuf_2
X_09824_ net738 net578 vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__and2_1
Xfanout425 net427 vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__buf_2
Xfanout436 _02523_ vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__clkbuf_4
Xfanout469 top.controller.state_reg\[2\] vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__buf_2
XANTENNA__05738__B1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout458 net462 vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__buf_2
X_06967_ top.findLeastValue.val2\[0\] net149 net122 _03625_ vssd1 vssd1 vccd1 vccd1
+ _01942_ sky130_fd_sc_hd__o22a_1
X_09755_ net736 net576 vssd1 vssd1 vccd1 vccd1 _00369_ sky130_fd_sc_hd__and2_1
X_09686_ net784 net624 vssd1 vssd1 vccd1 vccd1 _00300_ sky130_fd_sc_hd__and2_1
X_05918_ _02453_ _02888_ vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__nand2_1
X_08706_ _04555_ _04897_ vssd1 vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__or2_2
XANTENNA_fanout659_A net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06898_ top.compVal\[34\] top.findLeastValue.val1\[34\] net165 vssd1 vssd1 vccd1
+ vccd1 _03591_ sky130_fd_sc_hd__mux2_1
X_08637_ top.cb_syn.cb_length\[3\] _04847_ vssd1 vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_68_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05849_ top.compVal\[18\] net168 net154 top.WB.CPU_DAT_O\[18\] vssd1 vssd1 vccd1
+ vccd1 _02293_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_81_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout447_X net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout826_A net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08568_ net1349 top.cb_syn.char_path_n\[8\] net225 vssd1 vssd1 vccd1 vccd1 _01526_
+ sky130_fd_sc_hd__mux2_1
X_07519_ top.cb_syn.char_path_n\[120\] top.cb_syn.char_path_n\[119\] top.cb_syn.char_path_n\[118\]
+ top.cb_syn.char_path_n\[117\] net401 net352 vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_12_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08499_ net1186 top.cb_syn.char_path_n\[77\] net221 vssd1 vssd1 vccd1 vccd1 _01595_
+ sky130_fd_sc_hd__mux2_1
X_10530_ net859 net699 vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__and2_1
X_10461_ net723 net563 vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__and2_1
XFILLER_108_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_108_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07966__A1 _02763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07510__S0 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06841__S _03424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10392_ net756 net596 vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__and2_1
XFILLER_108_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_104_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold490 top.hTree.tree_reg\[10\] vssd1 vssd1 vccd1 vccd1 net1443 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11013_ clknet_leaf_4_clk _01561_ _00368_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07718__A1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07672__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11491__Q top.findLeastValue.val1\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11846_ clknet_leaf_117_clk _02362_ _01201_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[24\]
+ sky130_fd_sc_hd__dfrtp_4
X_11777_ clknet_leaf_55_clk _02310_ _01132_ vssd1 vssd1 vccd1 vccd1 top.histogram.init_edge
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_4_11_0_clk_X clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10728_ clknet_leaf_118_clk _01327_ _00147_ vssd1 vssd1 vccd1 vccd1 top.path\[104\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload13 clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clkload13/Y sky130_fd_sc_hd__clkinvlp_4
X_10659_ clknet_leaf_114_clk _01258_ _00078_ vssd1 vssd1 vccd1 vccd1 top.path\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload35 clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 clkload35/X sky130_fd_sc_hd__clkbuf_4
Xclkload24 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 clkload24/X sky130_fd_sc_hd__clkbuf_8
Xclkload68 clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 clkload68/Y sky130_fd_sc_hd__bufinv_16
Xclkload46 clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 clkload46/Y sky130_fd_sc_hd__clkinv_4
Xclkload57 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 clkload57/Y sky130_fd_sc_hd__inv_4
XANTENNA__09628__A net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload79 clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 clkload79/Y sky130_fd_sc_hd__inv_6
XANTENNA__07709__B2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_110_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08382__A1 top.cb_syn.char_path_n\[101\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07870_ top.hTree.tree_reg\[14\] top.findLeastValue.sum\[14\] net247 vssd1 vssd1
+ vccd1 vccd1 _04402_ sky130_fd_sc_hd__mux2_1
XFILLER_110_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06821_ top.findLeastValue.val1\[9\] net130 net114 net1713 vssd1 vssd1 vccd1 vccd1
+ _02017_ sky130_fd_sc_hd__o22a_1
X_09540_ net732 net572 vssd1 vssd1 vccd1 vccd1 _00154_ sky130_fd_sc_hd__and2_1
X_06752_ _03528_ _03529_ _03530_ vssd1 vssd1 vccd1 vccd1 _03540_ sky130_fd_sc_hd__or3_1
X_05703_ net10 net417 net359 top.WB.CPU_DAT_O\[17\] vssd1 vssd1 vccd1 vccd1 _02355_
+ sky130_fd_sc_hd__a22o_1
X_09471_ net747 net587 vssd1 vssd1 vccd1 vccd1 _00085_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_104_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10021__B net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08422_ top.cb_syn.char_path_n\[45\] top.cb_syn.char_path_n\[46\] top.cb_syn.char_path_n\[47\]
+ top.cb_syn.char_path_n\[48\] net514 net510 vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_47_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06683_ _03468_ _03469_ _03470_ vssd1 vssd1 vccd1 vccd1 _03471_ sky130_fd_sc_hd__a21o_1
XANTENNA__05499__A2 _02603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06926__S net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05634_ top.histogram.sram_out\[8\] net363 net419 top.hTree.node_reg\[8\] _02716_
+ vssd1 vssd1 vccd1 vccd1 _02717_ sky130_fd_sc_hd__a221o_1
XFILLER_36_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout142_A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05565_ _02657_ _02658_ net472 vssd1 vssd1 vccd1 vccd1 _02659_ sky130_fd_sc_hd__o21a_1
X_08353_ top.cb_syn.char_path_n\[69\] net391 net330 top.cb_syn.char_path_n\[70\] net438
+ vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__a221o_1
XANTENNA__08437__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08284_ top.cb_syn.char_path_n\[27\] net206 _04669_ vssd1 vssd1 vccd1 vccd1 _01673_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_63_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07304_ _03787_ _03935_ _03786_ vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__a21bo_1
XFILLER_20_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06448__A1 _03269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05496_ net1133 net139 _02601_ net175 vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__a22o_1
Xclkload7 clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clkload7/Y sky130_fd_sc_hd__clkinvlp_4
X_07235_ _03668_ _03883_ vssd1 vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__nand2_1
XANTENNA__08842__C1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07166_ _03822_ _03823_ vssd1 vssd1 vccd1 vccd1 _03824_ sky130_fd_sc_hd__nor2_1
XANTENNA__05671__A2 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06117_ top.TRN_char_index\[6\] _02973_ _02988_ vssd1 vssd1 vccd1 vccd1 _02989_ sky130_fd_sc_hd__o21a_1
X_07097_ top.findLeastValue.val1\[2\] top.findLeastValue.val2\[2\] vssd1 vssd1 vccd1
+ vccd1 _03755_ sky130_fd_sc_hd__or2_1
X_06048_ net1326 _02592_ net160 vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__a21o_1
XFILLER_105_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout211 _04565_ vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout776_A net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout222 net224 vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout397_X net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout200 net203 vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__buf_2
XFILLER_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout233 net234 vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__clkbuf_4
Xfanout244 net245 vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__buf_2
Xfanout255 net256 vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__buf_2
X_07999_ top.cb_syn.count\[4\] _02512_ _02513_ top.cb_syn.count\[3\] _04501_ vssd1
+ vssd1 vccd1 vccd1 _04502_ sky130_fd_sc_hd__o221a_1
X_09807_ net791 net631 vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__and2_1
Xfanout266 net267 vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08373__B2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout288 _03324_ vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__buf_2
Xfanout277 _03658_ vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__buf_2
Xfanout299 _03172_ vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__clkbuf_4
X_09738_ net777 net617 vssd1 vssd1 vccd1 vccd1 _00352_ sky130_fd_sc_hd__and2_1
XFILLER_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09669_ net780 net620 vssd1 vssd1 vccd1 vccd1 _00283_ sky130_fd_sc_hd__and2_1
X_11700_ clknet_leaf_49_clk _02233_ _01055_ vssd1 vssd1 vccd1 vccd1 top.TRN_sram_complete
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07884__A0 top.findLeastValue.sum\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11631_ clknet_leaf_56_clk top.dut.bit_buf_next\[3\] _00986_ vssd1 vssd1 vccd1 vccd1
+ top.dut.bit_buf\[3\] sky130_fd_sc_hd__dfrtp_1
X_11562_ clknet_leaf_37_clk _02110_ _00917_ vssd1 vssd1 vccd1 vccd1 top.header_synthesis.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10513_ net821 net661 vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__and2_1
X_11493_ clknet_leaf_86_clk _02041_ _00848_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[33\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10444_ net751 net591 vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__and2_1
X_10375_ net854 net694 vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__and2_1
XFILLER_97_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__08498__S net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11829_ clknet_leaf_115_clk _02345_ _01184_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_05350_ top.cw1\[0\] vssd1 vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__inv_2
XANTENNA__07627__A0 top.findLeastValue.least1\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_112_Right_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload113 clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 clkload113/Y sky130_fd_sc_hd__bufinv_16
Xclkload102 clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 clkload102/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__06850__A1 top.findLeastValue.least2\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05653__A2 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07020_ _03676_ _03677_ vssd1 vssd1 vccd1 vccd1 _03678_ sky130_fd_sc_hd__and2_1
XANTENNA__09077__B net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08971_ top.WB.CPU_DAT_O\[21\] net1385 net321 vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__mux2_1
XFILLER_114_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09805__B net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold19 top.hTree.node_reg\[0\] vssd1 vssd1 vccd1 vccd1 net972 sky130_fd_sc_hd__dlygate4sd3_1
X_07922_ net425 _04442_ _04443_ net258 vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_110_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07606__A net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07853_ net441 net1444 net253 top.findLeastValue.sum\[18\] _04388_ vssd1 vssd1 vccd1
+ vccd1 _01823_ sky130_fd_sc_hd__a221o_1
XFILLER_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06804_ top.findLeastValue.val1\[26\] net129 net113 top.compVal\[26\] vssd1 vssd1
+ vccd1 vccd1 _02034_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07784_ top.findLeastValue.sum\[31\] top.hTree.tree_reg\[31\] net280 vssd1 vssd1
+ vccd1 vccd1 _04333_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06735_ _02422_ top.findLeastValue.val2\[28\] _03511_ _03522_ vssd1 vssd1 vccd1 vccd1
+ _03523_ sky130_fd_sc_hd__o22a_1
X_09523_ net733 net573 vssd1 vssd1 vccd1 vccd1 _00137_ sky130_fd_sc_hd__and2_1
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_09454_ net869 net709 vssd1 vssd1 vccd1 vccd1 _00068_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout357_A _02926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06666_ _03449_ _03450_ _03453_ _03448_ vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__a22o_1
XFILLER_36_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08405_ top.cb_syn.char_path_n\[27\] top.cb_syn.char_path_n\[28\] net515 vssd1 vssd1
+ vccd1 vccd1 _04764_ sky130_fd_sc_hd__mux2_1
X_09385_ net1005 net240 _05266_ _05267_ vssd1 vssd1 vccd1 vccd1 _01442_ sky130_fd_sc_hd__a22o_1
X_05617_ net1384 net138 _02702_ net174 vssd1 vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__a22o_1
XFILLER_12_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_fanout145_X net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08336_ net517 net210 _04695_ vssd1 vssd1 vccd1 vccd1 _01647_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout524_A net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06597_ _03327_ _03330_ _03385_ _03328_ vssd1 vssd1 vccd1 vccd1 _03386_ sky130_fd_sc_hd__or4b_1
X_05548_ net456 top.hTree.node_reg\[54\] net361 net420 top.hTree.node_reg\[22\] vssd1
+ vssd1 vccd1 vccd1 _02645_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_22_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05479_ _02552_ _02558_ _02571_ _02586_ vssd1 vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__nor4_1
XANTENNA__08291__B1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout312_X net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08267_ top.cb_syn.char_path_n\[36\] net380 net340 top.cb_syn.char_path_n\[34\] net184
+ vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__a221o_1
XFILLER_117_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__05796__A net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06841__A1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08198_ top.cb_syn.char_path_n\[70\] net201 _04626_ vssd1 vssd1 vccd1 vccd1 _01716_
+ sky130_fd_sc_hd__o21a_1
X_07218_ _03839_ _03842_ _03841_ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_76_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07149_ _03783_ _03784_ _03793_ _03799_ vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__or4_1
XFILLER_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Left_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10160_ net820 net660 vssd1 vssd1 vccd1 vccd1 _00774_ sky130_fd_sc_hd__and2_1
X_10091_ net827 net667 vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__and2_1
XFILLER_47_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10993_ clknet_leaf_24_clk _01541_ _00348_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05580__B2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_52_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07251__A _03817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11614_ clknet_leaf_63_clk _02162_ _00969_ vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__dfrtp_1
XFILLER_11_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_clkbuf_leaf_67_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11545_ clknet_leaf_0_clk _02093_ _00900_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11476_ clknet_leaf_100_clk _02024_ _00831_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[16\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__05635__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10427_ net874 net714 vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_110_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08585__A1 top.cb_syn.char_index\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10358_ net871 net711 vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__and2_1
X_10289_ net724 net564 vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__and2_1
Xteam_05_880 vssd1 vssd1 vccd1 vccd1 team_05_880/HI ADR_O[0] sky130_fd_sc_hd__conb_1
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xteam_05_891 vssd1 vssd1 vccd1 vccd1 team_05_891/HI gpio_out[6] sky130_fd_sc_hd__conb_1
XFILLER_93_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07860__S net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire325_A _05035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_69_Left_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07848__B1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06520_ top.histogram.total\[1\] _03272_ net1608 vssd1 vssd1 vccd1 vccd1 _03314_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06451_ top.histogram.total\[3\] top.histogram.total\[2\] top.histogram.total\[1\]
+ top.histogram.total\[0\] vssd1 vssd1 vccd1 vccd1 _03274_ sky130_fd_sc_hd__and4_1
XFILLER_34_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_05402_ top.cb_syn.zeroes\[6\] vssd1 vssd1 vccd1 vccd1 _02510_ sky130_fd_sc_hd__inv_2
X_09170_ top.histogram.state\[6\] net295 _05164_ net1472 vssd1 vssd1 vccd1 vccd1 _00035_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_60_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06382_ net1048 net299 vssd1 vssd1 vccd1 vccd1 _03226_ sky130_fd_sc_hd__nand2_1
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05333_ top.compVal\[8\] vssd1 vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_122_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_122_clk
+ sky130_fd_sc_hd__clkbuf_8
X_08121_ top.cb_syn.char_path_n\[109\] net373 net333 top.cb_syn.char_path_n\[107\]
+ net178 vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__a221o_1
XANTENNA__09088__A _03172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08052_ net439 _04541_ net246 vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_78_Left_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07003_ top.findLeastValue.val1\[38\] top.findLeastValue.val2\[38\] vssd1 vssd1 vccd1
+ vccd1 _03661_ sky130_fd_sc_hd__nand2_1
XANTENNA__10027__A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06999__X _03657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09816__A net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08954_ top.WB.CPU_DAT_O\[19\] top.cb_syn.h_element\[51\] net369 vssd1 vssd1 vccd1
+ vccd1 _01356_ sky130_fd_sc_hd__mux2_1
X_07905_ top.hTree.tree_reg\[7\] top.findLeastValue.sum\[7\] net247 vssd1 vssd1 vccd1
+ vccd1 _04430_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout474_A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08885_ net1653 _05057_ vssd1 vssd1 vccd1 vccd1 _01460_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_71_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08423__S1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07836_ net485 _04373_ vssd1 vssd1 vccd1 vccd1 _04375_ sky130_fd_sc_hd__or2_1
XFILLER_112_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_84_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout262_X net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07767_ net430 _04318_ _04319_ net266 vssd1 vssd1 vccd1 vccd1 _04320_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_27_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05562__B2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout739_A net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06718_ _02489_ top.compVal\[24\] _02425_ top.findLeastValue.val2\[25\] vssd1 vssd1
+ vccd1 vccd1 _03506_ sky130_fd_sc_hd__o2bb2a_1
X_09506_ net758 net598 vssd1 vssd1 vccd1 vccd1 _00120_ sky130_fd_sc_hd__and2_1
X_07698_ top.findLeastValue.least2\[2\] top.hTree.tree_reg\[48\] net281 vssd1 vssd1
+ vccd1 vccd1 _04264_ sky130_fd_sc_hd__mux2_1
X_09437_ net970 vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__clkbuf_1
X_06649_ top.compVal\[45\] top.compVal\[44\] _03435_ _03437_ vssd1 vssd1 vccd1 vccd1
+ _03438_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout527_X net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09368_ net975 net238 net216 _04314_ vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_113_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_113_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09299_ net433 _05233_ vssd1 vssd1 vccd1 vccd1 _05234_ sky130_fd_sc_hd__or2_1
X_08319_ top.cb_syn.char_path_n\[10\] net378 net337 top.cb_syn.char_path_n\[8\] net182
+ vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__a221o_1
X_11330_ clknet_leaf_52_clk _01878_ _00685_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.curr_index\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05617__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_11261_ clknet_leaf_105_clk _01809_ _00616_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11192_ clknet_leaf_42_clk _01740_ _00547_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[94\]
+ sky130_fd_sc_hd__dfrtp_2
X_10212_ net825 net665 vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__and2_1
X_10143_ net825 net665 vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__and2_1
XFILLER_0_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10074_ net852 net692 vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__and2_1
XANTENNA_input35_A gpio_in[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08077__A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10976_ clknet_leaf_12_clk _01524_ _00331_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06309__B net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_104_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_104_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08350__S0 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold308 net85 vssd1 vssd1 vccd1 vccd1 net1261 sky130_fd_sc_hd__dlygate4sd3_1
X_11528_ clknet_leaf_5_clk _02076_ _00883_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11459_ clknet_leaf_66_clk _02007_ _00814_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.wipe_the_char_1
+ sky130_fd_sc_hd__dfrtp_1
Xhold319 top.histogram.sram_out\[18\] vssd1 vssd1 vccd1 vccd1 net1272 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07855__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05951_ top.WB.CPU_DAT_O\[4\] net1341 net307 vssd1 vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__mux2_1
X_08670_ _02528_ net1568 _04872_ vssd1 vssd1 vccd1 vccd1 _01490_ sky130_fd_sc_hd__mux2_1
X_05882_ net450 net556 net478 vssd1 vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__and3_1
XANTENNA__07590__S _04144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07621_ top.hTree.tree_reg\[63\] net486 net285 vssd1 vssd1 vccd1 vccd1 _04202_ sky130_fd_sc_hd__or3b_1
XFILLER_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05544__B2 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07552_ _02934_ _04141_ _04142_ vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__and3_1
XANTENNA__10310__A net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06503_ _03306_ net1617 vssd1 vssd1 vccd1 vccd1 _02088_ sky130_fd_sc_hd__nor2_1
X_07483_ top.cb_syn.cb_length\[0\] top.cb_syn.i\[0\] vssd1 vssd1 vccd1 vccd1 _04074_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_52_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06434_ top.header_synthesis.count\[3\] _03260_ _03259_ vssd1 vssd1 vccd1 vccd1 _03261_
+ sky130_fd_sc_hd__a21oi_1
X_09222_ _05192_ vssd1 vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__inv_2
XANTENNA__05847__A2 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06934__S net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_86_Left_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09153_ net463 _05113_ _05130_ top.sram_interface.word_cnt\[14\] vssd1 vssd1 vccd1
+ vccd1 _05159_ sky130_fd_sc_hd__o31a_1
X_06365_ top.hist_data_o\[18\] _03186_ vssd1 vssd1 vccd1 vccd1 _03215_ sky130_fd_sc_hd__nor2_1
XANTENNA__09310__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08104_ top.cb_syn.char_path_n\[117\] net204 _04579_ vssd1 vssd1 vccd1 vccd1 _01763_
+ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout222_A net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05316_ top.compVal\[26\] vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__inv_2
X_09084_ top.histogram.eof_n top.histogram.state\[0\] top.histogram.state\[3\] top.histogram.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__or4_1
X_06296_ _02562_ _02937_ _03155_ net469 _03160_ vssd1 vssd1 vccd1 vccd1 _03161_ sky130_fd_sc_hd__a221o_1
XANTENNA__11849__Q top.WB.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08035_ top.cb_syn.wait_cycle net540 net529 _04527_ net431 vssd1 vssd1 vccd1 vccd1
+ _04530_ sky130_fd_sc_hd__a221o_1
XFILLER_89_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout689_A net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09986_ net864 net704 vssd1 vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout856_A net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout477_X net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_95_Left_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08937_ top.WB.CPU_DAT_O\[17\] net1333 net371 vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08868_ net411 _05040_ vssd1 vssd1 vccd1 vccd1 _05047_ sky130_fd_sc_hd__nor2_1
X_07819_ top.findLeastValue.sum\[24\] top.hTree.tree_reg\[24\] net278 vssd1 vssd1
+ vccd1 vccd1 _04361_ sky130_fd_sc_hd__mux2_1
X_08799_ net432 _04980_ _04981_ vssd1 vssd1 vccd1 vccd1 _04982_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_84_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10830_ clknet_leaf_77_clk _01416_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_10761_ clknet_leaf_44_clk _01360_ _00180_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10692_ clknet_leaf_112_clk _01291_ _00111_ vssd1 vssd1 vccd1 vccd1 top.path\[68\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05838__A2 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05601__X _02689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08788__A1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05687__C _02759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06799__B1 net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11313_ clknet_leaf_84_clk _01861_ _00668_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_113_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_11244_ clknet_leaf_75_clk _01792_ _00599_ vssd1 vssd1 vccd1 vccd1 top.hTree.closing
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_95_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09201__A2 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11175_ clknet_leaf_10_clk _01723_ _00530_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[77\]
+ sky130_fd_sc_hd__dfrtp_2
X_10126_ net839 net679 vssd1 vssd1 vccd1 vccd1 _00740_ sky130_fd_sc_hd__and2_1
X_10057_ net849 net689 vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__and2_1
XANTENNA__08399__S0 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09191__A top.controller.fin_reg\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08173__C1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05526__B2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload0_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10959_ clknet_leaf_65_clk net958 _00314_ vssd1 vssd1 vccd1 vccd1 top.controller.fin_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_90_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05511__X _02614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06150_ top.hist_addr\[2\] top.hist_addr\[1\] top.hist_addr\[0\] top.hist_addr\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__a31o_1
X_06081_ top.sram_interface.init_counter\[9\] _02947_ vssd1 vssd1 vccd1 vccd1 _02954_
+ sky130_fd_sc_hd__xnor2_1
Xhold105 top.hTree.node_reg\[40\] vssd1 vssd1 vccd1 vccd1 net1058 sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 top.cb_syn.char_path\[38\] vssd1 vssd1 vccd1 vccd1 net1069 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 top.sram_interface.word_cnt\[4\] vssd1 vssd1 vccd1 vccd1 net1102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 top.path\[86\] vssd1 vssd1 vccd1 vccd1 net1080 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 top.cb_syn.char_path\[41\] vssd1 vssd1 vccd1 vccd1 net1091 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout618 net619 vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__clkbuf_2
X_09840_ net800 net640 vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__and2_1
Xfanout629 net630 vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__clkbuf_2
Xfanout607 net647 vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__clkbuf_2
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09771_ net782 net622 vssd1 vssd1 vccd1 vccd1 _00385_ sky130_fd_sc_hd__and2_1
XANTENNA__08951__A1 top.cb_syn.h_element\[54\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06983_ _03630_ _03635_ _03640_ net424 vssd1 vssd1 vccd1 vccd1 _03641_ sky130_fd_sc_hd__a31o_1
XANTENNA__10024__B net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08722_ top.cb_syn.i\[2\] _04899_ vssd1 vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__xnor2_1
X_05934_ top.WB.CPU_DAT_O\[21\] net1392 net304 vssd1 vssd1 vccd1 vccd1 _02255_ sky130_fd_sc_hd__mux2_1
XANTENNA__05461__A_N net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08653_ top.cb_syn.cb_length\[2\] _04859_ net210 vssd1 vssd1 vccd1 vccd1 _01494_
+ sky130_fd_sc_hd__mux2_1
X_05865_ top.compVal\[2\] net170 net156 top.WB.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1
+ _02277_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout172_A _02782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08584_ top.cb_syn.h_element\[59\] top.cb_syn.h_element\[50\] net532 vssd1 vssd1
+ vccd1 vccd1 _04811_ sky130_fd_sc_hd__mux2_1
X_05796_ net447 _02529_ vssd1 vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__nor2_1
X_07604_ _02454_ _02801_ vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_37_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07535_ top.cb_syn.cb_length\[6\] _02517_ _04064_ vssd1 vssd1 vccd1 vccd1 _04126_
+ sky130_fd_sc_hd__o21ai_1
X_07466_ top.cb_syn.cb_length\[1\] top.cb_syn.i\[1\] vssd1 vssd1 vccd1 vccd1 _04057_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout437_A _02523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06417_ top.header_synthesis.count\[2\] top.header_synthesis.count\[0\] _03247_ vssd1
+ vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__and3_1
X_09205_ top.CB_read_complete top.cb_syn.setup _02527_ top.CB_write_complete vssd1
+ vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__a211oi_1
XFILLER_22_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07397_ top.dut.bits_in_buf\[3\] _03997_ vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout604_A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09136_ net556 _05142_ _05143_ _05147_ vssd1 vssd1 vccd1 vccd1 _00051_ sky130_fd_sc_hd__a211o_1
X_06348_ top.hist_data_o\[25\] _03191_ _03197_ vssd1 vssd1 vccd1 vccd1 _03205_ sky130_fd_sc_hd__o21ba_1
X_09067_ top.hist_addr\[0\] _05090_ _05091_ top.TRN_char_index\[0\] vssd1 vssd1 vccd1
+ vccd1 _01248_ sky130_fd_sc_hd__a22o_1
X_06279_ top.cb_syn.char_index\[0\] net561 net478 vssd1 vssd1 vccd1 vccd1 _03145_
+ sky130_fd_sc_hd__o21ai_1
X_08018_ top.cb_syn.count\[6\] _04516_ _04520_ _04519_ net1412 vssd1 vssd1 vccd1 vccd1
+ _01790_ sky130_fd_sc_hd__a32o_1
Xhold650 top.cb_syn.zero_count\[5\] vssd1 vssd1 vccd1 vccd1 net1603 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold661 top.hist_data_o\[29\] vssd1 vssd1 vccd1 vccd1 net1614 sky130_fd_sc_hd__dlygate4sd3_1
Xhold672 top.hist_data_o\[17\] vssd1 vssd1 vccd1 vccd1 net1625 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold683 top.histogram.total\[8\] vssd1 vssd1 vccd1 vccd1 net1636 sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 top.histogram.total\[9\] vssd1 vssd1 vccd1 vccd1 net1647 sky130_fd_sc_hd__dlygate4sd3_1
X_09969_ net797 net637 vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__and2_1
XANTENNA__08942__A1 top.cb_syn.h_element\[63\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06953__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05756__B2 top.WB.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08155__C1 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06839__S _03424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05508__B2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07902__C1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08170__A2 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11862_ clknet_leaf_115_clk _02378_ _01217_ vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__dfrtp_1
X_10813_ clknet_leaf_105_clk _01399_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_11793_ clknet_leaf_73_clk _00018_ _01148_ vssd1 vssd1 vccd1 vccd1 top.hTree.state\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10744_ clknet_leaf_120_clk _01343_ _00163_ vssd1 vssd1 vccd1 vccd1 top.path\[120\]
+ sky130_fd_sc_hd__dfrtp_1
X_10675_ clknet_leaf_123_clk _01274_ _00094_ vssd1 vssd1 vccd1 vccd1 top.path\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10109__B net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_107_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_11227_ clknet_leaf_42_clk _01775_ _00582_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.end_cnt\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_11158_ clknet_leaf_19_clk _01706_ _00513_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[60\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__05747__A1 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08394__C1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10109_ net822 net662 vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__and2_1
XFILLER_0_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11089_ clknet_leaf_24_clk _01637_ _00444_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[119\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05506__X _02610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05650_ _02728_ _02729_ vssd1 vssd1 vccd1 vccd1 _02730_ sky130_fd_sc_hd__or2_1
X_05581_ top.cb_syn.char_path\[80\] net551 net542 top.cb_syn.char_path\[48\] vssd1
+ vssd1 vccd1 vccd1 _02672_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_34_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09110__A1 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09110__B2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07320_ _03711_ _03946_ vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__nand2_1
X_07251_ _03817_ _03820_ _03829_ vssd1 vssd1 vccd1 vccd1 _03896_ sky130_fd_sc_hd__and3_1
X_06202_ _03069_ _03070_ net470 vssd1 vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__o21ai_1
X_07182_ top.findLeastValue.val1\[40\] top.findLeastValue.val2\[40\] vssd1 vssd1 vccd1
+ vccd1 _03840_ sky130_fd_sc_hd__or2_1
X_06133_ top.cw2\[6\] _03003_ vssd1 vssd1 vccd1 vccd1 _03005_ sky130_fd_sc_hd__and2_1
XANTENNA__09413__A2 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10019__B net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08847__S1 top.translation.index\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06064_ net1051 net142 net137 vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__a21o_1
Xfanout404 _03987_ vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__buf_2
XANTENNA__08385__C1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09823_ net738 net578 vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__and2_1
Xfanout448 _02455_ vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__clkbuf_2
Xfanout426 net427 vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__clkbuf_2
Xfanout437 _02523_ vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__clkbuf_4
Xfanout415 net416 vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__buf_2
XFILLER_98_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout459 net461 vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__buf_2
XANTENNA_fanout387_A net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06966_ top.compVal\[0\] top.findLeastValue.val1\[0\] net164 vssd1 vssd1 vccd1 vccd1
+ _03625_ sky130_fd_sc_hd__mux2_1
X_09754_ net736 net576 vssd1 vssd1 vccd1 vccd1 _00368_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout175_X net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05917_ _02847_ _02883_ _02886_ _02887_ vssd1 vssd1 vccd1 vccd1 _02888_ sky130_fd_sc_hd__or4b_1
X_09685_ net784 net624 vssd1 vssd1 vccd1 vccd1 _00299_ sky130_fd_sc_hd__and2_1
X_08705_ _02933_ _04871_ _04896_ vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout554_A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06897_ top.findLeastValue.val2\[35\] net151 net125 _03590_ vssd1 vssd1 vccd1 vccd1
+ _01977_ sky130_fd_sc_hd__o22a_1
X_08636_ top.cb_syn.cb_length\[2\] _02927_ _04563_ vssd1 vssd1 vccd1 vccd1 _04847_
+ sky130_fd_sc_hd__or3_1
XANTENNA__08152__A2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05848_ top.compVal\[19\] net168 net154 top.WB.CPU_DAT_O\[19\] vssd1 vssd1 vccd1
+ vccd1 _02294_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_93_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_93_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout342_X net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05779_ _02797_ _02798_ vssd1 vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout819_A net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08567_ net1193 top.cb_syn.char_path_n\[9\] net225 vssd1 vssd1 vccd1 vccd1 _01527_
+ sky130_fd_sc_hd__mux2_1
X_07518_ top.cb_syn.char_path_n\[116\] top.cb_syn.char_path_n\[115\] top.cb_syn.char_path_n\[114\]
+ top.cb_syn.char_path_n\[113\] net400 net351 vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__mux4_1
X_08498_ net1210 top.cb_syn.char_path_n\[78\] net224 vssd1 vssd1 vccd1 vccd1 _01596_
+ sky130_fd_sc_hd__mux2_1
X_07449_ top.dut.bits_in_buf_next\[1\] _04035_ _04038_ _04041_ _04000_ vssd1 vssd1
+ vccd1 vccd1 _04042_ sky130_fd_sc_hd__a221o_1
XANTENNA__07663__A1 top.findLeastValue.least1\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout607_X net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10460_ net723 net563 vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__and2_1
X_09119_ top.sram_interface.word_cnt\[13\] net469 net1102 _05135_ vssd1 vssd1 vccd1
+ vccd1 _00047_ sky130_fd_sc_hd__a22o_1
XANTENNA__09404__A2 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10391_ net755 net595 vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__and2_1
XANTENNA__07510__S1 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold480 top.hTree.tree_reg\[8\] vssd1 vssd1 vccd1 vccd1 net1433 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold491 top.hTree.tree_reg\[18\] vssd1 vssd1 vccd1 vccd1 net1444 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08376__C1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11012_ clknet_leaf_11_clk _01560_ _00367_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08391__A2 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_84_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_60_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11845_ clknet_leaf_117_clk _02361_ _01200_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[23\]
+ sky130_fd_sc_hd__dfrtp_4
X_11776_ clknet_leaf_65_clk _02309_ _01131_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.write_counter_FLV\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07701__B _04266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07654__A1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07654__B2 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10727_ clknet_leaf_113_clk _01326_ _00146_ vssd1 vssd1 vccd1 vccd1 top.path\[103\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload14 clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clkload14/X sky130_fd_sc_hd__clkbuf_8
Xclkload25 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 clkload25/Y sky130_fd_sc_hd__bufinv_16
X_10658_ clknet_leaf_114_clk _01257_ _00077_ vssd1 vssd1 vccd1 vccd1 top.path\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload69 clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 clkload69/Y sky130_fd_sc_hd__inv_8
Xclkload47 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 clkload47/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload58 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 clkload58/X sky130_fd_sc_hd__clkbuf_4
X_10589_ net747 net587 vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__and2_1
XANTENNA__09628__B net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload36 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 clkload36/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__07501__S1 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08906__A1 _04187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__08382__A2 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06917__B1 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06820_ top.findLeastValue.val1\[10\] net130 net114 net1718 vssd1 vssd1 vccd1 vccd1
+ _02018_ sky130_fd_sc_hd__o22a_1
XFILLER_110_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06751_ _02411_ top.findLeastValue.val2\[38\] _03537_ _03538_ vssd1 vssd1 vccd1 vccd1
+ _03539_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_75_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08134__A2 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05702_ net11 net417 net359 top.WB.CPU_DAT_O\[18\] vssd1 vssd1 vccd1 vccd1 _02356_
+ sky130_fd_sc_hd__a22o_1
X_06682_ _02441_ top.findLeastValue.val2\[8\] top.findLeastValue.val2\[7\] _02442_
+ vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__a22o_1
X_09470_ net750 net590 vssd1 vssd1 vccd1 vccd1 _00084_ sky130_fd_sc_hd__and2_1
XFILLER_36_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08421_ net510 _04778_ _04779_ vssd1 vssd1 vccd1 vccd1 _04780_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_47_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07893__B2 top.findLeastValue.sum\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05633_ top.hTree.node_reg\[40\] net310 _02715_ net473 vssd1 vssd1 vccd1 vccd1 _02716_
+ sky130_fd_sc_hd__a22o_1
X_05564_ top.cb_syn.char_path\[19\] net557 net312 top.cb_syn.char_path\[115\] vssd1
+ vssd1 vccd1 vccd1 _02658_ sky130_fd_sc_hd__a22o_1
X_08352_ _02506_ top.cb_syn.char_path_n\[72\] _04710_ net509 vssd1 vssd1 vccd1 vccd1
+ _04711_ sky130_fd_sc_hd__o211a_1
X_08283_ top.cb_syn.char_path_n\[28\] net385 net345 top.cb_syn.char_path_n\[26\] net189
+ vssd1 vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__a221o_1
X_05495_ top.histogram.sram_out\[31\] net365 _02598_ _02600_ vssd1 vssd1 vccd1 vccd1
+ _02601_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_63_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07303_ _03811_ _03920_ _03783_ vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__o21ba_1
XANTENNA__06448__A2 _03270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout135_A net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07234_ _03668_ _03883_ vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__or2_1
Xclkload8 clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clkload8/Y sky130_fd_sc_hd__inv_6
XANTENNA__06942__S net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout302_A net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07165_ top.findLeastValue.val1\[34\] top.findLeastValue.val2\[34\] vssd1 vssd1 vccd1
+ vccd1 _03823_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_115_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06116_ top.TRN_char_index\[6\] _02973_ _02565_ vssd1 vssd1 vccd1 vccd1 _02988_ sky130_fd_sc_hd__a21oi_1
X_07096_ top.findLeastValue.val1\[0\] top.findLeastValue.val2\[0\] _03750_ _03749_
+ vssd1 vssd1 vccd1 vccd1 _03754_ sky130_fd_sc_hd__a31o_1
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06047_ net466 top.histogram.eof_n _02534_ net1047 vssd1 vssd1 vccd1 vccd1 _02173_
+ sky130_fd_sc_hd__a31o_1
Xfanout201 net202 vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__buf_2
Xfanout223 net224 vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09554__A net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout234 net235 vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__clkbuf_4
Xfanout245 _05260_ vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__buf_2
XANTENNA_fanout769_A net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout256 _04191_ vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout671_A net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07998_ top.cb_syn.count\[3\] _02513_ _04498_ _04500_ vssd1 vssd1 vccd1 vccd1 _04501_
+ sky130_fd_sc_hd__a22o_1
X_09806_ net789 net629 vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__and2_1
XFILLER_74_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout267 _04189_ vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__clkbuf_2
Xfanout278 _04198_ vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__clkbuf_4
X_09737_ net777 net617 vssd1 vssd1 vccd1 vccd1 _00351_ sky130_fd_sc_hd__and2_1
X_06949_ top.findLeastValue.val2\[9\] net149 net122 _03616_ vssd1 vssd1 vccd1 vccd1
+ _01951_ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_66_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout557_X net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09668_ net780 net620 vssd1 vssd1 vccd1 vccd1 _00282_ sky130_fd_sc_hd__and2_1
X_08619_ net1559 _04836_ _04837_ _04835_ vssd1 vssd1 vccd1 vccd1 _01506_ sky130_fd_sc_hd__a22o_1
X_09599_ net856 net696 vssd1 vssd1 vccd1 vccd1 _00213_ sky130_fd_sc_hd__and2_1
X_11630_ clknet_leaf_55_clk top.dut.bit_buf_next\[2\] _00985_ vssd1 vssd1 vccd1 vccd1
+ top.dut.bit_buf\[2\] sky130_fd_sc_hd__dfrtp_1
X_11561_ clknet_leaf_37_clk _02109_ _00916_ vssd1 vssd1 vccd1 vccd1 top.header_synthesis.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07636__B2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05647__B1 _02727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10512_ net813 net653 vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__and2_1
X_11492_ clknet_leaf_86_clk _02040_ _00847_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[32\]
+ sky130_fd_sc_hd__dfstp_2
X_10443_ net751 net591 vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__and2_1
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10374_ net855 net695 vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__and2_1
XFILLER_108_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_108_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08061__A1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07495__S0 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09010__A0 top.WB.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout790 net791 vssd1 vssd1 vccd1 vccd1 net790 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_57_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_45_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07875__A1 top.findLeastValue.sum\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05886__B1 top.cb_syn.h_element\[54\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11828_ clknet_leaf_114_clk _02344_ _01183_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_81_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_11759_ clknet_leaf_100_clk _02292_ _01114_ vssd1 vssd1 vccd1 vccd1 top.compVal\[17\]
+ sky130_fd_sc_hd__dfrtp_2
Xclkload103 clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 clkload103/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__06850__A2 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload114 clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 clkload114/Y sky130_fd_sc_hd__inv_6
XFILLER_115_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08052__A1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07486__S0 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06063__B1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08970_ top.WB.CPU_DAT_O\[22\] net1430 net321 vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__mux2_1
X_07921_ net482 _04441_ vssd1 vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__or2_1
XANTENNA__09001__A0 top.WB.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07606__B _04188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07852_ net428 _04386_ _04387_ net261 vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__o211a_1
Xinput1 ACK_I vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_1
X_06803_ top.findLeastValue.val1\[27\] net129 net113 net494 vssd1 vssd1 vccd1 vccd1
+ _02035_ sky130_fd_sc_hd__o22a_1
XFILLER_28_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_48_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_clk sky130_fd_sc_hd__clkbuf_8
X_07783_ net443 net1541 net254 net1726 _04332_ vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__a221o_1
X_09522_ net741 net581 vssd1 vssd1 vccd1 vccd1 _00136_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_65_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06734_ _03506_ _03510_ _03513_ _03512_ _03509_ vssd1 vssd1 vccd1 vccd1 _03522_ sky130_fd_sc_hd__o311a_1
X_09453_ net860 net700 vssd1 vssd1 vccd1 vccd1 _00067_ sky130_fd_sc_hd__and2_1
X_06665_ _03452_ vssd1 vssd1 vccd1 vccd1 _03453_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout252_A net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08404_ net511 _04761_ _04762_ vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__a21oi_1
X_09384_ top.hTree.nulls\[48\] net405 net244 vssd1 vssd1 vccd1 vccd1 _05267_ sky130_fd_sc_hd__o21a_1
X_05616_ top.hTree.node_reg\[43\] net310 _02700_ _02701_ vssd1 vssd1 vccd1 vccd1 _02702_
+ sky130_fd_sc_hd__a211o_1
X_08335_ top.cb_syn.char_path_n\[2\] net389 net193 net535 vssd1 vssd1 vccd1 vccd1
+ _04695_ sky130_fd_sc_hd__a211o_1
XFILLER_52_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06596_ _02422_ top.findLeastValue.val1\[28\] net496 _02425_ _03384_ vssd1 vssd1
+ vccd1 vccd1 _03385_ sky130_fd_sc_hd__a221o_1
X_05547_ _02642_ _02643_ net476 vssd1 vssd1 vccd1 vccd1 _02644_ sky130_fd_sc_hd__o21a_1
XANTENNA__05629__B1 _02712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout138_X net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05478_ _02453_ _02581_ _02585_ vssd1 vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__a21oi_1
X_08266_ top.cb_syn.char_path_n\[36\] net201 _04660_ vssd1 vssd1 vccd1 vccd1 _01682_
+ sky130_fd_sc_hd__o21a_1
X_08197_ top.cb_syn.char_path_n\[71\] net380 net339 top.cb_syn.char_path_n\[69\] net184
+ vssd1 vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__a221o_1
X_07217_ net271 _03868_ _03871_ net276 net1585 vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__a32o_1
XFILLER_106_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08043__A1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07148_ _03802_ _03805_ vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_76_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07079_ top.findLeastValue.val1\[7\] top.findLeastValue.val2\[7\] vssd1 vssd1 vccd1
+ vccd1 _03737_ sky130_fd_sc_hd__and2_1
X_10090_ net832 net672 vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__and2_1
XFILLER_59_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_39_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_8
X_10992_ clknet_leaf_24_clk _01540_ _00347_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06847__S _03424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05580__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold729_A top.findLeastValue.sum\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05604__X _02692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09059__B1 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_106_Left_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11613_ clknet_leaf_62_clk _02161_ _00968_ vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__dfrtp_1
XFILLER_42_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11544_ clknet_leaf_0_clk _02092_ _00899_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06832__A2 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_11475_ clknet_leaf_99_clk _02023_ _00830_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[15\]
+ sky130_fd_sc_hd__dfstp_1
X_10426_ net874 net714 vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_115_Left_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10357_ net872 net712 vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__and2_1
XANTENNA__07793__B1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10288_ net727 net567 vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__and2_1
Xteam_05_881 vssd1 vssd1 vccd1 vccd1 team_05_881/HI ADR_O[1] sky130_fd_sc_hd__conb_1
Xteam_05_892 vssd1 vssd1 vccd1 vccd1 team_05_892/HI gpio_out[7] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_49_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06899__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07848__A1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07848__B2 top.findLeastValue.sum\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06450_ top.histogram.total\[2\] top.histogram.total\[1\] _03272_ vssd1 vssd1 vccd1
+ vccd1 _03273_ sky130_fd_sc_hd__and3_1
X_05401_ top.cb_syn.zeroes\[7\] vssd1 vssd1 vccd1 vccd1 _02509_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_60_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06381_ _03178_ _03181_ top.hist_data_o\[12\] vssd1 vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__a21oi_1
XANTENNA__05897__A net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08120_ top.cb_syn.char_path_n\[109\] net196 _04587_ vssd1 vssd1 vccd1 vccd1 _01755_
+ sky130_fd_sc_hd__o21a_1
X_05332_ top.compVal\[9\] vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__inv_2
X_08051_ _04542_ _04544_ vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__or2_1
XANTENNA__10308__A net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07002_ top.findLeastValue.val1\[39\] top.findLeastValue.val2\[39\] vssd1 vssd1 vccd1
+ vccd1 _03660_ sky130_fd_sc_hd__xor2_1
XFILLER_115_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09816__B net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08953_ top.WB.CPU_DAT_O\[20\] top.cb_syn.h_element\[52\] net369 vssd1 vssd1 vccd1
+ vccd1 _01357_ sky130_fd_sc_hd__mux2_1
XFILLER_102_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07904_ top.findLeastValue.sum\[7\] top.hTree.tree_reg\[7\] net283 vssd1 vssd1 vccd1
+ vccd1 _04429_ sky130_fd_sc_hd__mux2_1
XFILLER_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08884_ net294 _05053_ top.sram_interface.TRN_counter\[0\] vssd1 vssd1 vccd1 vccd1
+ _05057_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_71_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout467_A top.controller.state_reg\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07835_ top.findLeastValue.sum\[21\] _04373_ net394 vssd1 vssd1 vccd1 vccd1 _04374_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__08448__A net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05562__A2 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07766_ net490 _04317_ vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_27_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09505_ net758 net598 vssd1 vssd1 vccd1 vccd1 _00119_ sky130_fd_sc_hd__and2_1
X_06717_ _02419_ top.findLeastValue.val2\[31\] top.findLeastValue.val2\[30\] _02420_
+ vssd1 vssd1 vccd1 vccd1 _03505_ sky130_fd_sc_hd__a22o_1
X_09436_ net971 vssd1 vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__clkbuf_1
X_07697_ net265 _04262_ _04263_ net1020 net446 vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout255_X net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06648_ top.compVal\[35\] top.compVal\[34\] top.compVal\[33\] top.compVal\[32\] vssd1
+ vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout422_X net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09367_ net974 net242 net218 _04318_ vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__a22o_1
X_06579_ _02439_ top.findLeastValue.val1\[10\] top.findLeastValue.val1\[9\] _02440_
+ vssd1 vssd1 vccd1 vccd1 _03368_ sky130_fd_sc_hd__a22o_1
X_09298_ top.histogram.total\[6\] top.histogram.total\[7\] top.translation.index\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__mux2_1
X_08318_ top.cb_syn.char_path_n\[10\] net196 _04686_ vssd1 vssd1 vccd1 vccd1 _01656_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__06814__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08249_ top.cb_syn.char_path_n\[45\] net373 net333 top.cb_syn.char_path_n\[43\] net178
+ vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__a221o_1
XFILLER_108_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_fanout791_X net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11260_ clknet_leaf_89_clk _01808_ _00615_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11191_ clknet_leaf_18_clk _01739_ _00546_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[93\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_79_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10211_ net825 net665 vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__and2_1
X_10142_ net825 net665 vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__and2_1
X_10073_ net852 net692 vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_7_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_89_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input28_A DAT_I[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10975_ clknet_leaf_14_clk _01523_ _00330_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_94_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08255__A1 top.cb_syn.char_path_n\[42\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08350__S1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06805__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11527_ clknet_leaf_5_clk _02075_ _00882_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10128__A net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11458_ clknet_leaf_72_clk _02006_ _00813_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least2\[8\]
+ sky130_fd_sc_hd__dfstp_2
Xhold309 top.cb_syn.char_path\[101\] vssd1 vssd1 vccd1 vccd1 net1262 sky130_fd_sc_hd__dlygate4sd3_1
X_10409_ net794 net634 vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__and2_1
X_11389_ clknet_leaf_83_clk _01937_ _00744_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_05950_ top.WB.CPU_DAT_O\[5\] net1434 net306 vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__mux2_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05881_ top.sram_interface.zero_cnt\[0\] _02854_ _02853_ vssd1 vssd1 vccd1 vccd1
+ _02271_ sky130_fd_sc_hd__mux2_1
X_07620_ net486 _04200_ vssd1 vssd1 vccd1 vccd1 _04201_ sky130_fd_sc_hd__nand2_1
XANTENNA__05544__A2 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07551_ _02554_ _02861_ _02858_ vssd1 vssd1 vccd1 vccd1 _04142_ sky130_fd_sc_hd__a21bo_1
XFILLER_19_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__10310__B net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06502_ top.histogram.total\[12\] _03281_ net1616 vssd1 vssd1 vccd1 vccd1 _03307_
+ sky130_fd_sc_hd__a21oi_1
X_07482_ _04056_ _04057_ vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_52_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06433_ top.header_synthesis.count\[2\] top.header_synthesis.count\[1\] top.header_synthesis.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__or3_1
X_09221_ top.header_synthesis.start _03261_ _04917_ vssd1 vssd1 vccd1 vccd1 _05192_
+ sky130_fd_sc_hd__or3b_1
X_09152_ net459 net1652 _02774_ net546 _05158_ vssd1 vssd1 vccd1 vccd1 _00042_ sky130_fd_sc_hd__a221o_1
X_06364_ net1239 _03214_ net302 vssd1 vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08103_ top.cb_syn.char_path_n\[118\] net383 net342 top.cb_syn.char_path_n\[116\]
+ net187 vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__a221o_1
X_05315_ net494 vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__inv_2
X_09083_ top.histogram.state\[2\] top.histogram.state\[5\] top.histogram.state\[7\]
+ top.histogram.state\[6\] vssd1 vssd1 vccd1 vccd1 _05104_ sky130_fd_sc_hd__or4_1
X_06295_ top.cb_syn.curr_index\[1\] _02558_ _03159_ net460 vssd1 vssd1 vccd1 vccd1
+ _03160_ sky130_fd_sc_hd__a22o_1
XANTENNA__05777__D top.findLeastValue.least2\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout215_A net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08034_ net529 _04527_ vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__nand2_1
XANTENNA__06950__S net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07618__Y _04199_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_51_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09985_ net846 net686 vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout584_A net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08936_ top.WB.CPU_DAT_O\[18\] net1211 net371 vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout372_X net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08867_ _05045_ _05046_ top.translation.index\[5\] vssd1 vssd1 vccd1 vccd1 _01467_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout849_A net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_66_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07524__A3 top.cb_syn.char_path_n\[101\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07818_ net441 net1539 net252 top.findLeastValue.sum\[25\] _04360_ vssd1 vssd1 vccd1
+ vccd1 _01830_ sky130_fd_sc_hd__a221o_1
XFILLER_45_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08798_ top.path\[28\] net408 net326 top.path\[29\] net521 vssd1 vssd1 vccd1 vccd1
+ _04981_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_84_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07749_ top.findLeastValue.sum\[38\] top.hTree.tree_reg\[38\] net284 vssd1 vssd1
+ vccd1 vccd1 _04305_ sky130_fd_sc_hd__mux2_1
X_10760_ clknet_leaf_43_clk _01359_ _00179_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[54\]
+ sky130_fd_sc_hd__dfrtp_2
X_09419_ top.hTree.nulls\[60\] net407 net245 vssd1 vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__o21a_1
X_10691_ clknet_leaf_112_clk _01290_ _00110_ vssd1 vssd1 vccd1 vccd1 top.path\[67\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06799__A1 top.findLeastValue.val1\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11312_ clknet_leaf_46_clk _01860_ _00667_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[55\]
+ sky130_fd_sc_hd__dfrtp_1
X_11243_ clknet_leaf_40_clk _01791_ _00598_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.check_right
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_106_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_19_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07748__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06161__A top.cb_syn.char_index\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11174_ clknet_leaf_4_clk _01722_ _00529_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[76\]
+ sky130_fd_sc_hd__dfrtp_2
X_10125_ net839 net679 vssd1 vssd1 vccd1 vccd1 _00739_ sky130_fd_sc_hd__and2_1
X_10056_ net858 net698 vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__and2_1
XANTENNA__08399__S1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09191__B top.controller.fin_reg\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08173__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05526__A2 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07920__A0 top.findLeastValue.sum\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10958_ clknet_leaf_69_clk net955 _00313_ vssd1 vssd1 vccd1 vccd1 top.controller.fin_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10889_ clknet_leaf_111_clk _01466_ _00244_ vssd1 vssd1 vccd1 vccd1 top.translation.index\[4\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__06981__D top.findLeastValue.val2\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_06080_ net1309 net143 _02953_ net159 vssd1 vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__a22o_1
Xhold117 top.cb_syn.char_path\[31\] vssd1 vssd1 vccd1 vccd1 net1070 sky130_fd_sc_hd__dlygate4sd3_1
Xhold106 top.path\[22\] vssd1 vssd1 vccd1 vccd1 net1059 sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 top.cb_syn.char_path\[30\] vssd1 vssd1 vccd1 vccd1 net1092 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold128 top.path\[31\] vssd1 vssd1 vccd1 vccd1 net1081 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout619 net626 vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__buf_1
XFILLER_98_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout608 net609 vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08400__B2 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_107_Right_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09770_ net782 net622 vssd1 vssd1 vccd1 vccd1 _00384_ sky130_fd_sc_hd__and2_1
X_06982_ _03636_ _03637_ _03638_ _03639_ vssd1 vssd1 vccd1 vccd1 _03640_ sky130_fd_sc_hd__and4_1
X_08721_ _04901_ _04905_ _04909_ _04898_ top.cb_syn.i\[3\] vssd1 vssd1 vccd1 vccd1
+ _01476_ sky130_fd_sc_hd__a32o_1
X_05933_ top.WB.CPU_DAT_O\[22\] net1202 net304 vssd1 vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__mux2_1
X_08652_ _04856_ _04858_ vssd1 vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__xnor2_1
XFILLER_66_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07603_ _02454_ _02801_ vssd1 vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__and2_2
X_05864_ top.compVal\[3\] net170 net156 top.WB.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1
+ _02278_ sky130_fd_sc_hd__a22o_1
XANTENNA__05415__A net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08583_ _04810_ top.cb_syn.char_index\[5\] _04807_ vssd1 vssd1 vccd1 vccd1 _01515_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__06010__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05795_ top.hTree.state\[6\] top.hTree.state\[9\] _02806_ vssd1 vssd1 vccd1 vccd1
+ _02815_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout165_A net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07534_ _04123_ _04124_ vssd1 vssd1 vccd1 vccd1 _04125_ sky130_fd_sc_hd__or2_1
XFILLER_81_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07465_ top.cb_syn.cb_length\[0\] top.cb_syn.i\[0\] vssd1 vssd1 vccd1 vccd1 _04056_
+ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_17_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_06416_ top.header_synthesis.count\[4\] top.header_synthesis.count\[3\] top.header_synthesis.count\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03247_ sky130_fd_sc_hd__and3_1
X_09204_ net1515 net257 _05181_ _03324_ vssd1 vssd1 vccd1 vccd1 _00019_ sky130_fd_sc_hd__a22o_1
X_07396_ _02405_ _03995_ vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__nor2_1
X_09135_ _05145_ _05146_ _02877_ vssd1 vssd1 vccd1 vccd1 _05147_ sky130_fd_sc_hd__or3b_1
X_06347_ net1301 _03204_ net302 vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__mux2_1
X_09066_ top.hist_addr\[1\] _05090_ _05091_ top.TRN_char_index\[1\] vssd1 vssd1 vccd1
+ vccd1 _01249_ sky130_fd_sc_hd__a22o_1
X_06278_ top.cb_syn.max_index\[2\] _03025_ _03027_ top.hTree.nullSumIndex\[1\] vssd1
+ vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__a22o_1
XANTENNA__09147__D_N net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout799_A net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08017_ net538 net476 _04507_ vssd1 vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__and3_2
XFILLER_118_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold651 top.hist_data_o\[27\] vssd1 vssd1 vccd1 vccd1 net1604 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold662 top.hist_data_o\[26\] vssd1 vssd1 vccd1 vccd1 net1615 sky130_fd_sc_hd__dlygate4sd3_1
Xhold640 top.findLeastValue.sum\[28\] vssd1 vssd1 vccd1 vccd1 net1593 sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 top.hist_addr\[3\] vssd1 vssd1 vccd1 vccd1 net1637 sky130_fd_sc_hd__dlygate4sd3_1
Xhold673 top.hist_data_o\[25\] vssd1 vssd1 vccd1 vccd1 net1626 sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 top.findLeastValue.sum\[18\] vssd1 vssd1 vccd1 vccd1 net1648 sky130_fd_sc_hd__dlygate4sd3_1
X_09968_ net797 net637 vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__and2_1
XFILLER_103_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08919_ _04180_ _04188_ _05072_ vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__o21ai_1
X_09899_ net790 net630 vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__and2_1
XANTENNA__05508__A2 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_84_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11861_ clknet_leaf_100_clk _02377_ _01216_ vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__dfrtp_1
X_11792_ clknet_leaf_74_clk _00027_ _01147_ vssd1 vssd1 vccd1 vccd1 top.hTree.state\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10812_ clknet_leaf_105_clk _01398_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_10743_ clknet_leaf_2_clk _01342_ _00162_ vssd1 vssd1 vccd1 vccd1 top.path\[119\]
+ sky130_fd_sc_hd__dfrtp_1
X_10674_ clknet_leaf_122_clk _01273_ _00093_ vssd1 vssd1 vccd1 vccd1 top.path\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05692__B2 top.WB.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11226_ clknet_leaf_28_clk _01774_ _00581_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.curr_path\[127\]
+ sky130_fd_sc_hd__dfrtp_1
X_11157_ clknet_leaf_27_clk _01705_ _00512_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[59\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_95_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10108_ net812 net652 vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__and2_1
X_11088_ clknet_leaf_23_clk _01636_ _00443_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[118\]
+ sky130_fd_sc_hd__dfrtp_1
X_10039_ net836 net676 vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_106_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05580_ net1235 net138 _02671_ net174 vssd1 vssd1 vccd1 vccd1 _02387_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_34_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08854__D1 net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07250_ net272 _03894_ _03895_ net277 net1613 vssd1 vssd1 vccd1 vccd1 _01929_ sky130_fd_sc_hd__a32o_1
X_06201_ _03040_ _03065_ _03068_ _02574_ vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__a2bb2o_1
X_07181_ _03837_ _03838_ vssd1 vssd1 vccd1 vccd1 _03839_ sky130_fd_sc_hd__and2_1
XANTENNA__05683__B2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06132_ _03003_ vssd1 vssd1 vccd1 vccd1 _03004_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_57_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_117_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06063_ net1041 net141 net137 vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__a21o_1
XANTENNA__06005__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout405 net406 vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__buf_2
Xfanout438 _02505_ vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__clkbuf_4
X_09822_ net738 net578 vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__and2_1
Xfanout427 net428 vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__clkbuf_2
Xfanout416 _02759_ vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__clkbuf_4
Xfanout449 _02418_ vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__buf_2
X_09753_ net740 net580 vssd1 vssd1 vccd1 vccd1 _00367_ sky130_fd_sc_hd__and2_1
XANTENNA__09316__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08704_ _04127_ _04129_ vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout282_A _04198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06965_ top.findLeastValue.val2\[1\] net149 net122 _03624_ vssd1 vssd1 vccd1 vccd1
+ _01943_ sky130_fd_sc_hd__o22a_1
X_05916_ _02760_ _02848_ _02850_ _02885_ vssd1 vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__and4_1
X_09684_ net799 net639 vssd1 vssd1 vccd1 vccd1 _00298_ sky130_fd_sc_hd__and2_1
X_06896_ top.compVal\[35\] top.findLeastValue.val1\[35\] net165 vssd1 vssd1 vccd1
+ vccd1 _03590_ sky130_fd_sc_hd__mux2_1
X_08635_ top.cb_syn.cb_length\[3\] _04844_ vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__and2_1
XANTENNA__09840__A net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05847_ top.compVal\[20\] net168 net154 top.WB.CPU_DAT_O\[20\] vssd1 vssd1 vccd1
+ vccd1 _02295_ sky130_fd_sc_hd__a22o_1
XFILLER_42_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout168_X net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08566_ net1113 top.cb_syn.char_path_n\[10\] net221 vssd1 vssd1 vccd1 vccd1 _01528_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07517_ _04102_ _04107_ _04069_ vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__mux2_1
X_05778_ top.findLeastValue.least2\[6\] top.findLeastValue.least2\[5\] top.findLeastValue.least2\[4\]
+ top.findLeastValue.least2\[7\] vssd1 vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__or4b_1
XANTENNA__09051__S net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08497_ net1160 top.cb_syn.char_path_n\[79\] net223 vssd1 vssd1 vccd1 vccd1 _01597_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07448_ top.dut.bit_buf\[0\] net38 net722 vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__mux2_1
XANTENNA__07663__A2 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07379_ _02494_ net153 net127 _03983_ vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__a2bb2o_1
X_09118_ net460 net423 _02937_ vssd1 vssd1 vccd1 vccd1 _05135_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_79_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10390_ net757 net597 vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__and2_1
XFILLER_2_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09049_ net1298 top.WB.CPU_DAT_O\[8\] net293 vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_92_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold470 _01838_ vssd1 vssd1 vccd1 vccd1 net1423 sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 top.path\[37\] vssd1 vssd1 vccd1 vccd1 net1434 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07179__A1 _03817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold492 _01823_ vssd1 vssd1 vccd1 vccd1 net1445 sky130_fd_sc_hd__dlygate4sd3_1
X_11011_ clknet_leaf_11_clk _01559_ _00366_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input10_A DAT_I[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07887__C1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06154__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11844_ clknet_leaf_115_clk _02360_ _01199_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07351__B2 top.findLeastValue.sum\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11775_ clknet_leaf_65_clk _02308_ _01130_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.write_counter_FLV\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10726_ clknet_leaf_113_clk _01325_ _00145_ vssd1 vssd1 vccd1 vccd1 top.path\[102\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_110_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_101_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10657_ clknet_leaf_116_clk _01256_ _00076_ vssd1 vssd1 vccd1 vccd1 top.path\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05665__B2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload26 clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 clkload26/Y sky130_fd_sc_hd__inv_8
Xclkload15 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 clkload15/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload48 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 clkload48/Y sky130_fd_sc_hd__inv_8
Xclkload59 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 clkload59/Y sky130_fd_sc_hd__clkinv_1
Xclkload37 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 clkload37/Y sky130_fd_sc_hd__clkinv_2
X_10588_ net747 net587 vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__and2_1
XANTENNA__09925__A net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11209_ clknet_leaf_6_clk _01757_ _00564_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[111\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05517__X _02619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08975__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06750_ _03526_ _03527_ _03528_ _03533_ vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__nand4_1
X_05701_ net12 net417 net359 top.WB.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1 _02357_
+ sky130_fd_sc_hd__a22o_1
X_06681_ _02442_ top.findLeastValue.val2\[7\] top.findLeastValue.val2\[6\] _02443_
+ vssd1 vssd1 vccd1 vccd1 _03469_ sky130_fd_sc_hd__o22a_1
X_08420_ top.cb_syn.char_path_n\[41\] net391 net330 top.cb_syn.char_path_n\[42\] net508
+ vssd1 vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_47_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05632_ _02713_ _02714_ vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__or2_1
X_05563_ top.cb_syn.char_path\[83\] net551 net542 top.cb_syn.char_path\[51\] vssd1
+ vssd1 vccd1 vccd1 _02657_ sky130_fd_sc_hd__a22o_1
X_08351_ net513 top.cb_syn.char_path_n\[71\] vssd1 vssd1 vccd1 vccd1 _04710_ sky130_fd_sc_hd__or2_1
X_08282_ top.cb_syn.char_path_n\[28\] net207 _04668_ vssd1 vssd1 vccd1 vccd1 _01674_
+ sky130_fd_sc_hd__o21a_1
X_05494_ net456 top.hTree.node_reg\[63\] net362 net422 top.hTree.node_reg\[31\] vssd1
+ vssd1 vccd1 vccd1 _02600_ sky130_fd_sc_hd__a32o_1
XANTENNA__07645__A2 _04199_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07302_ net1716 net273 net268 _03934_ vssd1 vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__a22o_1
XFILLER_20_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_07233_ _03669_ _03877_ vssd1 vssd1 vccd1 vccd1 _03883_ sky130_fd_sc_hd__nand2_1
Xclkload9 clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clkload9/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_119_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout128_A net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07164_ _03821_ vssd1 vssd1 vccd1 vccd1 _03822_ sky130_fd_sc_hd__inv_2
X_06115_ top.cb_syn.char_index\[6\] _02963_ vssd1 vssd1 vccd1 vccd1 _02987_ sky130_fd_sc_hd__or2_1
X_07095_ _03752_ vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__inv_2
XANTENNA__07802__C1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06046_ net530 _02935_ _02936_ net1564 vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout497_A top.findLeastValue.histo_index\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08358__B1 top.cb_syn.end_cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout202 net203 vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__buf_2
Xfanout246 _04538_ vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__clkbuf_2
Xfanout235 _04805_ vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__buf_2
XFILLER_86_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout224 _04805_ vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09046__S net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09554__B net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07997_ top.cb_syn.count\[2\] _02514_ _02515_ top.cb_syn.count\[1\] _04499_ vssd1
+ vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__a221o_1
X_09805_ net791 net631 vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout285_X net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout257 _04190_ vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__buf_2
Xfanout279 _04198_ vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout664_A net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout268 net269 vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__buf_2
XANTENNA_input2_A DAT_I[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09736_ net770 net610 vssd1 vssd1 vccd1 vccd1 _00350_ sky130_fd_sc_hd__and2_1
XANTENNA__05592__B1 _02681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06948_ top.compVal\[9\] top.findLeastValue.val1\[9\] net164 vssd1 vssd1 vccd1 vccd1
+ _03616_ sky130_fd_sc_hd__mux2_1
X_09667_ net780 net620 vssd1 vssd1 vccd1 vccd1 _00281_ sky130_fd_sc_hd__and2_1
XANTENNA__09322__A2 _05255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08618_ top.cb_syn.num_lefts\[7\] _04834_ vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout452_X net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout831_A net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_06879_ top.findLeastValue.val2\[44\] net150 net123 _03581_ vssd1 vssd1 vccd1 vccd1
+ _01986_ sky130_fd_sc_hd__o22a_1
X_09598_ net850 net690 vssd1 vssd1 vccd1 vccd1 _00212_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout717_X net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08549_ net1108 top.cb_syn.char_path_n\[27\] net231 vssd1 vssd1 vccd1 vccd1 _01545_
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_11560_ clknet_leaf_37_clk _02108_ _00915_ vssd1 vssd1 vccd1 vccd1 top.header_synthesis.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06844__B1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05647__B2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10511_ net827 net667 vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__and2_1
X_11491_ clknet_leaf_97_clk _02039_ _00846_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[31\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_108_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10442_ net754 net594 vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__and2_1
XFILLER_40_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10373_ net855 net695 vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__and2_1
XANTENNA__07495__S1 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout780 net786 vssd1 vssd1 vccd1 vccd1 net780 sky130_fd_sc_hd__clkbuf_2
XFILLER_92_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout791 net806 vssd1 vssd1 vccd1 vccd1 net791 sky130_fd_sc_hd__clkbuf_2
XANTENNA__05583__B1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11827_ clknet_leaf_100_clk _02343_ _01182_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_11758_ clknet_leaf_115_clk _02291_ _01113_ vssd1 vssd1 vccd1 vccd1 top.compVal\[16\]
+ sky130_fd_sc_hd__dfrtp_2
X_10709_ clknet_leaf_1_clk _01308_ _00128_ vssd1 vssd1 vccd1 vccd1 top.path\[85\]
+ sky130_fd_sc_hd__dfrtp_1
X_11689_ clknet_leaf_62_clk _02222_ _01044_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload104 clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 clkload104/Y sky130_fd_sc_hd__clkinv_4
Xclkload115 clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 clkload115/Y sky130_fd_sc_hd__inv_6
XANTENNA__06850__A3 _03547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07159__B _03782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07486__S1 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07920_ top.findLeastValue.sum\[4\] _04441_ net395 vssd1 vssd1 vccd1 vccd1 _04442_
+ sky130_fd_sc_hd__mux2_1
X_07851_ net483 _04385_ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__or2_1
XANTENNA__05574__B1 _02666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07782_ net430 _04330_ _04331_ net263 vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__o211a_1
Xinput2 DAT_I[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
X_06802_ top.findLeastValue.val1\[28\] net129 net113 net1699 vssd1 vssd1 vccd1 vccd1
+ _02036_ sky130_fd_sc_hd__o22a_1
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06733_ _03500_ _03504_ _03520_ vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__a21o_1
X_09521_ net740 net580 vssd1 vssd1 vccd1 vccd1 _00135_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_65_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09452_ net848 net688 vssd1 vssd1 vccd1 vccd1 _00066_ sky130_fd_sc_hd__and2_1
XFILLER_51_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06664_ _02409_ top.findLeastValue.val2\[41\] _03449_ _03451_ vssd1 vssd1 vccd1 vccd1
+ _03452_ sky130_fd_sc_hd__a211o_1
XANTENNA__09068__A1 top.CB_write_complete vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08403_ top.cb_syn.char_path_n\[17\] net392 net331 top.cb_syn.char_path_n\[18\] net506
+ vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__a221o_1
X_09383_ net405 _04266_ vssd1 vssd1 vccd1 vccd1 _05266_ sky130_fd_sc_hd__nand2_1
X_06595_ top.compVal\[24\] top.findLeastValue.val1\[24\] vssd1 vssd1 vccd1 vccd1 _03384_
+ sky130_fd_sc_hd__xor2_1
X_05615_ top.histogram.sram_out\[11\] net363 net419 top.hTree.node_reg\[11\] vssd1
+ vssd1 vccd1 vccd1 _02701_ sky130_fd_sc_hd__a22o_1
X_05546_ top.cb_syn.char_path\[22\] net559 net314 top.cb_syn.char_path\[118\] vssd1
+ vssd1 vccd1 vccd1 _02643_ sky130_fd_sc_hd__a22o_1
X_08334_ top.cb_syn.char_path_n\[2\] net202 _04694_ vssd1 vssd1 vccd1 vccd1 _01648_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__05629__B2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05477_ net450 top.histogram.wr_r_en\[1\] net366 _02580_ _02584_ vssd1 vssd1 vccd1
+ vccd1 _02585_ sky130_fd_sc_hd__a311o_1
X_08265_ top.cb_syn.char_path_n\[37\] net380 net339 top.cb_syn.char_path_n\[35\] net184
+ vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__a221o_1
X_07216_ _03853_ _03856_ _03867_ vssd1 vssd1 vccd1 vccd1 _03871_ sky130_fd_sc_hd__nand3_1
X_08196_ top.cb_syn.char_path_n\[71\] net200 _04625_ vssd1 vssd1 vccd1 vccd1 _01717_
+ sky130_fd_sc_hd__o21a_1
X_07147_ _03803_ _03804_ vssd1 vssd1 vccd1 vccd1 _03805_ sky130_fd_sc_hd__and2_1
XFILLER_106_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout879_A net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout781_A net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07078_ _03735_ vssd1 vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__inv_2
X_06029_ net1707 top.WB.CPU_DAT_O\[6\] net355 vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__mux2_1
XFILLER_59_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05565__B1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10991_ clknet_leaf_23_clk _01539_ _00346_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_62_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09719_ net758 net598 vssd1 vssd1 vccd1 vccd1 _00333_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_87_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09059__A1 _03270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11612_ clknet_leaf_63_clk _02160_ _00967_ vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__dfrtp_1
XFILLER_43_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06817__B1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11543_ clknet_leaf_0_clk _02091_ _00898_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11474_ clknet_leaf_99_clk _02022_ _00829_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[14\]
+ sky130_fd_sc_hd__dfstp_1
X_10425_ net874 net714 vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__and2_1
X_10356_ net874 net714 vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__and2_1
XANTENNA__07793__A1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08990__A0 top.WB.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07707__B _04271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10287_ net724 net564 vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__and2_1
XFILLER_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xteam_05_893 vssd1 vssd1 vccd1 vccd1 team_05_893/HI gpio_out[8] sky130_fd_sc_hd__conb_1
Xteam_05_882 vssd1 vssd1 vccd1 vccd1 team_05_882/HI ADR_O[27] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_49_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05556__B1 _02651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05859__B2 top.WB.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05400_ top.cb_syn.char_index\[0\] vssd1 vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__inv_2
XANTENNA__07869__S net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06380_ net1436 _03224_ net300 vssd1 vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05331_ top.compVal\[10\] vssd1 vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__inv_2
XANTENNA__06808__B1 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06074__A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08050_ net439 _04543_ net246 vssd1 vssd1 vccd1 vccd1 _04544_ sky130_fd_sc_hd__a21oi_1
XFILLER_115_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10308__B net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07001_ top.findLeastValue.val1\[44\] top.findLeastValue.val2\[44\] vssd1 vssd1 vccd1
+ vccd1 _03659_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_112_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08430__C1 _02504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08981__A0 top.WB.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08952_ top.WB.CPU_DAT_O\[21\] net1542 net370 vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__mux2_1
X_08883_ top.sram_interface.TRN_counter\[2\] _05054_ _05056_ _02563_ vssd1 vssd1 vccd1
+ vccd1 _01461_ sky130_fd_sc_hd__a22o_1
X_07903_ net442 net1433 net252 top.findLeastValue.sum\[8\] _04428_ vssd1 vssd1 vccd1
+ vccd1 _01813_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_71_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07834_ top.findLeastValue.sum\[21\] top.hTree.tree_reg\[21\] net278 vssd1 vssd1
+ vccd1 vccd1 _04373_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout195_A net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05547__B1 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06948__S net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout362_A _02583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07765_ top.findLeastValue.sum\[35\] _04317_ net396 vssd1 vssd1 vccd1 vccd1 _04318_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07696_ net491 _04259_ vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__or2_1
X_06716_ _03494_ _03503_ _03489_ vssd1 vssd1 vccd1 vccd1 _03504_ sky130_fd_sc_hd__a21oi_1
X_09504_ net759 net599 vssd1 vssd1 vccd1 vccd1 _00118_ sky130_fd_sc_hd__and2_1
X_09435_ net1027 vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__clkbuf_1
X_06647_ top.compVal\[39\] top.compVal\[38\] top.compVal\[37\] top.compVal\[36\] vssd1
+ vssd1 vccd1 vccd1 _03436_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout627_A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout248_X net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07779__S net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout150_X net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09366_ net984 net243 net218 _04322_ vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__a22o_1
X_06578_ _03364_ _03365_ _03366_ vssd1 vssd1 vccd1 vccd1 _03367_ sky130_fd_sc_hd__a21o_1
X_09297_ net298 _04007_ vssd1 vssd1 vccd1 vccd1 top.dut.bit_buf_next\[13\] sky130_fd_sc_hd__and2_1
X_05529_ _02627_ _02628_ net476 vssd1 vssd1 vccd1 vccd1 _02629_ sky130_fd_sc_hd__o21a_1
X_08317_ top.cb_syn.char_path_n\[11\] net374 net334 top.cb_syn.char_path_n\[9\] net179
+ vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__a221o_1
X_08248_ top.cb_syn.char_path_n\[45\] net195 _04651_ vssd1 vssd1 vccd1 vccd1 _01691_
+ sky130_fd_sc_hd__o21a_1
X_08179_ top.cb_syn.char_path_n\[80\] net376 net336 top.cb_syn.char_path_n\[78\] net181
+ vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__a221o_1
X_10210_ net826 net666 vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__and2_1
XANTENNA__06027__A1 top.WB.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11190_ clknet_leaf_19_clk _01738_ _00545_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[92\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08972__A0 top.WB.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10141_ net830 net670 vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__and2_1
X_10072_ net863 net703 vssd1 vssd1 vccd1 vccd1 _00686_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_7_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05538__B1 _02636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08639__A net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07543__A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10974_ clknet_leaf_14_clk _01522_ _00329_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06446__X _03269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05710__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09189__B _04188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11526_ clknet_leaf_55_clk _02074_ _00881_ vssd1 vssd1 vccd1 vccd1 top.controller.fin_HG
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10128__B net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11457_ clknet_leaf_69_clk _02005_ _00812_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least2\[7\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__06018__A1 top.WB.CPU_DAT_O\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10408_ net794 net634 vssd1 vssd1 vccd1 vccd1 _01022_ sky130_fd_sc_hd__and2_1
X_11388_ clknet_leaf_83_clk _01936_ _00743_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[40\]
+ sky130_fd_sc_hd__dfrtp_1
X_10339_ net794 net634 vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__and2_1
XFILLER_3_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08963__A0 top.WB.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09933__A net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05529__B1 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05880_ _02855_ _02856_ vssd1 vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__nor2_1
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05525__X _02626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07550_ _04140_ _04138_ _04137_ _04131_ vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__and4b_1
XANTENNA__07740__X _04298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06501_ net1531 _03306_ _03282_ vssd1 vssd1 vccd1 vccd1 _02089_ sky130_fd_sc_hd__o21ba_1
XANTENNA__08983__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09220_ _05191_ vssd1 vssd1 vccd1 vccd1 _00014_ sky130_fd_sc_hd__inv_2
X_07481_ _04054_ _04058_ vssd1 vssd1 vccd1 vccd1 _04072_ sky130_fd_sc_hd__xor2_4
XFILLER_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06432_ top.header_synthesis.count\[7\] top.header_synthesis.count\[6\] top.header_synthesis.count\[5\]
+ top.header_synthesis.count\[4\] vssd1 vssd1 vccd1 vccd1 _03259_ sky130_fd_sc_hd__or4_1
XANTENNA__05701__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09151_ _02937_ _05110_ top.sram_interface.word_cnt\[13\] vssd1 vssd1 vccd1 vccd1
+ _05158_ sky130_fd_sc_hd__o21a_1
X_06363_ top.hist_data_o\[19\] _03187_ vssd1 vssd1 vccd1 vccd1 _03214_ sky130_fd_sc_hd__xor2_1
XANTENNA__08246__A2 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_8_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09082_ top.histogram.eof_n top.dut.out_valid _03320_ net295 net449 vssd1 vssd1 vccd1
+ vccd1 _05103_ sky130_fd_sc_hd__a41o_1
X_08102_ top.cb_syn.char_path_n\[118\] net204 _04578_ vssd1 vssd1 vccd1 vccd1 _01764_
+ sky130_fd_sc_hd__o21a_1
X_05314_ top.compVal\[28\] vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_32_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08033_ _04527_ vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__inv_2
X_06294_ top.cb_syn.max_index\[1\] _03025_ _03027_ top.hTree.nullSumIndex\[0\] vssd1
+ vssd1 vccd1 vccd1 _03159_ sky130_fd_sc_hd__a22o_1
XANTENNA__06008__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout208_A net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06009__A1 top.WB.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08954__A0 top.WB.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09984_ net803 net643 vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__and2_1
XFILLER_103_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08935_ top.WB.CPU_DAT_O\[19\] net1347 net371 vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout577_A net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08866_ _02789_ _05042_ vssd1 vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__or2_1
X_07817_ net427 _04358_ _04359_ net259 vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__o211a_1
XANTENNA__09054__S net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08797_ top.path\[30\] top.path\[31\] net525 vssd1 vssd1 vccd1 vccd1 _04980_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout365_X net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout744_A net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07748_ net443 net1533 net255 top.findLeastValue.sum\[39\] _04304_ vssd1 vssd1 vccd1
+ vccd1 _01844_ sky130_fd_sc_hd__a221o_1
XANTENNA__05940__A0 top.WB.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07679_ net263 _04247_ _04248_ net1022 net446 vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__a32o_1
XFILLER_13_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_09418_ net407 _04211_ vssd1 vssd1 vccd1 vccd1 _05289_ sky130_fd_sc_hd__nand2_1
X_10690_ clknet_leaf_112_clk _01289_ _00109_ vssd1 vssd1 vccd1 vccd1 top.path\[66\]
+ sky130_fd_sc_hd__dfrtp_1
X_09349_ net1025 net238 net216 _04390_ vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__a22o_1
X_11311_ clknet_leaf_77_clk _01859_ _00666_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06799__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08641__B net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11242_ clknet_leaf_32_clk _01790_ _00597_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_95_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08945__A0 top.WB.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11173_ clknet_leaf_3_clk _01721_ _00528_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[75\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_input40_A gpio_in[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10124_ net839 net679 vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__and2_1
XFILLER_88_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10055_ net846 net686 vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__and2_1
XFILLER_87_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05931__A0 top.WB.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10957_ clknet_leaf_65_clk net954 _00312_ vssd1 vssd1 vccd1 vccd1 top.controller.fin_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10888_ clknet_leaf_111_clk _01465_ _00243_ vssd1 vssd1 vccd1 vccd1 top.translation.index\[3\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_8_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold107 net55 vssd1 vssd1 vccd1 vccd1 net1060 sky130_fd_sc_hd__dlygate4sd3_1
X_11509_ clknet_leaf_70_clk _02057_ _00864_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least1\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_8_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xhold129 top.path\[94\] vssd1 vssd1 vccd1 vccd1 net1082 sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 top.hTree.node_reg\[11\] vssd1 vssd1 vccd1 vccd1 net1071 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08936__A0 top.WB.CPU_DAT_O\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout609 net612 vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07735__X _04294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06981_ top.findLeastValue.val2\[34\] top.findLeastValue.val2\[33\] top.findLeastValue.val2\[32\]
+ top.findLeastValue.val2\[31\] vssd1 vssd1 vccd1 vccd1 _03639_ sky130_fd_sc_hd__and4_1
X_08720_ top.cb_syn.i\[2\] top.cb_syn.i\[1\] top.cb_syn.i\[0\] top.cb_syn.i\[3\] vssd1
+ vssd1 vccd1 vccd1 _04909_ sky130_fd_sc_hd__a31o_1
X_05932_ top.WB.CPU_DAT_O\[23\] net1257 net304 vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__mux2_1
X_08651_ _04563_ _04801_ _04857_ vssd1 vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__and3_1
XANTENNA__09361__B1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05863_ top.compVal\[4\] net170 net157 top.WB.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1
+ _02279_ sky130_fd_sc_hd__a22o_1
X_07602_ net1475 _04186_ _04144_ vssd1 vssd1 vccd1 vccd1 _01872_ sky130_fd_sc_hd__mux2_1
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_08582_ top.cb_syn.h_element\[60\] top.cb_syn.h_element\[51\] net533 vssd1 vssd1
+ vccd1 vccd1 _04810_ sky130_fd_sc_hd__mux2_1
X_05794_ top.sram_interface.counter_HTREE\[0\] top.hTree.state\[2\] _02805_ _02813_
+ top.WorR vssd1 vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_37_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07533_ _04054_ _04070_ net402 vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__nand3_1
XFILLER_81_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07464_ top.cb_syn.i\[1\] top.cb_syn.cb_length\[1\] vssd1 vssd1 vccd1 vccd1 _04055_
+ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_17_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06415_ _02540_ top.header_synthesis.start _03245_ vssd1 vssd1 vccd1 vccd1 _03246_
+ sky130_fd_sc_hd__a21boi_1
X_09203_ _02809_ _04188_ _05177_ net489 vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__a22o_1
X_07395_ _03996_ vssd1 vssd1 vccd1 vccd1 top.dut.bits_in_buf_next\[2\] sky130_fd_sc_hd__inv_2
X_09134_ net468 top.sram_interface.word_cnt\[7\] _02776_ _05144_ net548 vssd1 vssd1
+ vccd1 vccd1 _05146_ sky130_fd_sc_hd__a32o_1
XFILLER_108_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07522__S0 _04072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06346_ top.hist_data_o\[26\] _03197_ _03192_ vssd1 vssd1 vccd1 vccd1 _03204_ sky130_fd_sc_hd__o21ba_1
X_09065_ top.hist_addr\[2\] _05090_ _05091_ top.TRN_char_index\[2\] vssd1 vssd1 vccd1
+ vccd1 _01250_ sky130_fd_sc_hd__a22o_1
X_06277_ net561 _02563_ top.TRN_char_index\[0\] vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout113_X net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08016_ _04507_ _04518_ _04509_ vssd1 vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__a21o_1
XANTENNA__09049__S net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold630 top.hTree.tree_reg\[0\] vssd1 vssd1 vccd1 vccd1 net1583 sky130_fd_sc_hd__dlygate4sd3_1
Xhold641 top.hist_data_o\[28\] vssd1 vssd1 vccd1 vccd1 net1594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold652 top.hist_data_o\[24\] vssd1 vssd1 vccd1 vccd1 net1605 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08927__A0 top.WB.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold663 top.histogram.total\[13\] vssd1 vssd1 vccd1 vccd1 net1616 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold696 top.dut.out\[0\] vssd1 vssd1 vccd1 vccd1 net1649 sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 top.cb_syn.i\[4\] vssd1 vssd1 vccd1 vccd1 net1638 sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 top.findLeastValue.sum\[40\] vssd1 vssd1 vccd1 vccd1 net1627 sky130_fd_sc_hd__dlygate4sd3_1
X_09967_ net778 net618 vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout861_A net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08918_ _05072_ top.cb_syn.max_index\[2\] vssd1 vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__nand2b_1
XFILLER_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06953__A2 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09898_ net782 net622 vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__and2_1
XANTENNA__09352__B1 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08849_ top.translation.index\[6\] _05031_ _04976_ vssd1 vssd1 vccd1 vccd1 _05032_
+ sky130_fd_sc_hd__o21ba_1
XFILLER_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11860_ clknet_leaf_115_clk _02376_ _01215_ vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__dfrtp_1
X_11791_ clknet_leaf_72_clk _00026_ _01146_ vssd1 vssd1 vccd1 vccd1 top.hTree.state\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10811_ clknet_leaf_83_clk _01397_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_10742_ clknet_leaf_2_clk _01341_ _00161_ vssd1 vssd1 vccd1 vccd1 top.path\[118\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10955__Q top.controller.fin_reg\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06156__B net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10673_ clknet_leaf_122_clk _01272_ _00092_ vssd1 vssd1 vccd1 vccd1 top.path\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05692__A2 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05444__A2 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11225_ clknet_leaf_27_clk _01773_ _00580_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[127\]
+ sky130_fd_sc_hd__dfrtp_1
X_11156_ clknet_leaf_25_clk _01704_ _00511_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08394__B2 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11087_ clknet_leaf_23_clk _01635_ _00442_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[117\]
+ sky130_fd_sc_hd__dfrtp_1
X_10107_ net819 net659 vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__and2_1
X_10038_ net837 net677 vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_106_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06992__D top.findLeastValue.val1\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_50_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08854__C1 top.controller.state_reg\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06200_ _02572_ _03004_ _03066_ _02550_ net500 vssd1 vssd1 vccd1 vccd1 _03069_ sky130_fd_sc_hd__a32o_1
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07180_ _03672_ _03836_ _03675_ _03674_ vssd1 vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__o211a_1
XANTENNA__05683__A2 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06131_ top.cw2\[5\] top.cw2\[4\] _03001_ vssd1 vssd1 vccd1 vccd1 _03003_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_65_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07504__S0 _04072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06062_ net1052 net142 net137 vssd1 vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_57_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout439 _02498_ vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkload12_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout406 net407 vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__buf_2
Xfanout428 _02535_ vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__buf_2
XANTENNA__08385__B2 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09821_ net738 net578 vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__and2_1
Xfanout417 net418 vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08501__S net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09752_ net758 net598 vssd1 vssd1 vccd1 vccd1 _00366_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_123_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08703_ net439 _04895_ _04894_ vssd1 vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__mux2_1
XFILLER_104_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__08137__A1 top.cb_syn.char_path_n\[101\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06964_ top.compVal\[1\] top.findLeastValue.val1\[1\] net164 vssd1 vssd1 vccd1 vccd1
+ _03624_ sky130_fd_sc_hd__mux2_1
X_05915_ top.sram_interface.init_counter\[10\] _02582_ _02884_ top.sram_interface.init_counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02886_ sky130_fd_sc_hd__or4b_1
X_09683_ net799 net639 vssd1 vssd1 vccd1 vccd1 _00297_ sky130_fd_sc_hd__and2_1
XFILLER_104_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout275_A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06895_ top.findLeastValue.val2\[36\] net151 net123 _03589_ vssd1 vssd1 vccd1 vccd1
+ _01978_ sky130_fd_sc_hd__o22a_1
XANTENNA__06021__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08634_ _04844_ vssd1 vssd1 vccd1 vccd1 _04845_ sky130_fd_sc_hd__inv_2
XANTENNA__09840__B net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06956__S net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05846_ top.compVal\[21\] net168 net154 top.WB.CPU_DAT_O\[21\] vssd1 vssd1 vccd1
+ vccd1 _02296_ sky130_fd_sc_hd__a22o_1
XANTENNA__07641__A net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05777_ top.findLeastValue.least2\[3\] top.findLeastValue.least2\[2\] top.findLeastValue.least2\[1\]
+ top.findLeastValue.least2\[0\] vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__or4_1
X_08565_ net1216 top.cb_syn.char_path_n\[11\] net220 vssd1 vssd1 vccd1 vccd1 _01529_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07516_ _04103_ _04104_ _04105_ _04106_ _04072_ _04071_ vssd1 vssd1 vccd1 vccd1 _04107_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout442_A net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_18_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08496_ net1158 top.cb_syn.char_path_n\[80\] net223 vssd1 vssd1 vccd1 vccd1 _01598_
+ sky130_fd_sc_hd__mux2_1
X_07447_ net1623 top.dut.out_valid_next _04002_ _04021_ _04040_ vssd1 vssd1 vccd1
+ vccd1 _01881_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout707_A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06871__B2 top.findLeastValue.histo_index\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07378_ top.cw1\[0\] _03423_ _03553_ top.findLeastValue.histo_index\[0\] vssd1 vssd1
+ vccd1 vccd1 _03983_ sky130_fd_sc_hd__a22o_1
X_09117_ _02570_ _05134_ _05087_ vssd1 vssd1 vccd1 vccd1 _00046_ sky130_fd_sc_hd__or3b_1
X_06329_ top.hist_data_o\[26\] top.hist_data_o\[25\] _03191_ vssd1 vssd1 vccd1 vccd1
+ _03192_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_79_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09048_ net1277 top.WB.CPU_DAT_O\[9\] net293 vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout697_X net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold460 net68 vssd1 vssd1 vccd1 vccd1 net1413 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold471 top.hTree.node_reg\[20\] vssd1 vssd1 vccd1 vccd1 net1424 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08411__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08376__B2 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold482 top.path\[60\] vssd1 vssd1 vccd1 vccd1 net1435 sky130_fd_sc_hd__dlygate4sd3_1
Xhold493 top.path\[73\] vssd1 vssd1 vccd1 vccd1 net1446 sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ clknet_leaf_11_clk _01558_ _00365_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_57_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09089__C1 _02581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11843_ clknet_leaf_116_clk _02359_ _01198_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_14_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11774_ clknet_leaf_65_clk _02307_ _01129_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.write_counter_FLV\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10725_ clknet_leaf_112_clk _01324_ _00144_ vssd1 vssd1 vccd1 vccd1 top.path\[101\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10656_ clknet_leaf_114_clk _01255_ _00075_ vssd1 vssd1 vccd1 vccd1 top.path\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05665__A2 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload16 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 clkload16/Y sky130_fd_sc_hd__inv_6
XANTENNA__06075__C1 _02949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload49 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 clkload49/Y sky130_fd_sc_hd__inv_6
Xclkload38 clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 clkload38/Y sky130_fd_sc_hd__clkinv_2
Xclkload27 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 clkload27/Y sky130_fd_sc_hd__inv_8
X_10587_ net746 net586 vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__and2_1
XANTENNA__09925__B net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08367__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11208_ clknet_leaf_6_clk _01756_ _00563_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[110\]
+ sky130_fd_sc_hd__dfrtp_1
X_11139_ clknet_leaf_11_clk _01687_ _00494_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[41\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_36_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05700_ net14 net415 net308 top.WB.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 _02358_
+ sky130_fd_sc_hd__o22a_1
X_06680_ _03465_ _03466_ _03467_ vssd1 vssd1 vccd1 vccd1 _03468_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_19_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05631_ top.cb_syn.char_path\[8\] net558 net313 top.cb_syn.char_path\[104\] vssd1
+ vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__a22o_1
X_08350_ top.cb_syn.char_path_n\[65\] top.cb_syn.char_path_n\[66\] top.cb_syn.char_path_n\[67\]
+ top.cb_syn.char_path_n\[68\] net513 net509 vssd1 vssd1 vccd1 vccd1 _04709_ sky130_fd_sc_hd__mux4_1
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05562_ net1261 net139 _02656_ net175 vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__a22o_1
X_07301_ _03923_ _03933_ vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__nor2_1
X_08281_ top.cb_syn.char_path_n\[29\] net385 net344 top.cb_syn.char_path_n\[27\] net189
+ vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__a221o_1
X_05493_ net462 net550 vssd1 vssd1 vccd1 vccd1 _02599_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_63_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08842__A2 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07232_ net271 _03879_ _03882_ net276 net1659 vssd1 vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_119_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07163_ top.findLeastValue.val1\[34\] top.findLeastValue.val2\[34\] vssd1 vssd1 vccd1
+ vccd1 _03821_ sky130_fd_sc_hd__nand2_1
X_06114_ top.TRN_char_index\[6\] _02977_ _02985_ vssd1 vssd1 vccd1 vccd1 _02986_ sky130_fd_sc_hd__o21a_1
XANTENNA__06016__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07094_ top.findLeastValue.val1\[0\] top.findLeastValue.val2\[0\] _03750_ vssd1 vssd1
+ vccd1 vccd1 _03752_ sky130_fd_sc_hd__and3_1
X_06045_ net536 _02935_ vssd1 vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__nand2_1
Xfanout203 net211 vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout214 net215 vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__buf_2
X_09804_ net790 net630 vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout392_A net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout225 net226 vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__clkbuf_4
Xfanout247 net249 vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__clkbuf_4
Xfanout236 net237 vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__buf_2
X_07996_ top.cb_syn.count\[1\] _02515_ _02516_ top.cb_syn.count\[0\] vssd1 vssd1 vccd1
+ vccd1 _04499_ sky130_fd_sc_hd__o22a_1
Xfanout269 _03864_ vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__clkbuf_4
Xfanout258 net259 vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__buf_2
X_09735_ net771 net611 vssd1 vssd1 vccd1 vccd1 _00349_ sky130_fd_sc_hd__and2_1
XANTENNA__05592__B2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06947_ top.findLeastValue.val2\[10\] net147 net121 _03615_ vssd1 vssd1 vccd1 vccd1
+ _01952_ sky130_fd_sc_hd__o22a_1
X_09666_ net803 net643 vssd1 vssd1 vccd1 vccd1 _00280_ sky130_fd_sc_hd__and2_1
XFILLER_67_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout278_X net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout657_A net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08617_ net439 _02527_ _04834_ _04826_ vssd1 vssd1 vccd1 vccd1 _04836_ sky130_fd_sc_hd__a31o_1
X_06878_ top.compVal\[44\] top.findLeastValue.val1\[44\] net165 vssd1 vssd1 vccd1
+ vccd1 _03581_ sky130_fd_sc_hd__mux2_1
X_09597_ net851 net691 vssd1 vssd1 vccd1 vccd1 _00211_ sky130_fd_sc_hd__and2_1
X_05829_ _02838_ _02841_ vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout445_X net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout824_A net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08548_ net1164 top.cb_syn.char_path_n\[28\] net231 vssd1 vssd1 vccd1 vccd1 _01546_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout612_X net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08479_ net1266 top.cb_syn.char_path_n\[97\] net234 vssd1 vssd1 vccd1 vccd1 _01615_
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_25_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05647__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10510_ net816 net656 vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__and2_1
X_11490_ clknet_leaf_81_clk _02038_ _00845_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[30\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_109_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10441_ net847 net687 vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__and2_1
XANTENNA__08597__A1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10372_ net854 net694 vssd1 vssd1 vccd1 vccd1 _00986_ sky130_fd_sc_hd__and2_1
XANTENNA__06285__A1_N net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08349__A1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold290 net84 vssd1 vssd1 vccd1 vccd1 net1243 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout781 net786 vssd1 vssd1 vccd1 vccd1 net781 sky130_fd_sc_hd__buf_1
Xfanout770 net771 vssd1 vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__clkbuf_2
Xfanout792 net806 vssd1 vssd1 vccd1 vccd1 net792 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06780__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ clknet_leaf_115_clk _02342_ _01181_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_60_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11757_ clknet_leaf_101_clk _02290_ _01112_ vssd1 vssd1 vccd1 vccd1 top.compVal\[15\]
+ sky130_fd_sc_hd__dfrtp_4
X_10708_ clknet_leaf_2_clk _01307_ _00127_ vssd1 vssd1 vccd1 vccd1 top.path\[84\]
+ sky130_fd_sc_hd__dfrtp_1
X_11688_ clknet_leaf_62_clk _02221_ _01043_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload105 clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 clkload105/Y sky130_fd_sc_hd__bufinv_16
Xclkload116 clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 clkload116/Y sky130_fd_sc_hd__inv_8
X_10639_ clknet_leaf_74_clk _00048_ _00058_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.word_cnt\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09936__A net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07850_ top.findLeastValue.sum\[18\] _04385_ net395 vssd1 vssd1 vccd1 vccd1 _04386_
+ sky130_fd_sc_hd__mux2_1
XFILLER_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07563__A2 _04144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07781_ net490 _04329_ vssd1 vssd1 vccd1 vccd1 _04331_ sky130_fd_sc_hd__or2_1
X_06801_ top.findLeastValue.val1\[29\] net129 net113 net1669 vssd1 vssd1 vccd1 vccd1
+ _02037_ sky130_fd_sc_hd__o22a_1
XANTENNA__07890__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05574__B2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput3 DAT_I[10] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
X_06732_ _03516_ _03518_ _03519_ vssd1 vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__or3_1
X_09520_ net740 net580 vssd1 vssd1 vccd1 vccd1 _00134_ sky130_fd_sc_hd__and2_1
XFILLER_83_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_09451_ net848 net688 vssd1 vssd1 vccd1 vccd1 _00065_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_65_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06663_ top.compVal\[42\] _02483_ _03450_ vssd1 vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__o21ai_1
X_08402_ top.cb_syn.char_path_n\[19\] top.cb_syn.char_path_n\[20\] net515 vssd1 vssd1
+ vccd1 vccd1 _04761_ sky130_fd_sc_hd__mux2_1
X_09382_ net992 net240 _05264_ _05265_ vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__a22o_1
X_06594_ _02423_ top.findLeastValue.val1\[27\] top.findLeastValue.val1\[26\] _02424_
+ _03333_ vssd1 vssd1 vccd1 vccd1 _03383_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05614_ _02698_ _02699_ net472 vssd1 vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__o21a_1
X_05545_ top.cb_syn.char_path\[86\] net553 net544 top.cb_syn.char_path\[54\] vssd1
+ vssd1 vccd1 vccd1 _02642_ sky130_fd_sc_hd__a22o_1
X_08333_ top.cb_syn.char_path_n\[3\] net381 net340 net517 net185 vssd1 vssd1 vccd1
+ vccd1 _04694_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout140_A _02595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08371__S0 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08264_ top.cb_syn.char_path_n\[37\] net201 _04659_ vssd1 vssd1 vccd1 vccd1 _01683_
+ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout238_A net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05629__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05476_ top.sram_interface.word_cnt\[5\] top.sram_interface.word_cnt\[13\] net362
+ net459 vssd1 vssd1 vccd1 vccd1 _02584_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout405_A net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10057__A net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08195_ top.cb_syn.char_path_n\[72\] net379 net338 top.cb_syn.char_path_n\[70\] net183
+ vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__a221o_1
XFILLER_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07215_ net271 _03869_ _03870_ net276 net1703 vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__a32o_1
X_07146_ top.findLeastValue.val1\[22\] top.findLeastValue.val2\[22\] vssd1 vssd1 vccd1
+ vccd1 _03804_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_76_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07787__C1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07077_ _03731_ _03733_ _03734_ vssd1 vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__and3_1
XANTENNA__09057__S net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06028_ net1485 top.WB.CPU_DAT_O\[7\] net355 vssd1 vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout774_A net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout395_X net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07979_ net1488 net534 _04482_ vssd1 vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__mux2_1
X_09718_ net742 net582 vssd1 vssd1 vccd1 vccd1 _00332_ sky130_fd_sc_hd__and2_1
X_10990_ clknet_leaf_23_clk _01538_ _00345_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09649_ net780 net620 vssd1 vssd1 vccd1 vccd1 _00263_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_87_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ clknet_leaf_64_clk _02159_ _00966_ vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_116_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_116_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_42_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11542_ clknet_leaf_0_clk _02090_ _00897_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_109_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11473_ clknet_leaf_99_clk _02021_ _00828_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[13\]
+ sky130_fd_sc_hd__dfstp_1
X_10424_ net873 net713 vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__and2_1
XANTENNA__08660__A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10355_ net872 net712 vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__and2_1
X_10286_ net726 net566 vssd1 vssd1 vccd1 vccd1 _00900_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_29_Left_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xteam_05_894 vssd1 vssd1 vccd1 vccd1 team_05_894/HI gpio_out[9] sky130_fd_sc_hd__conb_1
Xteam_05_883 vssd1 vssd1 vccd1 vccd1 team_05_883/HI ADR_O[30] sky130_fd_sc_hd__conb_1
XANTENNA__05556__B2 _02589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_1_Left_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11809_ clknet_leaf_97_clk _02326_ _01164_ vssd1 vssd1 vccd1 vccd1 top.compVal\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_38_Left_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_107_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_107_clk
+ sky130_fd_sc_hd__clkbuf_8
X_05330_ top.compVal\[11\] vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_60_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06284__A2 _02767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06074__B net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05492__B1 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07000_ net287 _03657_ vssd1 vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__and2_2
XANTENNA__06090__A top.cb_syn.char_index\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08951_ top.WB.CPU_DAT_O\[22\] top.cb_syn.h_element\[54\] net370 vssd1 vssd1 vccd1
+ vccd1 _01359_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_47_Left_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08882_ _02891_ _05055_ _05054_ vssd1 vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__a21oi_1
X_07902_ net427 _04426_ _04427_ net259 vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__o211a_1
XFILLER_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_clkbuf_4_4_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07833_ net441 net1588 net253 top.findLeastValue.sum\[22\] _04372_ vssd1 vssd1 vccd1
+ vccd1 _01827_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout188_A net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07764_ top.findLeastValue.sum\[35\] top.hTree.tree_reg\[35\] net280 vssd1 vssd1
+ vccd1 vccd1 _04317_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07695_ net491 _04261_ vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__nand2_1
XFILLER_52_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06715_ _03495_ _03502_ _03491_ vssd1 vssd1 vccd1 vccd1 _03503_ sky130_fd_sc_hd__a21o_1
X_09503_ net749 net589 vssd1 vssd1 vccd1 vccd1 _00117_ sky130_fd_sc_hd__and2_1
X_09434_ net1017 vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_56_Left_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06964__S net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06646_ top.compVal\[43\] top.compVal\[42\] top.compVal\[41\] top.compVal\[40\] vssd1
+ vssd1 vccd1 vccd1 _03435_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout355_A net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout143_X net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09365_ net1006 net240 net216 _04326_ vssd1 vssd1 vccd1 vccd1 _01427_ sky130_fd_sc_hd__a22o_1
X_06577_ _02441_ top.findLeastValue.val1\[8\] top.findLeastValue.val1\[7\] _02442_
+ vssd1 vssd1 vccd1 vccd1 _03366_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout522_A top.translation.index\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09296_ net298 _04003_ vssd1 vssd1 vccd1 vccd1 top.dut.bit_buf_next\[12\] sky130_fd_sc_hd__and2_1
X_05528_ top.cb_syn.char_path\[25\] net559 net314 top.cb_syn.char_path\[121\] vssd1
+ vssd1 vccd1 vccd1 _02628_ sky130_fd_sc_hd__a22o_1
X_08316_ top.cb_syn.char_path_n\[11\] net196 _04685_ vssd1 vssd1 vccd1 vccd1 _01657_
+ sky130_fd_sc_hd__o21a_1
X_05459_ net495 _02418_ vssd1 vssd1 vccd1 vccd1 _02567_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08247_ top.cb_syn.char_path_n\[46\] net373 net333 top.cb_syn.char_path_n\[44\] net178
+ vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__a221o_1
XANTENNA__07795__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout408_X net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_106_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_EDGE_ROW_65_Left_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08178_ top.cb_syn.char_path_n\[80\] net202 _04616_ vssd1 vssd1 vccd1 vccd1 _01726_
+ sky130_fd_sc_hd__o21a_1
XFILLER_97_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07129_ top.findLeastValue.val1\[18\] top.findLeastValue.val2\[18\] vssd1 vssd1 vccd1
+ vccd1 _03787_ sky130_fd_sc_hd__or2_1
X_10140_ net830 net670 vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__and2_1
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10071_ net850 net690 vssd1 vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_7_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06983__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05538__B2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07543__B net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold734_A top.findLeastValue.sum\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10958__Q top.controller.fin_reg\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_74_Left_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10973_ clknet_leaf_15_clk _01521_ _00328_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09250__S net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05710__B2 top.WB.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11525_ clknet_leaf_66_clk _02073_ _00880_ vssd1 vssd1 vccd1 vccd1 top.controller.fin_FLV
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09204__A2 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11456_ clknet_leaf_71_clk _02004_ _00811_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least2\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08412__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10407_ net792 net632 vssd1 vssd1 vccd1 vccd1 _01021_ sky130_fd_sc_hd__and2_1
X_11387_ clknet_leaf_87_clk _01935_ _00742_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05487__A_N net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10338_ net794 net634 vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__and2_1
XANTENNA__09933__B net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10269_ net735 net575 vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__and2_1
XFILLER_93_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07480_ _04059_ _04070_ vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__xnor2_4
X_06500_ top.histogram.total\[13\] top.histogram.total\[12\] _03281_ vssd1 vssd1 vccd1
+ vccd1 _03306_ sky130_fd_sc_hd__and3_1
XANTENNA__05541__X _02639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06431_ net1495 _03258_ _03254_ vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__o21a_1
XANTENNA__05701__B2 top.WB.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09150_ net459 net546 top.sram_interface.word_cnt\[2\] net468 _05157_ vssd1 vssd1
+ vccd1 vccd1 _00041_ sky130_fd_sc_hd__a221o_1
X_06362_ net1138 _03213_ net302 vssd1 vssd1 vccd1 vccd1 _02135_ sky130_fd_sc_hd__mux2_1
X_06293_ _03020_ _03157_ top.histogram.init vssd1 vssd1 vccd1 vccd1 _03158_ sky130_fd_sc_hd__a21o_1
X_09081_ _02568_ _05101_ vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__nor2_1
X_08101_ top.cb_syn.char_path_n\[119\] net383 net342 top.cb_syn.char_path_n\[117\]
+ net187 vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__a221o_1
X_05313_ top.compVal\[29\] vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_32_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08032_ top.cb_syn.end_cond top.CB_write_complete vssd1 vssd1 vccd1 vccd1 _04527_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_116_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__08403__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_09983_ net785 net625 vssd1 vssd1 vccd1 vccd1 _00597_ sky130_fd_sc_hd__and2_1
XFILLER_89_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07757__A2 _04310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06024__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08934_ top.WB.CPU_DAT_O\[20\] net1296 net371 vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__mux2_1
XANTENNA__06965__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08167__C1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout472_A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08865_ _02519_ _02789_ _05040_ vssd1 vssd1 vccd1 vccd1 _05045_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08182__A2 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07816_ net484 _04357_ vssd1 vssd1 vccd1 vccd1 _04359_ sky130_fd_sc_hd__or2_1
X_08796_ top.path\[24\] net408 _04978_ vssd1 vssd1 vccd1 vccd1 _04979_ sky130_fd_sc_hd__o21a_1
X_07747_ net429 _04302_ _04303_ net261 vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout737_A net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07678_ net489 _04244_ vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09417_ net990 net242 _05287_ _05288_ vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_51_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06629_ top.compVal\[38\] _02463_ _03404_ _03417_ _03395_ vssd1 vssd1 vccd1 vccd1
+ _03418_ sky130_fd_sc_hd__o221a_1
X_09348_ net997 net238 net216 _04394_ vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__a22o_1
XFILLER_8_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09279_ _05228_ _05229_ vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_zero_count\[6\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__08922__B net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11310_ clknet_leaf_77_clk _01858_ _00665_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_113_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_11241_ clknet_leaf_30_clk _01789_ _00596_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10245__A net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11172_ clknet_leaf_3_clk _01720_ _00527_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[74\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_106_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_10123_ net840 net680 vssd1 vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__and2_1
XFILLER_0_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05759__B2 top.WB.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10054_ net837 net677 vssd1 vssd1 vccd1 vccd1 _00668_ sky130_fd_sc_hd__and2_1
XANTENNA_input33_A DAT_I[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_82_Left_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08173__A2 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09370__B2 _04306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__09122__A1 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10956_ clknet_leaf_40_clk net956 _00311_ vssd1 vssd1 vccd1 vccd1 top.controller.fin_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10887_ clknet_leaf_111_clk _01464_ _00242_ vssd1 vssd1 vccd1 vccd1 top.translation.index\[2\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_91_Left_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold108 top.WB.curr_state\[2\] vssd1 vssd1 vccd1 vccd1 net1061 sky130_fd_sc_hd__dlygate4sd3_1
X_11508_ clknet_leaf_69_clk _02056_ _00863_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least1\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_8_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold119 top.path\[10\] vssd1 vssd1 vccd1 vccd1 net1072 sky130_fd_sc_hd__dlygate4sd3_1
X_11439_ clknet_leaf_89_clk _01987_ _00794_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[45\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__08397__C1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06947__B1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06980_ top.findLeastValue.val2\[38\] top.findLeastValue.val2\[37\] top.findLeastValue.val2\[36\]
+ top.findLeastValue.val2\[35\] vssd1 vssd1 vccd1 vccd1 _03638_ sky130_fd_sc_hd__and4_1
XANTENNA__05536__X _02635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05931_ top.WB.CPU_DAT_O\[24\] net1364 net305 vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__mux2_1
XFILLER_39_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08650_ top.cb_syn.cb_length\[0\] top.cb_syn.cb_length\[1\] vssd1 vssd1 vccd1 vccd1
+ _04857_ sky130_fd_sc_hd__nand2b_1
XANTENNA__08164__A2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05862_ top.compVal\[5\] net170 net156 top.WB.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1
+ _02280_ sky130_fd_sc_hd__a22o_1
X_07601_ net532 top.cb_syn.h_element\[46\] _04184_ _04185_ vssd1 vssd1 vccd1 vccd1
+ _04186_ sky130_fd_sc_hd__a211o_1
XFILLER_66_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08581_ _04809_ top.cb_syn.char_index\[6\] _04807_ vssd1 vssd1 vccd1 vccd1 _01516_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09113__A1 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05793_ _02459_ _02473_ vssd1 vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_37_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07532_ _04044_ _04045_ _04048_ _04057_ vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__or4b_1
X_07463_ _04052_ _04053_ vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_17_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_06414_ top.header_synthesis.write_num_lefts top.header_synthesis.write_char_path
+ vssd1 vssd1 vccd1 vccd1 _03245_ sky130_fd_sc_hd__or2_2
X_09202_ top.hTree.state\[3\] net264 _05162_ net1698 vssd1 vssd1 vccd1 vccd1 _00020_
+ sky130_fd_sc_hd__a22o_1
X_07394_ top.dut.bits_in_buf\[2\] _03984_ net403 net722 vssd1 vssd1 vccd1 vccd1 _03996_
+ sky130_fd_sc_hd__a22oi_4
X_09133_ net469 net562 top.sram_interface.word_cnt\[2\] net460 _02564_ vssd1 vssd1
+ vccd1 vccd1 _05145_ sky130_fd_sc_hd__a221o_1
XANTENNA__09416__A2 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06019__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06345_ net1259 _03203_ net303 vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__mux2_1
XANTENNA__08742__B top.TRN_sram_complete vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout220_A net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09064_ net1637 _05090_ _05091_ top.TRN_char_index\[3\] vssd1 vssd1 vccd1 vccd1 _01251_
+ sky130_fd_sc_hd__a22o_1
X_06276_ _02943_ _03140_ _03141_ net495 net467 vssd1 vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__o221a_1
XANTENNA__07522__S1 _04071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold620 top.cb_syn.zeroes\[3\] vssd1 vssd1 vccd1 vccd1 net1573 sky130_fd_sc_hd__dlygate4sd3_1
X_08015_ top.cb_syn.count\[6\] _04516_ vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__nand2_1
XFILLER_89_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xhold653 top.hTree.tree_reg\[38\] vssd1 vssd1 vccd1 vccd1 net1606 sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 top.hTree.tree_reg\[5\] vssd1 vssd1 vccd1 vccd1 net1584 sky130_fd_sc_hd__dlygate4sd3_1
Xhold642 top.hTree.tree_reg\[13\] vssd1 vssd1 vccd1 vccd1 net1595 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout687_A net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold686 top.findLeastValue.sum\[35\] vssd1 vssd1 vccd1 vccd1 net1639 sky130_fd_sc_hd__dlygate4sd3_1
Xhold675 top.compVal\[16\] vssd1 vssd1 vccd1 vccd1 net1628 sky130_fd_sc_hd__dlygate4sd3_1
Xhold664 _03307_ vssd1 vssd1 vccd1 vccd1 net1617 sky130_fd_sc_hd__dlygate4sd3_1
Xhold697 top.translation.totalEn vssd1 vssd1 vccd1 vccd1 net1650 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09966_ net778 net618 vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__and2_1
XANTENNA__07645__Y _04221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06402__A2 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09897_ net775 net615 vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__and2_1
X_08917_ top.cb_syn.max_index\[3\] _05082_ _05072_ vssd1 vssd1 vccd1 vccd1 _01389_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__08155__A2 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_96_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_96_clk sky130_fd_sc_hd__clkbuf_8
X_08848_ _05024_ _05030_ top.translation.index\[5\] vssd1 vssd1 vccd1 vccd1 _05031_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07363__B1 _03553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08779_ top.path\[121\] net328 _04961_ vssd1 vssd1 vccd1 vccd1 _04962_ sky130_fd_sc_hd__o21a_1
X_11790_ clknet_leaf_72_clk _00025_ _01145_ vssd1 vssd1 vccd1 vccd1 top.hTree.state\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10810_ clknet_leaf_83_clk _01396_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07666__A1 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07666__B2 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10741_ clknet_leaf_2_clk _01340_ _00160_ vssd1 vssd1 vccd1 vccd1 top.path\[117\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05677__B1 _02752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09407__A2 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10672_ clknet_leaf_122_clk _01271_ _00091_ vssd1 vssd1 vccd1 vccd1 top.path\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_20_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07513__S1 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11224_ clknet_leaf_28_clk _01772_ _00579_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[126\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_4_12_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08379__C1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11155_ clknet_leaf_26_clk _01703_ _00510_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08394__A2 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11086_ clknet_leaf_23_clk _01634_ _00441_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[116\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input36_X net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10106_ net812 net652 vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__and2_1
XANTENNA__07284__A _03782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10037_ net837 net677 vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_87_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10939_ clknet_leaf_35_clk _01494_ _00294_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.cb_length\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_44_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06634__Y _03423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_11_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_8
X_06130_ top.cw2\[4\] _03001_ vssd1 vssd1 vccd1 vccd1 _03002_ sky130_fd_sc_hd__nand2_1
XANTENNA__07504__S1 _04071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06061_ net1044 net141 net137 vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__a21o_1
XANTENNA__06093__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05840__B1 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout418 _02758_ vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__buf_2
Xfanout407 _02808_ vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__clkbuf_4
Xfanout429 net430 vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__buf_2
X_09820_ net735 net575 vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__and2_1
XFILLER_100_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06963_ top.findLeastValue.val2\[2\] net149 net122 _03623_ vssd1 vssd1 vccd1 vccd1
+ _01944_ sky130_fd_sc_hd__o22a_1
XANTENNA__08790__C1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09751_ net762 net602 vssd1 vssd1 vccd1 vccd1 _00365_ sky130_fd_sc_hd__and2_1
X_05914_ top.sram_interface.init_counter\[1\] top.sram_interface.init_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02885_ sky130_fd_sc_hd__nor2_1
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08702_ _02457_ _04536_ top.cb_syn.left_check vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__a21boi_1
Xclkbuf_leaf_78_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_clk sky130_fd_sc_hd__clkbuf_8
X_09682_ net797 net637 vssd1 vssd1 vccd1 vccd1 _00296_ sky130_fd_sc_hd__and2_1
XANTENNA__07481__X _04072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06894_ top.compVal\[36\] top.findLeastValue.val1\[36\] net165 vssd1 vssd1 vccd1
+ vccd1 _03589_ sky130_fd_sc_hd__mux2_1
X_08633_ top.cb_syn.cb_length\[2\] top.cb_syn.cb_length\[1\] top.cb_syn.cb_length\[0\]
+ _04563_ vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_68_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout170_A net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05845_ top.compVal\[22\] net168 net154 top.WB.CPU_DAT_O\[22\] vssd1 vssd1 vccd1
+ vccd1 _02297_ sky130_fd_sc_hd__a22o_1
X_05776_ top.findLeastValue.least1\[8\] _02795_ vssd1 vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout268_A net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08564_ net1143 top.cb_syn.char_path_n\[12\] net220 vssd1 vssd1 vccd1 vccd1 _01530_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__05442__A net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07515_ top.cb_syn.char_path_n\[80\] top.cb_syn.char_path_n\[79\] top.cb_syn.char_path_n\[78\]
+ top.cb_syn.char_path_n\[77\] net399 net350 vssd1 vssd1 vccd1 vccd1 _04106_ sky130_fd_sc_hd__mux4_1
XANTENNA__07648__B2 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08495_ net1281 top.cb_syn.char_path_n\[81\] net223 vssd1 vssd1 vccd1 vccd1 _01599_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__05659__B1 _02737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07446_ net354 top.dut.bits_in_buf_next\[0\] _04034_ _04039_ vssd1 vssd1 vccd1 vccd1
+ _04040_ sky130_fd_sc_hd__a31o_1
X_07377_ top.cw2\[1\] net134 _03547_ net127 _03982_ vssd1 vssd1 vccd1 vccd1 _01889_
+ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout602_A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09116_ net555 _05132_ _05133_ net541 vssd1 vssd1 vccd1 vccd1 _05134_ sky130_fd_sc_hd__a22o_1
X_06328_ top.hist_data_o\[24\] top.hist_data_o\[23\] _03190_ vssd1 vssd1 vccd1 vccd1
+ _03191_ sky130_fd_sc_hd__and3_1
X_09047_ net1072 top.WB.CPU_DAT_O\[10\] net293 vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__mux2_1
X_06259_ _02559_ _03123_ _03124_ _03125_ _03121_ vssd1 vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_79_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09584__A net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold450 top.hTree.tree_reg\[29\] vssd1 vssd1 vccd1 vccd1 net1403 sky130_fd_sc_hd__dlygate4sd3_1
Xhold472 top.path\[2\] vssd1 vssd1 vccd1 vccd1 net1425 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09022__A0 top.WB.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold461 top.path\[88\] vssd1 vssd1 vccd1 vccd1 net1414 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08376__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold494 top.path\[105\] vssd1 vssd1 vccd1 vccd1 net1447 sky130_fd_sc_hd__dlygate4sd3_1
Xhold483 top.histogram.sram_out\[13\] vssd1 vssd1 vccd1 vccd1 net1436 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07562__B1_N _04144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09949_ net738 net578 vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__and2_1
XANTENNA__08781__C1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout857_X net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_69_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08759__S0 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11842_ clknet_leaf_117_clk _02358_ _01197_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_33_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10966__Q top.cb_syn.char_index\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07639__A1 top.findLeastValue.least1\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11773_ clknet_leaf_103_clk _02306_ _01128_ vssd1 vssd1 vccd1 vccd1 top.compVal\[31\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_110_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10724_ clknet_leaf_112_clk _01323_ _00143_ vssd1 vssd1 vccd1 vccd1 top.path\[100\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06882__S net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10655_ clknet_leaf_59_clk _01254_ _00074_ vssd1 vssd1 vccd1 vccd1 top.hist_addr\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07498__S0 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload17 clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 clkload17/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__11797__Q top.controller.state_reg\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06075__B1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload39 clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 clkload39/Y sky130_fd_sc_hd__clkinv_2
Xclkload28 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 clkload28/Y sky130_fd_sc_hd__clkinv_2
XFILLER_5_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10586_ net746 net586 vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__and2_1
XFILLER_119_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__05822__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09013__A0 top.WB.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11207_ clknet_leaf_6_clk _01755_ _00562_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[109\]
+ sky130_fd_sc_hd__dfrtp_2
X_11138_ clknet_leaf_12_clk _01686_ _00493_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[40\]
+ sky130_fd_sc_hd__dfrtp_2
X_11069_ clknet_leaf_16_clk _01617_ _00424_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[99\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_0_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07327__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07878__B2 top.findLeastValue.sum\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05630_ top.cb_syn.char_path\[72\] net552 net543 top.cb_syn.char_path\[40\] vssd1
+ vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__a22o_1
XANTENNA__10876__Q top.cb_syn.curr_state\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09095__A3 _02899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05561_ top.histogram.sram_out\[20\] net364 _02654_ _02655_ vssd1 vssd1 vccd1 vccd1
+ _02656_ sky130_fd_sc_hd__a211o_1
X_07300_ _03794_ _03813_ _03922_ vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__and3_1
X_08280_ top.cb_syn.char_path_n\[29\] net206 _04667_ vssd1 vssd1 vccd1 vccd1 _01675_
+ sky130_fd_sc_hd__o21a_1
X_05492_ _02596_ _02597_ net477 vssd1 vssd1 vccd1 vccd1 _02598_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_63_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07231_ _03663_ _03878_ vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_119_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07162_ _03704_ _03816_ _03818_ _03819_ vssd1 vssd1 vccd1 vccd1 _03820_ sky130_fd_sc_hd__o211a_1
XANTENNA__06066__B1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06113_ top.TRN_char_index\[6\] _02977_ _02560_ vssd1 vssd1 vccd1 vccd1 _02985_ sky130_fd_sc_hd__a21oi_1
XFILLER_105_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07093_ top.findLeastValue.val1\[0\] top.findLeastValue.val2\[0\] vssd1 vssd1 vccd1
+ vccd1 _03751_ sky130_fd_sc_hd__nand2_1
X_06044_ _02457_ net517 _02934_ vssd1 vssd1 vccd1 vccd1 _02935_ sky130_fd_sc_hd__o21a_1
XANTENNA__08512__S net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09004__A0 top.WB.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout204 net211 vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__buf_2
XFILLER_115_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09803_ net783 net623 vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__and2_1
Xfanout226 net228 vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__clkbuf_4
Xfanout215 net217 vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__buf_2
Xfanout237 net239 vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__buf_1
X_07995_ top.cb_syn.count\[2\] _02514_ vssd1 vssd1 vccd1 vccd1 _04498_ sky130_fd_sc_hd__or2_1
Xfanout248 net249 vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__clkbuf_4
Xfanout259 net261 vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__clkbuf_4
X_09734_ net770 net610 vssd1 vssd1 vccd1 vccd1 _00348_ sky130_fd_sc_hd__and2_1
XFILLER_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05592__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06946_ top.compVal\[10\] top.findLeastValue.val1\[10\] net162 vssd1 vssd1 vccd1
+ vccd1 _03615_ sky130_fd_sc_hd__mux2_1
X_09665_ net784 net624 vssd1 vssd1 vccd1 vccd1 _00279_ sky130_fd_sc_hd__and2_1
XANTENNA__07652__A net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout552_A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06877_ top.findLeastValue.val2\[45\] net150 net125 _03580_ vssd1 vssd1 vccd1 vccd1
+ _01987_ sky130_fd_sc_hd__o22a_1
X_08616_ _04826_ _02527_ net439 vssd1 vssd1 vccd1 vccd1 _04835_ sky130_fd_sc_hd__and3b_2
X_05828_ top.sram_interface.write_counter_FLV\[0\] net289 net1635 vssd1 vssd1 vccd1
+ vccd1 _02841_ sky130_fd_sc_hd__a21oi_1
X_09596_ net851 net691 vssd1 vssd1 vccd1 vccd1 _00210_ sky130_fd_sc_hd__and2_1
X_08547_ net1076 top.cb_syn.char_path_n\[29\] net232 vssd1 vssd1 vccd1 vccd1 _01547_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout438_X net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_05759_ top.compVal\[35\] net172 net158 top.WB.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1
+ _02320_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout817_A net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08478_ net1359 top.cb_syn.char_path_n\[98\] net233 vssd1 vssd1 vccd1 vccd1 _01616_
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07429_ top.dut.bit_buf\[4\] net42 net720 vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__mux2_1
XANTENNA__05501__C1 _02605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10440_ net860 net700 vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__and2_1
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06057__B1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10371_ net855 net695 vssd1 vssd1 vccd1 vccd1 _00985_ sky130_fd_sc_hd__and2_1
Xhold280 top.cb_syn.char_path\[99\] vssd1 vssd1 vccd1 vccd1 net1233 sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 top.path\[107\] vssd1 vssd1 vccd1 vccd1 net1244 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout760 net762 vssd1 vssd1 vccd1 vccd1 net760 sky130_fd_sc_hd__clkbuf_2
Xfanout782 net786 vssd1 vssd1 vccd1 vccd1 net782 sky130_fd_sc_hd__clkbuf_2
Xfanout771 net772 vssd1 vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06780__A1 top.findLeastValue.least1\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout793 net806 vssd1 vssd1 vccd1 vccd1 net793 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_92_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05634__X _02717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_64_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06532__A1 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11825_ clknet_leaf_100_clk _02341_ _01180_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_26_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11756_ clknet_leaf_99_clk _02289_ _01111_ vssd1 vssd1 vccd1 vccd1 top.compVal\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10707_ clknet_leaf_4_clk _01306_ _00126_ vssd1 vssd1 vccd1 vccd1 top.path\[83\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_79_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11687_ clknet_leaf_62_clk _02220_ _01042_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_122_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06048__B1 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload106 clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 clkload106/Y sky130_fd_sc_hd__inv_6
Xclkload117 clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 clkload117/Y sky130_fd_sc_hd__clkinv_8
X_10638_ clknet_leaf_58_clk net1103 _00057_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.word_cnt\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09936__B net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10569_ net752 net592 vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_114_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_17_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05574__A2 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07780_ top.hTree.tree_reg\[32\] top.findLeastValue.sum\[32\] net250 vssd1 vssd1
+ vccd1 vccd1 _04330_ sky130_fd_sc_hd__mux2_1
X_06800_ top.findLeastValue.val1\[30\] net129 net113 top.compVal\[30\] vssd1 vssd1
+ vccd1 vccd1 _02038_ sky130_fd_sc_hd__o22a_1
Xinput4 DAT_I[11] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
X_06731_ top.compVal\[25\] _02488_ _02489_ top.compVal\[24\] _03513_ vssd1 vssd1 vccd1
+ vccd1 _03519_ sky130_fd_sc_hd__a221o_1
X_09450_ net867 net707 vssd1 vssd1 vccd1 vccd1 _00064_ sky130_fd_sc_hd__and2_1
XANTENNA__06088__A top.cb_syn.char_index\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08401_ net508 _04751_ _04754_ _04759_ top.cb_syn.end_cnt\[4\] vssd1 vssd1 vccd1
+ vccd1 _04760_ sky130_fd_sc_hd__a311oi_2
X_06662_ _02408_ top.findLeastValue.val2\[43\] vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__nand2_1
X_09381_ top.hTree.nulls\[47\] net405 net244 vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__o21a_1
XFILLER_51_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06593_ _03352_ _03379_ _03380_ _03381_ vssd1 vssd1 vccd1 vccd1 _03382_ sky130_fd_sc_hd__a31o_1
X_05613_ top.cb_syn.char_path\[11\] net557 net312 top.cb_syn.char_path\[107\] vssd1
+ vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__a22o_1
X_05544_ net1354 net140 _02641_ net176 vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__a22o_1
X_08332_ top.cb_syn.char_path_n\[3\] net201 _04693_ vssd1 vssd1 vccd1 vccd1 _01649_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__06287__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08371__S1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08263_ top.cb_syn.char_path_n\[38\] net380 net339 top.cb_syn.char_path_n\[36\] net184
+ vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_22_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05475_ top.WorR _02536_ vssd1 vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__nor2_1
XFILLER_20_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_0_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07214_ _03851_ _03868_ _03850_ vssd1 vssd1 vccd1 vccd1 _03870_ sky130_fd_sc_hd__a21o_1
XANTENNA__10057__B net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08194_ top.cb_syn.char_path_n\[72\] net200 _04624_ vssd1 vssd1 vccd1 vccd1 _01718_
+ sky130_fd_sc_hd__o21a_1
XFILLER_106_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout300_A net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07145_ top.findLeastValue.val1\[22\] top.findLeastValue.val2\[22\] vssd1 vssd1 vccd1
+ vccd1 _03803_ sky130_fd_sc_hd__nand2_1
XANTENNA__09320__S0 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07076_ top.findLeastValue.val1\[9\] top.findLeastValue.val2\[9\] vssd1 vssd1 vccd1
+ vccd1 _03734_ sky130_fd_sc_hd__or2_1
X_06027_ net1618 top.WB.CPU_DAT_O\[8\] net355 vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__mux2_1
XFILLER_59_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07978_ _02932_ _04142_ _04481_ vssd1 vssd1 vccd1 vccd1 _04482_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout767_A net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09717_ net760 net600 vssd1 vssd1 vccd1 vccd1 _00331_ sky130_fd_sc_hd__and2_1
X_06929_ top.findLeastValue.val2\[19\] net146 net120 _03606_ vssd1 vssd1 vccd1 vccd1
+ _01961_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout555_X net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09648_ net780 net620 vssd1 vssd1 vccd1 vccd1 _00262_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_87_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09579_ net819 net659 vssd1 vssd1 vccd1 vccd1 _00193_ sky130_fd_sc_hd__and2_1
X_11610_ clknet_leaf_69_clk _02158_ _00965_ vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__dfrtp_1
XFILLER_30_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08417__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11541_ clknet_leaf_0_clk _02089_ _00896_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06817__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11472_ clknet_leaf_99_clk _02020_ _00827_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[12\]
+ sky130_fd_sc_hd__dfstp_1
X_10423_ net873 net713 vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__and2_1
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11140__Q top.cb_syn.char_path_n\[42\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10354_ net874 net714 vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__and2_1
XFILLER_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10285_ net725 net565 vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__and2_1
XANTENNA__06202__B1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_05_895 vssd1 vssd1 vccd1 vccd1 team_05_895/HI gpio_out[10] sky130_fd_sc_hd__conb_1
Xteam_05_884 vssd1 vssd1 vccd1 vccd1 team_05_884/HI ADR_O[31] sky130_fd_sc_hd__conb_1
XANTENNA__07950__A0 top.findLeastValue.least1\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05556__A2 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout590 net597 vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__clkbuf_2
XFILLER_93_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_clkload9_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11808_ clknet_leaf_90_clk _02325_ _01163_ vssd1 vssd1 vccd1 vccd1 top.compVal\[40\]
+ sky130_fd_sc_hd__dfrtp_2
X_11739_ clknet_leaf_66_clk _02272_ _01094_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.zero_cnt\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06808__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08430__A1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_102_Left_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08950_ top.WB.CPU_DAT_O\[23\] top.cb_syn.h_element\[55\] net369 vssd1 vssd1 vccd1
+ vccd1 _01360_ sky130_fd_sc_hd__mux2_1
XFILLER_102_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08881_ top.sram_interface.TRN_counter\[1\] top.sram_interface.TRN_counter\[0\] top.sram_interface.TRN_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05055_ sky130_fd_sc_hd__a21bo_1
X_07901_ net484 _04425_ vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__or2_1
XFILLER_111_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07832_ net428 _04370_ _04371_ net262 vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__o211a_1
X_07763_ net443 net1401 net255 top.findLeastValue.sum\[36\] _04316_ vssd1 vssd1 vccd1
+ vccd1 _01841_ sky130_fd_sc_hd__a221o_1
X_09502_ net750 net590 vssd1 vssd1 vccd1 vccd1 _00116_ sky130_fd_sc_hd__and2_1
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07694_ _02477_ net396 _04260_ vssd1 vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__o21a_1
X_06714_ _03488_ _03498_ _03501_ _02492_ top.compVal\[20\] vssd1 vssd1 vccd1 vccd1
+ _03502_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_27_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09433_ net959 vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_fanout250_A _04199_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06645_ _03430_ _03431_ _03433_ vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_111_Left_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout348_A net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09364_ net982 net242 net218 _04330_ vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__a22o_1
XFILLER_24_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05450__A net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06576_ _02442_ top.findLeastValue.val1\[7\] top.findLeastValue.val1\[6\] _02443_
+ vssd1 vssd1 vccd1 vccd1 _03365_ sky130_fd_sc_hd__o22a_1
X_08315_ top.cb_syn.char_path_n\[12\] net374 net334 top.cb_syn.char_path_n\[10\] net179
+ vssd1 vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__a221o_1
X_09295_ net298 _04004_ vssd1 vssd1 vccd1 vccd1 top.dut.bit_buf_next\[11\] sky130_fd_sc_hd__and2_1
X_05527_ top.cb_syn.char_path\[89\] net553 net544 top.cb_syn.char_path\[57\] vssd1
+ vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout515_A top.cb_syn.end_cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout136_X net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05458_ _02560_ _02565_ vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__nand2_1
XANTENNA__09857__A net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08246_ top.cb_syn.char_path_n\[46\] net196 _04650_ vssd1 vssd1 vccd1 vccd1 _01692_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__08761__A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08177_ top.cb_syn.char_path_n\[81\] net382 net341 top.cb_syn.char_path_n\[79\] net186
+ vssd1 vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__a221o_1
X_05389_ top.cb_syn.check_right vssd1 vssd1 vccd1 vccd1 _02497_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout303_X net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07128_ top.findLeastValue.val1\[18\] top.findLeastValue.val2\[18\] vssd1 vssd1 vccd1
+ vccd1 _03786_ sky130_fd_sc_hd__nand2_1
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08421__A1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07059_ top.findLeastValue.val1\[13\] top.findLeastValue.val2\[13\] vssd1 vssd1 vccd1
+ vccd1 _03717_ sky130_fd_sc_hd__and2_1
X_10070_ net851 net691 vssd1 vssd1 vccd1 vccd1 _00684_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_7_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_102_Right_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08185__B1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05538__A2 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10972_ clknet_leaf_16_clk _01520_ _00327_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_83_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05710__A2 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11524_ clknet_leaf_59_clk _02072_ _00879_ vssd1 vssd1 vccd1 vccd1 top.cw1\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_7_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06890__S net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11455_ clknet_leaf_71_clk _02003_ _00810_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least2\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_109_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_109_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10406_ net793 net633 vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__and2_1
X_11386_ clknet_leaf_87_clk _01934_ _00741_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_111_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10337_ net794 net634 vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__and2_1
X_10268_ net735 net575 vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__and2_1
X_10199_ net858 net698 vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_109_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06430_ top.header_synthesis.count\[3\] top.header_synthesis.count\[2\] _03256_ vssd1
+ vssd1 vccd1 vccd1 _03258_ sky130_fd_sc_hd__and3_1
XANTENNA__05701__A2 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08852__Y _05035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06361_ _03188_ _03212_ vssd1 vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__nor2_1
X_06292_ top.hist_addr\[1\] top.hist_addr\[0\] vssd1 vssd1 vccd1 vccd1 _03157_ sky130_fd_sc_hd__or2_1
X_09080_ top.histogram.init_edge _05089_ vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__or2_1
XANTENNA__09677__A net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08100_ top.cb_syn.char_path_n\[119\] net204 _04577_ vssd1 vssd1 vccd1 vccd1 _01765_
+ sky130_fd_sc_hd__o21a_1
X_05312_ top.compVal\[30\] vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_32_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput40 gpio_in[6] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__clkbuf_1
X_08031_ _04520_ _04509_ top.cb_syn.count\[0\] vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__mux2_1
XFILLER_116_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_73_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09982_ net781 net621 vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__and2_1
XFILLER_88_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08933_ top.WB.CPU_DAT_O\[21\] net1181 net371 vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__mux2_1
XFILLER_69_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10351__A net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07914__A0 top.findLeastValue.sum\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08864_ _02790_ _05042_ _05044_ _05041_ net1656 vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__o32a_1
XANTENNA__05445__A top.CB_write_complete vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07815_ top.hTree.tree_reg\[25\] top.findLeastValue.sum\[25\] net249 vssd1 vssd1
+ vccd1 vccd1 _04358_ sky130_fd_sc_hd__mux2_1
X_08795_ top.path\[25\] net326 _04977_ net432 net436 vssd1 vssd1 vccd1 vccd1 _04978_
+ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout465_A top.controller.state_reg\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07746_ net488 _04301_ vssd1 vssd1 vccd1 vccd1 _04303_ sky130_fd_sc_hd__or2_1
XFILLER_84_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05732__X _02767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout632_A net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout253_X net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07677_ net489 _04246_ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__nand2_1
X_09416_ top.hTree.nulls\[59\] net407 net245 vssd1 vssd1 vccd1 vccd1 _05288_ sky130_fd_sc_hd__o21a_1
XFILLER_52_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06628_ top.compVal\[36\] _02465_ _03390_ _03416_ _03402_ vssd1 vssd1 vccd1 vccd1
+ _03417_ sky130_fd_sc_hd__o221a_1
X_09347_ net1012 net238 net216 _04398_ vssd1 vssd1 vccd1 vccd1 _01409_ sky130_fd_sc_hd__a22o_1
X_06559_ _03344_ _03345_ _03346_ _03347_ vssd1 vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__o31a_1
X_09278_ _05213_ _05224_ top.cb_syn.zero_count\[6\] vssd1 vssd1 vccd1 vccd1 _05229_
+ sky130_fd_sc_hd__a21o_1
XFILLER_32_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08229_ top.cb_syn.char_path_n\[55\] net384 net343 top.cb_syn.char_path_n\[53\] net188
+ vssd1 vssd1 vccd1 vccd1 _04642_ sky130_fd_sc_hd__a221o_1
X_11240_ clknet_leaf_30_clk _01788_ _00595_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_106_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_95_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11171_ clknet_leaf_11_clk _01719_ _00526_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[73\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_106_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10122_ net840 net680 vssd1 vssd1 vccd1 vccd1 _00736_ sky130_fd_sc_hd__and2_1
XFILLER_95_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07554__B top.cb_syn.h_element\[63\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10053_ net845 net685 vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__and2_1
XANTENNA_input26_A DAT_I[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10955_ clknet_leaf_42_clk top.controller.fin_TRN _00310_ vssd1 vssd1 vccd1 vccd1
+ top.controller.fin_reg\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_73_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10886_ clknet_leaf_110_clk _01463_ _00241_ vssd1 vssd1 vccd1 vccd1 top.translation.index\[1\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__05695__B2 top.WB.CPU_DAT_O\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11507_ clknet_leaf_66_clk _02055_ _00862_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.wipe_the_char_2
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xhold109 top.cb_syn.end_cond vssd1 vssd1 vccd1 vccd1 net1062 sky130_fd_sc_hd__dlygate4sd3_1
X_11438_ clknet_leaf_89_clk _01986_ _00793_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[44\]
+ sky130_fd_sc_hd__dfstp_1
X_11369_ clknet_leaf_102_clk _01917_ _00724_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_05930_ top.WB.CPU_DAT_O\[25\] net1396 net305 vssd1 vssd1 vccd1 vccd1 _02259_ sky130_fd_sc_hd__mux2_1
XFILLER_39_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05861_ top.compVal\[6\] net171 net157 top.WB.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1
+ _02281_ sky130_fd_sc_hd__a22o_1
XFILLER_39_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08580_ top.cb_syn.h_element\[61\] top.cb_syn.h_element\[52\] net533 vssd1 vssd1
+ vccd1 vccd1 _04809_ sky130_fd_sc_hd__mux2_1
X_07600_ top.cb_syn.max_index\[1\] _04135_ _04183_ net537 vssd1 vssd1 vccd1 vccd1
+ _04185_ sky130_fd_sc_hd__a22o_1
X_07531_ top.cb_syn.h_element\[54\] _04121_ vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__nand2b_1
XANTENNA__09113__A2 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05792_ _02806_ _02807_ _02809_ _02811_ vssd1 vssd1 vccd1 vccd1 _02812_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07462_ top.cb_syn.cb_length\[2\] top.cb_syn.i\[2\] vssd1 vssd1 vccd1 vccd1 _04053_
+ sky130_fd_sc_hd__and2b_1
X_07393_ top.dut.bits_in_buf\[0\] top.dut.bits_in_buf\[1\] top.dut.bits_in_buf\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__nor3_1
X_09201_ top.hTree.state\[3\] net257 _05180_ vssd1 vssd1 vccd1 vccd1 _00021_ sky130_fd_sc_hd__a21o_1
X_06413_ _02456_ top.histogram.sram_out\[0\] net299 vssd1 vssd1 vccd1 vccd1 _02115_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09132_ net454 net463 _05112_ vssd1 vssd1 vccd1 vccd1 _05144_ sky130_fd_sc_hd__a21o_1
X_06344_ top.hist_data_o\[27\] _03192_ _03198_ vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__o21ba_1
XFILLER_108_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08515__S net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_06275_ top.hist_addr\[2\] _03020_ vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__xnor2_1
X_09063_ top.hist_addr\[4\] _05090_ _05091_ top.TRN_char_index\[4\] vssd1 vssd1 vccd1
+ vccd1 _01252_ sky130_fd_sc_hd__a22o_1
XANTENNA__07832__C1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08014_ _04516_ vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__inv_2
Xhold621 top.hTree.tree_reg\[15\] vssd1 vssd1 vccd1 vccd1 net1574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold610 _01821_ vssd1 vssd1 vccd1 vccd1 net1563 sky130_fd_sc_hd__dlygate4sd3_1
Xhold643 top.cb_syn.curr_index\[4\] vssd1 vssd1 vccd1 vccd1 net1596 sky130_fd_sc_hd__dlygate4sd3_1
Xhold654 top.hist_data_o\[10\] vssd1 vssd1 vccd1 vccd1 net1607 sky130_fd_sc_hd__dlygate4sd3_1
Xhold632 top.findLeastValue.sum\[42\] vssd1 vssd1 vccd1 vccd1 net1585 sky130_fd_sc_hd__dlygate4sd3_1
Xhold676 top.hTree.nullSumIndex\[4\] vssd1 vssd1 vccd1 vccd1 net1629 sky130_fd_sc_hd__dlygate4sd3_1
Xhold687 top.findLeastValue.sum\[29\] vssd1 vssd1 vccd1 vccd1 net1640 sky130_fd_sc_hd__dlygate4sd3_1
Xhold665 top.hist_data_o\[8\] vssd1 vssd1 vccd1 vccd1 net1618 sky130_fd_sc_hd__dlygate4sd3_1
Xhold698 top.cb_syn.num_lefts\[5\] vssd1 vssd1 vccd1 vccd1 net1651 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09965_ net779 net619 vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout582_A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09896_ net775 net615 vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__and2_1
X_08916_ _04174_ _05081_ vssd1 vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__xor2_1
X_08847_ _05019_ _05029_ _05000_ _04995_ net520 top.translation.index\[4\] vssd1 vssd1
+ vccd1 vccd1 _05030_ sky130_fd_sc_hd__mux4_1
XANTENNA__07363__B2 top.findLeastValue.histo_index\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout847_A net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08778_ top.path\[120\] net410 _04960_ net434 net520 vssd1 vssd1 vccd1 vccd1 _04961_
+ sky130_fd_sc_hd__o221a_1
X_07729_ top.findLeastValue.sum\[42\] top.hTree.tree_reg\[42\] net282 vssd1 vssd1
+ vccd1 vccd1 _04289_ sky130_fd_sc_hd__mux2_1
X_10740_ clknet_leaf_119_clk _01339_ _00159_ vssd1 vssd1 vccd1 vccd1 top.path\[116\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05677__B2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10671_ clknet_leaf_119_clk _01270_ _00090_ vssd1 vssd1 vccd1 vccd1 top.path\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11223_ clknet_leaf_30_clk _01771_ _00578_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[125\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08379__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09040__A1 top.WB.CPU_DAT_O\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11154_ clknet_leaf_26_clk _01702_ _00509_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[56\]
+ sky130_fd_sc_hd__dfrtp_1
X_11085_ clknet_leaf_23_clk _01633_ _00440_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[115\]
+ sky130_fd_sc_hd__dfrtp_1
X_10105_ net819 net659 vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__and2_1
X_10036_ net837 net677 vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__and2_1
XANTENNA__08396__A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10938_ clknet_leaf_34_clk _01493_ _00293_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.cb_length\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07657__A2 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08854__A1 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10869_ clknet_leaf_47_clk _01455_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_14_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06060_ net1060 net141 net137 vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_117_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08909__A2 _04187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__05547__X _02644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09031__A1 top.WB.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05840__B2 top.WB.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout408 _02788_ vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__clkbuf_4
Xfanout419 net421 vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__buf_2
XFILLER_86_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09750_ net760 net600 vssd1 vssd1 vccd1 vccd1 _00364_ sky130_fd_sc_hd__and2_1
X_06962_ top.compVal\[2\] top.findLeastValue.val1\[2\] net164 vssd1 vssd1 vccd1 vccd1
+ _03623_ sky130_fd_sc_hd__mux2_1
X_05913_ top.sram_interface.init_counter\[9\] top.sram_interface.init_counter\[8\]
+ top.sram_interface.init_counter\[7\] top.sram_interface.init_counter\[6\] vssd1
+ vssd1 vccd1 vccd1 _02884_ sky130_fd_sc_hd__or4_1
X_08701_ top.cb_syn.h_element\[63\] _02862_ _04534_ _04893_ vssd1 vssd1 vccd1 vccd1
+ _04894_ sky130_fd_sc_hd__or4_1
X_09681_ net783 net623 vssd1 vssd1 vccd1 vccd1 _00295_ sky130_fd_sc_hd__and2_1
XANTENNA__09334__A2 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08632_ _04835_ _04826_ top.cb_syn.num_lefts\[0\] vssd1 vssd1 vccd1 vccd1 _01499_
+ sky130_fd_sc_hd__mux2_1
X_06893_ top.findLeastValue.val2\[37\] net150 net125 _03588_ vssd1 vssd1 vccd1 vccd1
+ _01979_ sky130_fd_sc_hd__o22a_1
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05844_ top.compVal\[23\] net168 net154 top.WB.CPU_DAT_O\[23\] vssd1 vssd1 vccd1
+ vccd1 _02298_ sky130_fd_sc_hd__a22o_1
XFILLER_82_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05775_ _02793_ _02794_ vssd1 vssd1 vccd1 vccd1 _02795_ sky130_fd_sc_hd__nor2_1
XFILLER_54_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout163_A _03423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08563_ net1180 top.cb_syn.char_path_n\[13\] net220 vssd1 vssd1 vccd1 vccd1 _01531_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__05442__B net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08494_ net1188 top.cb_syn.char_path_n\[82\] net223 vssd1 vssd1 vccd1 vccd1 _01600_
+ sky130_fd_sc_hd__mux2_1
X_07514_ top.cb_syn.char_path_n\[76\] top.cb_syn.char_path_n\[75\] top.cb_syn.char_path_n\[74\]
+ top.cb_syn.char_path_n\[73\] net399 net350 vssd1 vssd1 vccd1 vccd1 _04105_ sky130_fd_sc_hd__mux4_1
XANTENNA__06538__B top.findLeastValue.val1\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07445_ top.dut.bits_in_buf_next\[1\] _04031_ _04037_ _04038_ _04000_ vssd1 vssd1
+ vccd1 vccd1 _04039_ sky130_fd_sc_hd__a221o_1
XFILLER_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05659__B2 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07376_ top.cw1\[1\] net167 _03553_ net503 vssd1 vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__a22o_1
X_09115_ _02451_ _02452_ net479 _02774_ vssd1 vssd1 vccd1 vccd1 _05133_ sky130_fd_sc_hd__a31o_1
X_06327_ top.hist_data_o\[22\] top.hist_data_o\[21\] _03188_ vssd1 vssd1 vccd1 vccd1
+ _03190_ sky130_fd_sc_hd__and3_1
X_06258_ top.TRN_char_index\[1\] _02565_ _03122_ net460 vssd1 vssd1 vccd1 vccd1 _03125_
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout216_X net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09046_ net1123 top.WB.CPU_DAT_O\[11\] net293 vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout797_A net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06189_ _02960_ _03058_ vssd1 vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__nor2_1
Xhold440 top.findLeastValue.wipe_the_char_2 vssd1 vssd1 vccd1 vccd1 net1393 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09584__B net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold451 top.hTree.tree_reg\[40\] vssd1 vssd1 vccd1 vccd1 net1404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 top.path\[34\] vssd1 vssd1 vccd1 vccd1 net1415 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout585_X net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold495 top.path\[38\] vssd1 vssd1 vccd1 vccd1 net1448 sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 top.path\[87\] vssd1 vssd1 vccd1 vccd1 net1437 sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 top.cb_syn.char_path\[107\] vssd1 vssd1 vccd1 vccd1 net1426 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05595__B1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09948_ net737 net577 vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__and2_1
X_09879_ net760 net600 vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__and2_1
XFILLER_73_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11841_ clknet_leaf_116_clk _02357_ _01196_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07639__A2 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11772_ clknet_leaf_104_clk _02305_ _01127_ vssd1 vssd1 vccd1 vccd1 top.compVal\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10723_ clknet_leaf_112_clk _01322_ _00142_ vssd1 vssd1 vccd1 vccd1 top.path\[99\]
+ sky130_fd_sc_hd__dfrtp_1
X_10654_ clknet_leaf_60_clk _01253_ _00073_ vssd1 vssd1 vccd1 vccd1 top.hist_addr\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10585_ net751 net591 vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__and2_1
XANTENNA__07498__S1 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload18 clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 clkload18/Y sky130_fd_sc_hd__bufinv_16
Xclkload29 clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 clkload29/Y sky130_fd_sc_hd__inv_6
XANTENNA__05822__B2 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11206_ clknet_leaf_5_clk _01754_ _00561_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[108\]
+ sky130_fd_sc_hd__dfrtp_2
X_11137_ clknet_leaf_12_clk _01685_ _00492_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05586__B1 _02676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11068_ clknet_leaf_16_clk _01616_ _00423_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[98\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07327__A1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10019_ net845 net685 vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_19_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05560_ net457 top.hTree.node_reg\[52\] net361 net420 top.hTree.node_reg\[20\] vssd1
+ vssd1 vccd1 vccd1 _02655_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_47_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05491_ top.cb_syn.char_path\[31\] net560 net315 top.cb_syn.char_path\[127\] vssd1
+ vssd1 vccd1 vccd1 _02597_ sky130_fd_sc_hd__a22o_1
XANTENNA__06838__B1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05510__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07230_ net271 _03880_ _03881_ net276 net1674 vssd1 vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_119_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07161_ _03688_ _03691_ _03703_ _03708_ _03687_ vssd1 vssd1 vccd1 vccd1 _03819_ sky130_fd_sc_hd__o221a_1
X_06112_ top.cb_syn.char_index\[6\] _02961_ vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__xor2_1
XANTENNA__07489__S1 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07092_ top.findLeastValue.val1\[1\] top.findLeastValue.val2\[1\] vssd1 vssd1 vccd1
+ vccd1 _03750_ sky130_fd_sc_hd__xor2_1
X_06043_ _02931_ _02933_ vssd1 vssd1 vccd1 vccd1 _02934_ sky130_fd_sc_hd__nor2_1
XFILLER_99_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xfanout205 net211 vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09802_ net782 net622 vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__and2_1
XANTENNA__05437__B net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout227 net228 vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__clkbuf_4
Xfanout216 net217 vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__buf_2
Xfanout238 net239 vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__buf_2
X_07994_ _02499_ top.cb_syn.zeroes\[7\] top.cb_syn.zeroes\[6\] _02500_ vssd1 vssd1
+ vccd1 vccd1 _04497_ sky130_fd_sc_hd__o22a_1
XFILLER_101_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xfanout249 _04199_ vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__clkbuf_4
XANTENNA__05577__B1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09733_ net770 net610 vssd1 vssd1 vccd1 vccd1 _00347_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout280_A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06945_ top.findLeastValue.val2\[11\] net147 net121 _03614_ vssd1 vssd1 vccd1 vccd1
+ _01953_ sky130_fd_sc_hd__o22a_1
X_09664_ net784 net624 vssd1 vssd1 vccd1 vccd1 _00278_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout378_A net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06876_ top.compVal\[45\] top.findLeastValue.val1\[45\] net165 vssd1 vssd1 vccd1
+ vccd1 _03580_ sky130_fd_sc_hd__mux2_1
X_08615_ top.cb_syn.num_lefts\[6\] _04832_ vssd1 vssd1 vccd1 vccd1 _04834_ sky130_fd_sc_hd__nand2_1
X_09595_ net851 net691 vssd1 vssd1 vccd1 vccd1 _00209_ sky130_fd_sc_hd__and2_1
X_05827_ top.sram_interface.write_counter_FLV\[0\] net290 vssd1 vssd1 vccd1 vccd1
+ _02840_ sky130_fd_sc_hd__nand2_1
XANTENNA__05453__A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout545_A net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout166_X net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08546_ net1092 top.cb_syn.char_path_n\[30\] net232 vssd1 vssd1 vccd1 vccd1 _01548_
+ sky130_fd_sc_hd__mux2_1
X_05758_ top.compVal\[36\] net172 net158 top.WB.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1
+ _02321_ sky130_fd_sc_hd__a22o_1
XFILLER_23_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_08477_ net1233 top.cb_syn.char_path_n\[99\] net227 vssd1 vssd1 vccd1 vccd1 _01617_
+ sky130_fd_sc_hd__mux2_1
X_05689_ net26 net415 net308 top.WB.CPU_DAT_O\[31\] vssd1 vssd1 vccd1 vccd1 _02369_
+ sky130_fd_sc_hd__o22a_1
X_07428_ top.dut.bits_in_buf_next\[1\] _04014_ _04024_ _04001_ vssd1 vssd1 vccd1 vccd1
+ _04025_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout500_X net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07359_ _03753_ net270 _03972_ net275 top.findLeastValue.sum\[1\] vssd1 vssd1 vccd1
+ vccd1 _01897_ sky130_fd_sc_hd__a32o_1
XFILLER_108_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10370_ net853 net693 vssd1 vssd1 vccd1 vccd1 _00984_ sky130_fd_sc_hd__and2_1
XFILLER_109_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09029_ net1226 top.WB.CPU_DAT_O\[28\] net292 vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__mux2_1
Xhold270 top.path\[74\] vssd1 vssd1 vccd1 vccd1 net1223 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold292 top.hTree.nulls\[60\] vssd1 vssd1 vccd1 vccd1 net1245 sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 top.path\[49\] vssd1 vssd1 vccd1 vccd1 net1234 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05568__B1 _02661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout750 net757 vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__clkbuf_2
Xfanout783 net786 vssd1 vssd1 vccd1 vccd1 net783 sky130_fd_sc_hd__buf_1
Xfanout772 net807 vssd1 vssd1 vccd1 vccd1 net772 sky130_fd_sc_hd__clkbuf_2
Xfanout794 net796 vssd1 vssd1 vccd1 vccd1 net794 sky130_fd_sc_hd__clkbuf_2
Xfanout761 net762 vssd1 vssd1 vccd1 vccd1 net761 sky130_fd_sc_hd__buf_1
XANTENNA__06780__A2 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ clknet_leaf_100_clk _02340_ _01179_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11755_ clknet_leaf_99_clk _02288_ _01110_ vssd1 vssd1 vccd1 vccd1 top.compVal\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10706_ clknet_leaf_4_clk _01305_ _00125_ vssd1 vssd1 vccd1 vccd1 top.path\[82\]
+ sky130_fd_sc_hd__dfrtp_1
X_11686_ clknet_leaf_61_clk _02219_ _01041_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload118 clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 clkload118/Y sky130_fd_sc_hd__inv_6
Xclkload107 clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 clkload107/Y sky130_fd_sc_hd__bufinv_16
X_10637_ clknet_leaf_49_clk _00046_ _00056_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.word_cnt\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_116_Right_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10568_ net808 net648 vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__and2_1
X_10499_ net752 net592 vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_114_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05559__B1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput5 DAT_I[12] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
X_06730_ _03510_ _03514_ _03517_ vssd1 vssd1 vccd1 vccd1 _03518_ sky130_fd_sc_hd__or3_1
XFILLER_37_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10887__Q top.translation.index\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06661_ _02408_ top.findLeastValue.val2\[43\] _02483_ top.compVal\[42\] vssd1 vssd1
+ vccd1 vccd1 _03449_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_37_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06088__B top.cb_syn.char_index\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08400_ _04756_ _04757_ _04758_ net505 net438 vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__o221a_1
XANTENNA__07899__S net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05612_ top.cb_syn.char_path\[75\] net551 net542 top.cb_syn.char_path\[43\] vssd1
+ vssd1 vccd1 vccd1 _02698_ sky130_fd_sc_hd__a22o_1
X_09380_ net405 _04271_ vssd1 vssd1 vccd1 vccd1 _05264_ sky130_fd_sc_hd__nand2_1
X_06592_ _03350_ _03351_ _03352_ _03348_ vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__o31ai_1
XFILLER_24_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05543_ top.histogram.sram_out\[23\] net365 _02639_ _02640_ vssd1 vssd1 vccd1 vccd1
+ _02641_ sky130_fd_sc_hd__a211o_1
X_08331_ top.cb_syn.char_path_n\[4\] net380 net339 top.cb_syn.char_path_n\[2\] net184
+ vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__a221o_1
X_05474_ net495 net467 vssd1 vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__nand2_1
X_08262_ top.cb_syn.char_path_n\[38\] net200 _04658_ vssd1 vssd1 vccd1 vccd1 _01684_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__05495__C1 _02600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07213_ _03850_ _03851_ _03868_ vssd1 vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__nand3_1
X_08193_ top.cb_syn.char_path_n\[73\] net379 net338 top.cb_syn.char_path_n\[71\] net183
+ vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__a221o_1
XANTENNA__08433__C1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07787__A1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09320__S1 top.translation.index\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07144_ _03800_ _03801_ vssd1 vssd1 vccd1 vccd1 _03802_ sky130_fd_sc_hd__and2_1
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07075_ top.findLeastValue.val1\[9\] top.findLeastValue.val2\[9\] vssd1 vssd1 vccd1
+ vccd1 _03733_ sky130_fd_sc_hd__nand2_1
XANTENNA__08984__A0 top.WB.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06026_ top.hist_data_o\[9\] top.WB.CPU_DAT_O\[9\] net355 vssd1 vssd1 vccd1 vccd1
+ _02184_ sky130_fd_sc_hd__mux2_1
XFILLER_101_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07977_ net534 _02526_ _04480_ vssd1 vssd1 vccd1 vccd1 _04481_ sky130_fd_sc_hd__a21o_1
XFILLER_87_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09716_ net765 net605 vssd1 vssd1 vccd1 vccd1 _00330_ sky130_fd_sc_hd__and2_1
X_06928_ top.compVal\[19\] top.findLeastValue.val1\[19\] net161 vssd1 vssd1 vccd1
+ vccd1 _03606_ sky130_fd_sc_hd__mux2_1
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09647_ net780 net620 vssd1 vssd1 vccd1 vccd1 _00261_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout450_X net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06859_ top.findLeastValue.histo_index\[7\] net497 net498 vssd1 vssd1 vccd1 vccd1
+ _03573_ sky130_fd_sc_hd__and3_1
XANTENNA__07711__A1 top.findLeastValue.least2\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09578_ net766 net606 vssd1 vssd1 vccd1 vccd1 _00192_ sky130_fd_sc_hd__and2_1
XFILLER_43_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07602__S _04144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08529_ net1286 top.cb_syn.char_path_n\[47\] net221 vssd1 vssd1 vccd1 vccd1 _01565_
+ sky130_fd_sc_hd__mux2_1
X_11540_ clknet_leaf_0_clk _02088_ _00895_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06726__B top.findLeastValue.val2\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11471_ clknet_leaf_96_clk _02019_ _00826_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[11\]
+ sky130_fd_sc_hd__dfstp_2
X_10422_ net873 net713 vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__and2_1
XFILLER_109_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10353_ net872 net712 vssd1 vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__and2_1
XANTENNA__08975__A0 top.WB.CPU_DAT_O\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10284_ net726 net566 vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__and2_1
XANTENNA__06888__S net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_05_885 vssd1 vssd1 vccd1 vccd1 team_05_885/HI gpio_oeb[1] sky130_fd_sc_hd__conb_1
XFILLER_116_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xteam_05_896 vssd1 vssd1 vccd1 vccd1 team_05_896/HI gpio_out[11] sky130_fd_sc_hd__conb_1
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout591 net594 vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__clkbuf_2
Xfanout580 net584 vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__clkbuf_2
XFILLER_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05713__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11807_ clknet_leaf_91_clk _02324_ _01162_ vssd1 vssd1 vccd1 vccd1 top.compVal\[39\]
+ sky130_fd_sc_hd__dfrtp_1
X_11738_ clknet_leaf_66_clk _02271_ _01093_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.zero_cnt\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08851__B top.TRN_sram_complete vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11669_ clknet_leaf_44_clk _02202_ _01024_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08415__C1 top.cb_syn.end_cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08966__A0 top.WB.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08880_ net294 _05053_ vssd1 vssd1 vccd1 vccd1 _05054_ sky130_fd_sc_hd__nor2_1
X_07900_ top.findLeastValue.sum\[8\] _04425_ net395 vssd1 vssd1 vccd1 vccd1 _04426_
+ sky130_fd_sc_hd__mux2_1
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05555__X _02651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07831_ net485 _04369_ vssd1 vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__or2_1
X_07762_ net430 _04314_ _04315_ net260 vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__o211a_1
XANTENNA__05952__A0 top.WB.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09501_ net750 net590 vssd1 vssd1 vccd1 vccd1 _00115_ sky130_fd_sc_hd__and2_1
X_07693_ net398 _04259_ vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__nand2_1
X_06713_ _03492_ _03497_ vssd1 vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__nand2_1
XFILLER_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09432_ net964 vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__clkbuf_1
XFILLER_92_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06644_ top.compVal\[19\] top.compVal\[18\] top.compVal\[17\] top.compVal\[16\] vssd1
+ vssd1 vccd1 vccd1 _03433_ sky130_fd_sc_hd__or4_1
XFILLER_24_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09363_ net1458 net242 net218 _04334_ vssd1 vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__a22o_1
X_06575_ _03361_ _03362_ _03363_ vssd1 vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__a21o_1
XFILLER_40_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05526_ net1325 net139 _02626_ net175 vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__a22o_1
X_08314_ top.cb_syn.char_path_n\[12\] net195 _04684_ vssd1 vssd1 vccd1 vccd1 _01658_
+ sky130_fd_sc_hd__o21a_1
X_09294_ _03988_ net298 vssd1 vssd1 vccd1 vccd1 top.dut.bit_buf_next\[10\] sky130_fd_sc_hd__and2_1
X_05457_ net464 _02563_ vssd1 vssd1 vccd1 vccd1 _02565_ sky130_fd_sc_hd__nand2_2
XANTENNA__09857__B net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08245_ top.cb_syn.char_path_n\[47\] net377 net336 top.cb_syn.char_path_n\[45\] net181
+ vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout410_A _02788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08406__C1 _02504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05388_ top.hTree.wait_cnt vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__inv_2
X_08176_ top.cb_syn.char_path_n\[81\] net202 _04615_ vssd1 vssd1 vccd1 vccd1 _01727_
+ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout129_X net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08957__A0 top.WB.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07127_ _03783_ _03784_ vssd1 vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_63_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout877_A net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07058_ top.findLeastValue.val1\[13\] top.findLeastValue.val2\[13\] vssd1 vssd1 vccd1
+ vccd1 _03716_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout498_X net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06009_ net1615 top.WB.CPU_DAT_O\[26\] net357 vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_7_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_78_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_121_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05943__A0 top.WB.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10971_ clknet_leaf_16_clk _01519_ _00326_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_54_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_16_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11523_ clknet_leaf_65_clk _02071_ _00878_ vssd1 vssd1 vccd1 vccd1 top.cw1\[6\] sky130_fd_sc_hd__dfrtp_1
X_11454_ clknet_leaf_71_clk _02002_ _00809_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least2\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_109_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08948__A0 top.WB.CPU_DAT_O\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10405_ net792 net632 vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__and2_1
XANTENNA__08412__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11385_ clknet_leaf_85_clk _01933_ _00740_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_111_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10336_ net801 net641 vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__and2_1
X_10267_ net853 net693 vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__and2_1
Xclkbuf_4_9_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_9_0_clk sky130_fd_sc_hd__clkbuf_8
X_10198_ net863 net703 vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__and2_1
XANTENNA__07923__B2 top.findLeastValue.sum\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05934__A0 top.WB.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_06360_ top.hist_data_o\[19\] _03187_ top.hist_data_o\[20\] vssd1 vssd1 vccd1 vccd1
+ _03212_ sky130_fd_sc_hd__a21oi_1
X_06291_ _02885_ _02910_ _02942_ vssd1 vssd1 vccd1 vccd1 _03156_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09677__B net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05311_ top.compVal\[31\] vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_32_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08030_ _04510_ _04520_ _04526_ _04509_ top.cb_syn.count\[1\] vssd1 vssd1 vccd1 vccd1
+ _01784_ sky130_fd_sc_hd__a32o_1
Xinput30 DAT_I[6] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_1
Xinput41 gpio_in[7] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08939__A0 top.WB.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08403__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09981_ net781 net621 vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__and2_1
XANTENNA__09693__A net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10632__A net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08932_ top.WB.CPU_DAT_O\[22\] net1528 net371 vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__mux2_1
XANTENNA__06965__A2 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout193_A net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10351__B net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06717__A2 top.findLeastValue.val2\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08863_ top.translation.index\[5\] _02789_ top.translation.index\[6\] vssd1 vssd1
+ vccd1 vccd1 _05044_ sky130_fd_sc_hd__o21a_1
XANTENNA__05445__B top.CB_read_complete vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07814_ top.findLeastValue.sum\[25\] top.hTree.tree_reg\[25\] net283 vssd1 vssd1
+ vccd1 vccd1 _04357_ sky130_fd_sc_hd__mux2_1
XANTENNA__05925__A0 top.WB.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08794_ top.path\[26\] top.path\[27\] net524 vssd1 vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout360_A _02761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07745_ top.hTree.tree_reg\[39\] top.findLeastValue.sum\[39\] net250 vssd1 vssd1
+ vccd1 vccd1 _04302_ sky130_fd_sc_hd__mux2_1
XFILLER_37_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout458_A net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07676_ _02474_ net397 _04245_ vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__o21a_1
X_09415_ _02808_ _04216_ vssd1 vssd1 vccd1 vccd1 _05287_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout625_A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06627_ _03394_ _03415_ _03392_ vssd1 vssd1 vccd1 vccd1 _03416_ sky130_fd_sc_hd__o21a_1
X_09346_ net1050 net239 net217 _04402_ vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__a22o_1
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06558_ _03339_ _03343_ _03342_ _03340_ vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__a211o_1
X_09277_ _05213_ _05227_ _05214_ vssd1 vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__a21o_1
X_05509_ top.cb_syn.char_path\[92\] net553 net544 top.cb_syn.char_path\[60\] vssd1
+ vssd1 vccd1 vccd1 _02612_ sky130_fd_sc_hd__a22o_1
XANTENNA__07525__S0 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06489_ _03287_ net1514 vssd1 vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__nor2_1
X_08228_ top.cb_syn.char_path_n\[55\] net205 _04641_ vssd1 vssd1 vccd1 vccd1 _01701_
+ sky130_fd_sc_hd__o21a_1
XFILLER_32_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08159_ top.cb_syn.char_path_n\[90\] net387 net346 top.cb_syn.char_path_n\[88\] net191
+ vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_95_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11170_ clknet_leaf_11_clk _01718_ _00525_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[72\]
+ sky130_fd_sc_hd__dfrtp_2
X_10121_ net840 net680 vssd1 vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__and2_1
XANTENNA__09355__B1 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10052_ net845 net685 vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__and2_1
XANTENNA__07905__A1 top.findLeastValue.sum\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input19_A DAT_I[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10954_ clknet_leaf_40_clk _01509_ _00309_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_found
+ sky130_fd_sc_hd__dfrtp_1
X_10885_ clknet_leaf_110_clk _01462_ _00240_ vssd1 vssd1 vccd1 vccd1 top.translation.index\[0\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__07516__S0 _04072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11506_ clknet_leaf_85_clk _02054_ _00861_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[46\]
+ sky130_fd_sc_hd__dfstp_1
X_11437_ clknet_leaf_90_clk _01985_ _00792_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[43\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__08397__A1 _02506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11368_ clknet_leaf_106_clk _01916_ _00723_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10319_ net763 net603 vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__and2_1
XFILLER_112_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__09346__B1 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11299_ clknet_leaf_82_clk net1353 _00654_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_112_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05860_ top.compVal\[7\] net171 net156 top.WB.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1
+ _02282_ sky130_fd_sc_hd__a22o_1
XFILLER_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05791_ net452 _02810_ vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__nor2_1
XFILLER_93_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07530_ _04097_ _04120_ _04065_ vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__mux2_1
XFILLER_35_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07461_ top.cb_syn.i\[2\] top.cb_syn.cb_length\[2\] vssd1 vssd1 vccd1 vccd1 _04052_
+ sky130_fd_sc_hd__and2b_1
XANTENNA__06221__A1_N top.findLeastValue.histo_index\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_22_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07392_ _03990_ _03993_ _03986_ vssd1 vssd1 vccd1 vccd1 _03994_ sky130_fd_sc_hd__mux2_1
X_09200_ net264 _05058_ _05059_ _02825_ vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_17_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06412_ net1483 net299 _03173_ _03244_ vssd1 vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__a22o_1
X_06343_ net1279 _03202_ net303 vssd1 vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__mux2_1
X_09131_ _02529_ _02773_ _02778_ net451 vssd1 vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__and4bb_1
XANTENNA__07507__S0 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09062_ net1530 _05090_ _05091_ top.TRN_char_index\[5\] vssd1 vssd1 vccd1 vccd1 _01253_
+ sky130_fd_sc_hd__a22o_1
X_06274_ _02911_ _03139_ vssd1 vssd1 vccd1 vccd1 _03140_ sky130_fd_sc_hd__nor2_1
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08013_ _02501_ _04515_ vssd1 vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__nor2_1
Xhold611 top.cb_syn.pulse_first vssd1 vssd1 vccd1 vccd1 net1564 sky130_fd_sc_hd__dlygate4sd3_1
Xhold600 _03296_ vssd1 vssd1 vccd1 vccd1 net1553 sky130_fd_sc_hd__dlygate4sd3_1
Xhold644 top.histogram.state\[1\] vssd1 vssd1 vccd1 vccd1 net1597 sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 top.hist_data_o\[21\] vssd1 vssd1 vccd1 vccd1 net1586 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08388__A1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold622 top.hTree.tree_reg\[28\] vssd1 vssd1 vccd1 vccd1 net1575 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08531__S net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold677 top.histogram.total\[16\] vssd1 vssd1 vccd1 vccd1 net1630 sky130_fd_sc_hd__dlygate4sd3_1
Xhold666 top.hist_data_o\[4\] vssd1 vssd1 vccd1 vccd1 net1619 sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 top.compVal\[31\] vssd1 vssd1 vccd1 vccd1 net1641 sky130_fd_sc_hd__dlygate4sd3_1
Xhold655 top.histogram.total\[2\] vssd1 vssd1 vccd1 vccd1 net1608 sky130_fd_sc_hd__dlygate4sd3_1
X_09964_ net778 net618 vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__and2_1
Xhold699 top.sram_interface.word_cnt\[6\] vssd1 vssd1 vccd1 vccd1 net1652 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07655__B net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08915_ _04179_ _04187_ vssd1 vssd1 vccd1 vccd1 _05081_ sky130_fd_sc_hd__nor2_1
X_09895_ net775 net615 vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout196_X net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08846_ _05026_ _05028_ vssd1 vssd1 vccd1 vccd1 _05029_ sky130_fd_sc_hd__nor2_1
XANTENNA__07899__A0 top.findLeastValue.sum\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07363__A2 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05989_ _02914_ _02919_ vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout742_A net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08777_ top.path\[122\] top.path\[123\] net525 vssd1 vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__mux2_1
XFILLER_38_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07728_ net440 net1522 net251 top.findLeastValue.sum\[43\] _04288_ vssd1 vssd1 vccd1
+ vccd1 _01848_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout530_X net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07659_ net489 _04230_ vssd1 vssd1 vccd1 vccd1 _04233_ sky130_fd_sc_hd__or2_1
XANTENNA__05677__A2 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10670_ clknet_leaf_119_clk _01269_ _00089_ vssd1 vssd1 vccd1 vccd1 top.path\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_09329_ net487 _02809_ net262 _00053_ vssd1 vssd1 vccd1 vccd1 _05260_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_97_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07823__B1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06626__B2 top.compVal\[33\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11222_ clknet_leaf_29_clk _01770_ _00577_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[124\]
+ sky130_fd_sc_hd__dfrtp_2
X_11153_ clknet_leaf_26_clk _01701_ _00508_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_88_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11084_ clknet_leaf_23_clk _01632_ _00439_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[114\]
+ sky130_fd_sc_hd__dfrtp_1
X_10104_ net816 net656 vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__and2_1
XFILLER_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10035_ net839 net679 vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__and2_1
XANTENNA__06896__S net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10937_ clknet_leaf_28_clk _01492_ _00292_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.cb_length\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08854__A2 top.header_synthesis.enable vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06865__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08918__A_N _05072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10868_ clknet_leaf_76_clk _01454_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_14_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10799_ clknet_leaf_53_clk _00001_ _00218_ vssd1 vssd1 vccd1 vccd1 top.WB.curr_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__06093__A2 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05840__A2 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07756__A net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout409 _02788_ vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__clkbuf_2
X_06961_ top.findLeastValue.val2\[3\] net149 net122 _03622_ vssd1 vssd1 vccd1 vccd1
+ _01945_ sky130_fd_sc_hd__o22a_1
XANTENNA__08790__A1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05912_ top.sram_interface.init_counter\[5\] top.sram_interface.init_counter\[4\]
+ top.sram_interface.init_counter\[3\] top.sram_interface.init_counter\[2\] vssd1
+ vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__or4_1
X_08700_ _02457_ net517 _02930_ vssd1 vssd1 vccd1 vccd1 _04893_ sky130_fd_sc_hd__or3b_1
X_09680_ net797 net637 vssd1 vssd1 vccd1 vccd1 _00294_ sky130_fd_sc_hd__and2_1
XFILLER_79_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08631_ _04827_ _04835_ _04843_ _04826_ top.cb_syn.num_lefts\[1\] vssd1 vssd1 vccd1
+ vccd1 _01500_ sky130_fd_sc_hd__a32o_1
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06892_ top.compVal\[37\] top.findLeastValue.val1\[37\] net165 vssd1 vssd1 vccd1
+ vccd1 _03588_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05843_ top.compVal\[24\] net169 net155 top.WB.CPU_DAT_O\[24\] vssd1 vssd1 vccd1
+ vccd1 _02299_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_68_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05774_ top.findLeastValue.least1\[6\] top.findLeastValue.least1\[5\] top.findLeastValue.least1\[4\]
+ top.findLeastValue.least1\[7\] vssd1 vssd1 vccd1 vccd1 _02794_ sky130_fd_sc_hd__or4b_1
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08562_ net1269 top.cb_syn.char_path_n\[14\] net220 vssd1 vssd1 vccd1 vccd1 _01532_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__11514__Q top.findLeastValue.least1\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08493_ net1196 top.cb_syn.char_path_n\[83\] net223 vssd1 vssd1 vccd1 vccd1 _01601_
+ sky130_fd_sc_hd__mux2_1
X_07513_ top.cb_syn.char_path_n\[72\] top.cb_syn.char_path_n\[71\] top.cb_syn.char_path_n\[70\]
+ top.cb_syn.char_path_n\[69\] net399 net350 vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__mux4_1
X_07444_ top.dut.bits_in_buf\[1\] top.dut.bits_in_buf_next\[0\] vssd1 vssd1 vccd1
+ vccd1 _04038_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout156_A net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08845__A2 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05659__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07375_ net1620 net134 _03547_ net127 _03981_ vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__a32o_1
XFILLER_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09114_ _05130_ _05131_ vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__or2_1
X_06326_ top.hist_data_o\[21\] _03188_ vssd1 vssd1 vccd1 vccd1 _03189_ sky130_fd_sc_hd__and2_1
XANTENNA__06084__A2 top.cb_syn.char_index\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06257_ top.TRN_char_index\[1\] top.TRN_char_index\[0\] vssd1 vssd1 vccd1 vccd1 _03124_
+ sky130_fd_sc_hd__nand2b_1
X_09045_ net1096 top.WB.CPU_DAT_O\[12\] net293 vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold430 net46 vssd1 vssd1 vccd1 vccd1 net1383 sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 top.dut.out\[5\] vssd1 vssd1 vccd1 vccd1 net1394 sky130_fd_sc_hd__dlygate4sd3_1
X_06188_ top.cb_syn.char_index\[4\] _02958_ vssd1 vssd1 vccd1 vccd1 _03058_ sky130_fd_sc_hd__nor2_1
Xhold452 _01845_ vssd1 vssd1 vccd1 vccd1 net1405 sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 top.path\[52\] vssd1 vssd1 vccd1 vccd1 net1416 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold496 top.cb_syn.char_path\[0\] vssd1 vssd1 vccd1 vccd1 net1449 sky130_fd_sc_hd__dlygate4sd3_1
Xhold474 top.hTree.tree_reg\[35\] vssd1 vssd1 vccd1 vccd1 net1427 sky130_fd_sc_hd__dlygate4sd3_1
Xhold485 top.hTree.tree_reg\[2\] vssd1 vssd1 vccd1 vccd1 net1438 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout480_X net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09947_ net737 net577 vssd1 vssd1 vccd1 vccd1 _00561_ sky130_fd_sc_hd__and2_1
XANTENNA__06792__B1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09878_ net760 net600 vssd1 vssd1 vccd1 vccd1 _00492_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout745_X net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08829_ top.path\[42\] top.path\[43\] net528 vssd1 vssd1 vccd1 vccd1 _05012_ sky130_fd_sc_hd__mux2_1
XFILLER_45_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11840_ clknet_leaf_117_clk _02356_ _01195_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08297__B1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11771_ clknet_leaf_102_clk _02304_ _01126_ vssd1 vssd1 vccd1 vccd1 top.compVal\[29\]
+ sky130_fd_sc_hd__dfrtp_2
X_10722_ clknet_leaf_112_clk _01321_ _00141_ vssd1 vssd1 vccd1 vccd1 top.path\[98\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10653_ clknet_leaf_60_clk _01252_ _00072_ vssd1 vssd1 vccd1 vccd1 top.hist_addr\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10584_ net747 net587 vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__and2_1
XANTENNA__06075__A2 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload19 clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 clkload19/Y sky130_fd_sc_hd__bufinv_16
X_11205_ clknet_leaf_6_clk _01753_ _00560_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[107\]
+ sky130_fd_sc_hd__dfrtp_2
X_11136_ clknet_leaf_12_clk _01684_ _00491_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[38\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_1_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__06783__B1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05586__B2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11067_ clknet_leaf_16_clk _01615_ _00422_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[97\]
+ sky130_fd_sc_hd__dfrtp_1
X_10018_ net822 net662 vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__and2_1
XFILLER_49_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_47_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11969_ net453 vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06299__C1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06302__A3 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05490_ top.cb_syn.char_path\[95\] net554 net545 top.cb_syn.char_path\[63\] vssd1
+ vssd1 vccd1 vccd1 _02596_ sky130_fd_sc_hd__a22o_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_63_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07160_ _03697_ _03700_ _03698_ _03695_ vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__a211o_1
X_06111_ _02582_ _02982_ vssd1 vssd1 vccd1 vccd1 _02983_ sky130_fd_sc_hd__nor2_1
X_07091_ top.findLeastValue.val1\[1\] top.findLeastValue.val2\[1\] vssd1 vssd1 vccd1
+ vccd1 _03749_ sky130_fd_sc_hd__and2_1
XFILLER_105_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06042_ net536 _02869_ net431 vssd1 vssd1 vccd1 vccd1 _02933_ sky130_fd_sc_hd__a21o_1
Xfanout206 net207 vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__buf_2
X_09801_ net782 net622 vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__and2_1
Xfanout228 _04805_ vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__clkbuf_2
Xfanout217 net219 vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__clkbuf_2
XFILLER_113_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07993_ _04492_ _04493_ _04495_ vssd1 vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__or3_1
XANTENNA__06774__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05437__C top.findLeastValue.histo_index\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09732_ net769 net609 vssd1 vssd1 vccd1 vccd1 _00346_ sky130_fd_sc_hd__and2_1
Xfanout239 _05261_ vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__buf_2
XANTENNA_clkload10_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06944_ top.compVal\[11\] top.findLeastValue.val1\[11\] net162 vssd1 vssd1 vccd1
+ vccd1 _03614_ sky130_fd_sc_hd__mux2_1
X_09663_ net784 net624 vssd1 vssd1 vccd1 vccd1 _00277_ sky130_fd_sc_hd__and2_1
XANTENNA__09206__A _02530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05734__A _02763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout273_A _03658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06875_ top.findLeastValue.val2\[46\] net150 net125 top.findLeastValue.val1\[46\]
+ vssd1 vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__o22a_1
X_08614_ _04832_ vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__inv_2
X_09594_ net850 net690 vssd1 vssd1 vccd1 vccd1 _00208_ sky130_fd_sc_hd__and2_1
X_05826_ net289 _02839_ _02838_ net1527 vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__05453__B net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08545_ net1070 top.cb_syn.char_path_n\[31\] net234 vssd1 vssd1 vccd1 vccd1 _01549_
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout159_X net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05757_ top.compVal\[37\] net172 net158 top.WB.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1
+ _02322_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout440_A net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08476_ net1187 top.cb_syn.char_path_n\[100\] net227 vssd1 vssd1 vccd1 vccd1 _01618_
+ sky130_fd_sc_hd__mux2_1
X_05688_ net416 _02760_ vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__nand2_1
X_07427_ net354 _04010_ vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout705_A net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout326_X net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07358_ _03750_ _03751_ vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__nand2b_1
X_06309_ _02568_ net454 top.histogram.state\[3\] vssd1 vssd1 vccd1 vccd1 _03172_ sky130_fd_sc_hd__or3b_2
X_07289_ _03795_ _03805_ _03924_ vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__nand3_1
X_09028_ net1172 top.WB.CPU_DAT_O\[29\] net292 vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__mux2_1
Xhold260 net70 vssd1 vssd1 vccd1 vccd1 net1213 sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 top.cb_syn.char_path\[56\] vssd1 vssd1 vccd1 vccd1 net1224 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09400__C1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold293 top.cb_syn.char_path\[126\] vssd1 vssd1 vccd1 vccd1 net1246 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 net81 vssd1 vssd1 vccd1 vccd1 net1235 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05568__B2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout751 net754 vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__clkbuf_2
Xfanout740 net744 vssd1 vssd1 vccd1 vccd1 net740 sky130_fd_sc_hd__clkbuf_2
Xfanout784 net785 vssd1 vssd1 vccd1 vccd1 net784 sky130_fd_sc_hd__clkbuf_2
Xfanout773 net774 vssd1 vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__clkbuf_2
Xfanout762 net767 vssd1 vssd1 vccd1 vccd1 net762 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout795 net796 vssd1 vssd1 vccd1 vccd1 net795 sky130_fd_sc_hd__clkbuf_2
XFILLER_73_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11823_ clknet_leaf_100_clk _02339_ _01178_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_103_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05740__A1 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_119_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_119_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11754_ clknet_leaf_99_clk _02287_ _01109_ vssd1 vssd1 vccd1 vccd1 top.compVal\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08690__B1 _04875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11685_ clknet_leaf_62_clk _02218_ _01040_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_24_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ clknet_leaf_1_clk _01304_ _00124_ vssd1 vssd1 vccd1 vccd1 top.path\[81\]
+ sky130_fd_sc_hd__dfrtp_1
X_10636_ clknet_leaf_73_clk _00045_ _00055_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.word_cnt\[2\]
+ sky130_fd_sc_hd__dfrtp_4
Xclkload119 clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 clkload119/Y sky130_fd_sc_hd__bufinv_16
Xclkload108 clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 clkload108/Y sky130_fd_sc_hd__inv_8
XFILLER_6_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10567_ net752 net592 vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__and2_1
X_10498_ net809 net649 vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_114_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11119_ clknet_leaf_24_clk _01667_ _00474_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[21\]
+ sky130_fd_sc_hd__dfrtp_2
Xinput6 DAT_I[13] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
X_06660_ _02409_ top.findLeastValue.val2\[41\] _02484_ top.compVal\[40\] vssd1 vssd1
+ vccd1 vccd1 _03448_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_65_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05611_ net1351 net138 _02697_ net174 vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__a22o_1
XFILLER_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06591_ _02433_ top.findLeastValue.val1\[16\] _03350_ _03351_ vssd1 vssd1 vccd1 vccd1
+ _03380_ sky130_fd_sc_hd__a211oi_1
X_05542_ net456 top.hTree.node_reg\[55\] net362 net420 top.hTree.node_reg\[23\] vssd1
+ vssd1 vccd1 vccd1 _02640_ sky130_fd_sc_hd__a32o_1
X_08330_ top.cb_syn.char_path_n\[4\] net200 _04692_ vssd1 vssd1 vccd1 vccd1 _01650_
+ sky130_fd_sc_hd__o21a_1
XFILLER_51_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05473_ _02417_ _02418_ vssd1 vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__nor2_2
XFILLER_60_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08261_ top.cb_syn.char_path_n\[39\] net379 net337 top.cb_syn.char_path_n\[37\] net182
+ vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__a221o_1
XFILLER_20_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07212_ _03856_ _03867_ _03853_ vssd1 vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__a21o_1
XFILLER_9_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08192_ top.cb_syn.char_path_n\[73\] net200 _04623_ vssd1 vssd1 vccd1 vccd1 _01719_
+ sky130_fd_sc_hd__o21a_1
X_07143_ top.findLeastValue.val1\[23\] top.findLeastValue.val2\[23\] vssd1 vssd1 vccd1
+ vccd1 _03801_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_76_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07074_ top.findLeastValue.val1\[9\] top.findLeastValue.val2\[9\] vssd1 vssd1 vccd1
+ vccd1 _03732_ sky130_fd_sc_hd__and2_1
XFILLER_105_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_06025_ net1607 top.WB.CPU_DAT_O\[10\] net356 vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__mux2_1
XFILLER_101_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout488_A net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07976_ _02871_ _04479_ vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__nor2_1
XFILLER_101_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05464__A net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09715_ net765 net605 vssd1 vssd1 vccd1 vccd1 _00329_ sky130_fd_sc_hd__and2_1
X_06927_ top.findLeastValue.val2\[20\] net146 net120 _03605_ vssd1 vssd1 vccd1 vccd1
+ _01962_ sky130_fd_sc_hd__o22a_1
X_09646_ net780 net620 vssd1 vssd1 vccd1 vccd1 _00260_ sky130_fd_sc_hd__and2_1
XANTENNA__09161__A1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06858_ net497 net498 _03570_ vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_2_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05809_ top.sram_interface.counter_HTREE\[2\] _02828_ vssd1 vssd1 vccd1 vccd1 _02829_
+ sky130_fd_sc_hd__and2_1
X_09577_ net766 net606 vssd1 vssd1 vccd1 vccd1 _00191_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout822_A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06789_ top.findLeastValue.val1\[41\] net131 net115 top.compVal\[41\] vssd1 vssd1
+ vccd1 vccd1 _02049_ sky130_fd_sc_hd__o22a_1
X_08528_ net1276 top.cb_syn.char_path_n\[48\] net223 vssd1 vssd1 vccd1 vccd1 _01566_
+ sky130_fd_sc_hd__mux2_1
X_08459_ net1267 top.cb_syn.char_path_n\[117\] net229 vssd1 vssd1 vccd1 vccd1 _01635_
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__05486__B1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11470_ clknet_leaf_96_clk _02018_ _00825_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[10\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_7_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10421_ net873 net713 vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__and2_1
X_10352_ net871 net711 vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__and2_1
XFILLER_3_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08727__A1 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10283_ net726 net566 vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xteam_05_886 vssd1 vssd1 vccd1 vccd1 team_05_886/HI gpio_out[0] sky130_fd_sc_hd__conb_1
Xteam_05_897 vssd1 vssd1 vccd1 vccd1 team_05_897/HI gpio_out[12] sky130_fd_sc_hd__conb_1
Xfanout581 net584 vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__clkbuf_2
Xfanout570 net571 vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__buf_1
Xfanout592 net594 vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09152__B2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08360__C1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06757__X _03545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05713__B2 top.WB.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05821__B net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11806_ clknet_leaf_91_clk _02323_ _01161_ vssd1 vssd1 vccd1 vccd1 top.compVal\[38\]
+ sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11737_ clknet_leaf_50_clk _02270_ _01092_ vssd1 vssd1 vccd1 vccd1 top.CB_write_complete
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_60_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11668_ clknet_leaf_44_clk _02201_ _01023_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10619_ net804 net644 vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__and2_1
X_11599_ clknet_leaf_62_clk _02147_ _00954_ vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07830_ top.hTree.tree_reg\[22\] top.findLeastValue.sum\[22\] net248 vssd1 vssd1
+ vccd1 vccd1 _04370_ sky130_fd_sc_hd__mux2_1
X_07761_ net490 _04313_ vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_16_Left_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06712_ _03483_ _03485_ _03486_ _03499_ vssd1 vssd1 vccd1 vccd1 _03500_ sky130_fd_sc_hd__a31o_1
X_09500_ net756 net596 vssd1 vssd1 vccd1 vccd1 _00114_ sky130_fd_sc_hd__and2_1
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07692_ top.findLeastValue.least2\[3\] top.hTree.tree_reg\[49\] net281 vssd1 vssd1
+ vccd1 vccd1 _04259_ sky130_fd_sc_hd__mux2_1
X_09431_ net968 vssd1 vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06901__B1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05704__B2 top.WB.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06643_ top.compVal\[23\] top.compVal\[22\] top.compVal\[21\] top.compVal\[20\] vssd1
+ vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__or4_1
X_09362_ net1088 net242 net218 _04338_ vssd1 vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__a22o_1
X_06574_ _02443_ top.findLeastValue.val1\[6\] top.findLeastValue.val1\[5\] _02444_
+ vssd1 vssd1 vccd1 vccd1 _03363_ sky130_fd_sc_hd__a22o_1
XFILLER_24_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05525_ top.histogram.sram_out\[26\] net365 _02624_ _02625_ vssd1 vssd1 vccd1 vccd1
+ _02626_ sky130_fd_sc_hd__a211o_1
X_08313_ top.cb_syn.char_path_n\[13\] net373 net333 top.cb_syn.char_path_n\[11\] net178
+ vssd1 vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__a221o_1
X_09293_ _03989_ net298 vssd1 vssd1 vccd1 vccd1 top.dut.bit_buf_next\[9\] sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_25_Left_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05456_ net464 _02563_ vssd1 vssd1 vccd1 vccd1 _02564_ sky130_fd_sc_hd__and2_1
X_08244_ top.cb_syn.char_path_n\[47\] net198 _04649_ vssd1 vssd1 vccd1 vccd1 _01693_
+ sky130_fd_sc_hd__o21a_1
X_05387_ top.hTree.tree_reg\[54\] vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__inv_2
X_08175_ top.cb_syn.char_path_n\[82\] net382 net341 top.cb_syn.char_path_n\[80\] net186
+ vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__a221o_1
X_07126_ top.findLeastValue.val1\[17\] top.findLeastValue.val2\[17\] vssd1 vssd1 vccd1
+ vccd1 _03784_ sky130_fd_sc_hd__and2_1
X_07057_ _03711_ _03712_ _03713_ vssd1 vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout772_A net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout393_X net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06008_ net1604 top.WB.CPU_DAT_O\[27\] net357 vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_7_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_34_Left_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout560_X net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07959_ net1470 _04469_ _04461_ vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__mux2_1
XANTENNA__05481__X _02589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10970_ clknet_leaf_42_clk _01518_ _00325_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09629_ net755 net595 vssd1 vssd1 vccd1 vccd1 _00243_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_26_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Left_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08645__B1 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_50_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_clk sky130_fd_sc_hd__clkbuf_8
Xwire212 net213 vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__clkbuf_1
X_11522_ clknet_leaf_63_clk _02070_ _00877_ vssd1 vssd1 vccd1 vccd1 top.cw1\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_109_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11453_ clknet_leaf_70_clk _02001_ _00808_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least2\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10404_ net792 net632 vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__and2_1
X_11384_ clknet_leaf_85_clk _01932_ _00739_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06959__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10335_ net801 net641 vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__and2_1
X_10266_ net865 net705 vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_52_Left_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05631__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08176__A2 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09373__B2 _04294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10197_ net858 net698 vssd1 vssd1 vccd1 vccd1 _00811_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_109_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_61_Left_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05698__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_41_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_61_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05310_ net466 vssd1 vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__inv_2
X_06290_ _02574_ _02991_ _03153_ _03154_ vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_32_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput31 DAT_I[7] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
Xinput20 DAT_I[26] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
Xinput42 gpio_in[8] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__buf_1
XANTENNA__06382__B net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09980_ net781 net621 vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__and2_1
XANTENNA__09693__B net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07611__A1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_70_Left_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08931_ top.WB.CPU_DAT_O\[23\] net1308 net371 vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__mux2_1
XANTENNA__10632__B net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08862_ _02791_ _05042_ top.translation.resEn _02785_ vssd1 vssd1 vccd1 vccd1 _01469_
+ sky130_fd_sc_hd__a2bb2o_1
X_07813_ net442 net1459 net256 top.findLeastValue.sum\[26\] _04356_ vssd1 vssd1 vccd1
+ vccd1 _01831_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_4_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09116__A1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout186_A net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08793_ top.translation.index\[5\] _04970_ _04971_ _04975_ top.translation.index\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__o311a_1
XANTENNA__09116__B2 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08529__S net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07744_ top.findLeastValue.sum\[39\] top.hTree.tree_reg\[39\] net284 vssd1 vssd1
+ vccd1 vccd1 _04301_ sky130_fd_sc_hd__mux2_1
X_07675_ net397 _04244_ vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_84_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09414_ net978 net241 _05285_ _05286_ vssd1 vssd1 vccd1 vccd1 _01452_ sky130_fd_sc_hd__a22o_1
XFILLER_13_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_06626_ top.compVal\[34\] _02467_ _02468_ top.compVal\[33\] _03389_ vssd1 vssd1 vccd1
+ vccd1 _03415_ sky130_fd_sc_hd__o221a_1
XANTENNA__09419__A2 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08627__B1 _04826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_32_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout239_X net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06557_ _02430_ top.findLeastValue.val1\[19\] vssd1 vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__and2_1
X_09345_ net1008 net236 net215 _04406_ vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__a22o_1
X_05508_ net1319 net139 _02611_ net175 vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__a22o_1
X_09276_ top.cb_syn.zero_count\[6\] _05224_ vssd1 vssd1 vccd1 vccd1 _05227_ sky130_fd_sc_hd__nand2_1
XANTENNA__07525__S1 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06488_ top.histogram.total\[20\] _03286_ net1513 vssd1 vssd1 vccd1 vccd1 _03301_
+ sky130_fd_sc_hd__a21oi_1
X_05439_ top.findLeastValue.histo_index\[7\] net497 _02545_ _02546_ vssd1 vssd1 vccd1
+ vccd1 _02547_ sky130_fd_sc_hd__or4_1
X_08227_ top.cb_syn.char_path_n\[56\] net384 net343 top.cb_syn.char_path_n\[54\] net188
+ vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__a221o_1
XFILLER_119_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout406_X net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05861__B1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08158_ net1706 net210 _04606_ vssd1 vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__o21a_1
XFILLER_4_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08089_ top.cb_syn.char_path_n\[125\] net385 net345 top.cb_syn.char_path_n\[123\]
+ net189 vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__a221o_1
X_07109_ _03746_ _03759_ _03766_ _03745_ _03744_ vssd1 vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_95_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05613__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10120_ net821 net661 vssd1 vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__and2_1
XANTENNA__08158__A2 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10051_ net846 net686 vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_99_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_99_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__06169__B2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06169__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold732_A top.findLeastValue.sum\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10953_ clknet_leaf_41_clk _01508_ _00308_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.setup
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__07669__A1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10884_ clknet_leaf_49_clk _01461_ _00239_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.TRN_counter\[2\]
+ sky130_fd_sc_hd__dfrtp_2
Xclkbuf_leaf_23_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07516__S1 _04071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_11505_ clknet_leaf_89_clk _02053_ _00860_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[45\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__05852__B1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11436_ clknet_leaf_89_clk _01984_ _00791_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[42\]
+ sky130_fd_sc_hd__dfstp_1
X_11367_ clknet_leaf_101_clk _01915_ _00722_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10318_ net763 net603 vssd1 vssd1 vccd1 vccd1 _00932_ sky130_fd_sc_hd__and2_1
XANTENNA__05604__B1 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11298_ clknet_leaf_82_clk net1510 _00653_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[41\]
+ sky130_fd_sc_hd__dfrtp_1
X_10249_ net866 net706 vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__and2_1
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05907__B2 _02875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07372__A3 _03547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05790_ top.sram_interface.counter_HTREE\[3\] top.sram_interface.counter_HTREE\[1\]
+ top.sram_interface.counter_HTREE\[0\] top.sram_interface.counter_HTREE\[2\] vssd1
+ vssd1 vccd1 vccd1 _02810_ sky130_fd_sc_hd__or4b_1
XFILLER_93_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_62_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07460_ top.cb_syn.cb_length\[3\] top.cb_syn.i\[3\] vssd1 vssd1 vccd1 vccd1 _04051_
+ sky130_fd_sc_hd__and2b_1
XFILLER_22_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07391_ _03991_ _03992_ net404 vssd1 vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06411_ top.hist_data_o\[1\] top.hist_data_o\[0\] net300 vssd1 vssd1 vccd1 vccd1
+ _03244_ sky130_fd_sc_hd__o21a_1
XFILLER_34_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06883__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06342_ top.hist_data_o\[28\] _03198_ _03193_ vssd1 vssd1 vccd1 vccd1 _03202_ sky130_fd_sc_hd__o21ba_1
X_09130_ _02763_ _02773_ _02899_ _05114_ vssd1 vssd1 vccd1 vccd1 _05142_ sky130_fd_sc_hd__o22ai_1
XANTENNA__07507__S1 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_14_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_8
X_09061_ net1665 _05090_ _05091_ top.TRN_char_index\[6\] vssd1 vssd1 vccd1 vccd1 _01254_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_77_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06273_ top.sram_interface.init_counter\[2\] _02910_ vssd1 vssd1 vccd1 vccd1 _03139_
+ sky130_fd_sc_hd__nor2_1
X_08012_ top.cb_syn.count\[4\] _04513_ vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_120_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05843__B1 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold612 top.header_synthesis.count\[5\] vssd1 vssd1 vccd1 vccd1 net1565 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xhold601 top.hTree.tree_reg\[20\] vssd1 vssd1 vccd1 vccd1 net1554 sky130_fd_sc_hd__dlygate4sd3_1
Xhold645 _00033_ vssd1 vssd1 vccd1 vccd1 net1598 sky130_fd_sc_hd__dlygate4sd3_1
Xhold634 top.hist_data_o\[22\] vssd1 vssd1 vccd1 vccd1 net1587 sky130_fd_sc_hd__dlygate4sd3_1
Xhold623 _01833_ vssd1 vssd1 vccd1 vccd1 net1576 sky130_fd_sc_hd__dlygate4sd3_1
Xhold656 top.cb_syn.cb_length\[5\] vssd1 vssd1 vccd1 vccd1 net1609 sky130_fd_sc_hd__dlygate4sd3_1
X_09963_ net779 net619 vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__and2_1
Xhold667 top.cw2\[2\] vssd1 vssd1 vccd1 vccd1 net1620 sky130_fd_sc_hd__dlygate4sd3_1
Xhold678 top.findLeastValue.sum\[36\] vssd1 vssd1 vccd1 vccd1 net1631 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold689 top.cb_syn.zero_count\[4\] vssd1 vssd1 vccd1 vccd1 net1642 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08914_ top.cb_syn.max_index\[4\] _05080_ _05072_ vssd1 vssd1 vccd1 vccd1 _01390_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07655__C net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09894_ net771 net611 vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_15_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07348__B1 _03966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08845_ top.path\[44\] net410 _05027_ vssd1 vssd1 vccd1 vccd1 _05028_ sky130_fd_sc_hd__o21a_1
X_08776_ net434 _04957_ _04958_ vssd1 vssd1 vccd1 vccd1 _04959_ sky130_fd_sc_hd__o21a_1
X_05988_ top.sram_interface.init_counter\[6\] _02907_ vssd1 vssd1 vccd1 vccd1 _02919_
+ sky130_fd_sc_hd__nor2_1
X_07727_ net425 _04286_ _04287_ net259 vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout356_X net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07658_ net489 _04231_ vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__nand2_1
XFILLER_53_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07589_ top.cb_syn.max_index\[3\] _04136_ _04172_ _04175_ vssd1 vssd1 vccd1 vccd1
+ _04176_ sky130_fd_sc_hd__o22a_1
XFILLER_80_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_8_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_8_0_clk sky130_fd_sc_hd__clkbuf_8
X_06609_ _02408_ top.findLeastValue.val1\[43\] vssd1 vssd1 vccd1 vccd1 _03398_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout523_X net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09328_ net847 net687 vssd1 vssd1 vccd1 vccd1 _00053_ sky130_fd_sc_hd__and2_1
XFILLER_40_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09259_ top.cb_syn.zero_count\[0\] top.cb_syn.zero_count\[1\] vssd1 vssd1 vccd1 vccd1
+ _05215_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_97_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07823__A1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_111_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_5_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09025__A0 top.WB.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_107_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_11221_ clknet_leaf_29_clk _01769_ _00576_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[123\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08379__A2 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11152_ clknet_leaf_22_clk _01700_ _00507_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[54\]
+ sky130_fd_sc_hd__dfrtp_1
X_10103_ net812 net652 vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__and2_1
XFILLER_76_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11083_ clknet_leaf_7_clk _01631_ _00438_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[113\]
+ sky130_fd_sc_hd__dfrtp_1
X_10034_ net837 net677 vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__and2_1
XANTENNA_input31_A DAT_I[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08839__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10936_ clknet_leaf_41_clk _01491_ _00291_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.wait_cycle
+ sky130_fd_sc_hd__dfstp_2
X_10867_ clknet_leaf_76_clk _01453_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_14_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10798_ clknet_leaf_39_clk _00000_ _00217_ vssd1 vssd1 vccd1 vccd1 top.WB.curr_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__09016__A0 top.WB.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11419_ clknet_leaf_104_clk _01967_ _00774_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[25\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_117_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09319__A1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06960_ top.compVal\[3\] top.findLeastValue.val1\[3\] net164 vssd1 vssd1 vccd1 vccd1
+ _03622_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_3_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_8
X_05911_ top.sram_interface.CB_write_counter\[0\] _02880_ _02881_ vssd1 vssd1 vccd1
+ vccd1 _02267_ sky130_fd_sc_hd__o21a_1
X_06891_ top.findLeastValue.val2\[38\] net150 net123 _03587_ vssd1 vssd1 vccd1 vccd1
+ _01980_ sky130_fd_sc_hd__o22a_1
X_08630_ top.cb_syn.num_lefts\[1\] top.cb_syn.num_lefts\[0\] vssd1 vssd1 vccd1 vccd1
+ _04843_ sky130_fd_sc_hd__or2_1
XANTENNA__06002__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05842_ top.compVal\[25\] net169 net155 top.WB.CPU_DAT_O\[25\] vssd1 vssd1 vccd1
+ vccd1 _02300_ sky130_fd_sc_hd__a22o_1
XFILLER_82_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05773_ top.findLeastValue.least1\[3\] top.findLeastValue.least1\[2\] top.findLeastValue.least1\[1\]
+ top.findLeastValue.least1\[0\] vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__or4_1
X_08561_ net1205 top.cb_syn.char_path_n\[15\] net221 vssd1 vssd1 vccd1 vccd1 _01533_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08492_ net1192 top.cb_syn.char_path_n\[84\] net233 vssd1 vssd1 vccd1 vccd1 _01602_
+ sky130_fd_sc_hd__mux2_1
X_07512_ top.cb_syn.char_path_n\[68\] top.cb_syn.char_path_n\[67\] top.cb_syn.char_path_n\[66\]
+ top.cb_syn.char_path_n\[65\] net399 net351 vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__mux4_1
X_07443_ top.dut.bit_buf\[1\] net39 net722 vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__mux2_1
XANTENNA__05513__C1 _02615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07711__S net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout149_A net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07374_ top.findLeastValue.histo_index\[2\] _03553_ _03980_ vssd1 vssd1 vccd1 vccd1
+ _03981_ sky130_fd_sc_hd__a21o_1
X_09113_ net455 net462 _05112_ vssd1 vssd1 vccd1 vccd1 _05131_ sky130_fd_sc_hd__a21o_1
X_06325_ top.hist_data_o\[20\] top.hist_data_o\[19\] _03187_ vssd1 vssd1 vccd1 vccd1
+ _03188_ sky130_fd_sc_hd__and3_1
X_06256_ top.TRN_char_index\[0\] top.TRN_char_index\[1\] vssd1 vssd1 vccd1 vccd1 _03123_
+ sky130_fd_sc_hd__nand2b_1
XANTENNA__06851__A net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08542__S net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09044_ net1068 top.WB.CPU_DAT_O\[13\] net292 vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__mux2_1
XANTENNA__09007__A0 top.WB.CPU_DAT_O\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold420 top.cb_syn.char_path\[55\] vssd1 vssd1 vccd1 vccd1 net1373 sky130_fd_sc_hd__dlygate4sd3_1
Xhold453 net89 vssd1 vssd1 vccd1 vccd1 net1406 sky130_fd_sc_hd__dlygate4sd3_1
X_06187_ _02560_ _02976_ _03054_ _03056_ _03053_ vssd1 vssd1 vccd1 vccd1 _03057_ sky130_fd_sc_hd__o311a_1
Xhold431 net75 vssd1 vssd1 vccd1 vccd1 net1384 sky130_fd_sc_hd__dlygate4sd3_1
Xhold442 net101 vssd1 vssd1 vccd1 vccd1 net1395 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_104_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_92_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout685_A net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold486 top.hTree.nulls\[63\] vssd1 vssd1 vccd1 vccd1 net1439 sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 top.cb_syn.char_path\[52\] vssd1 vssd1 vccd1 vccd1 net1417 sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 _01840_ vssd1 vssd1 vccd1 vccd1 net1428 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_8_Left_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold497 top.hTree.tree_reg\[17\] vssd1 vssd1 vccd1 vccd1 net1450 sky130_fd_sc_hd__dlygate4sd3_1
X_09946_ net737 net577 vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__and2_1
XANTENNA__05473__Y _02581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09877_ net760 net600 vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08828_ top.path\[46\] top.path\[47\] net525 vssd1 vssd1 vccd1 vccd1 _05011_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout640_X net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08759_ top.path\[96\] top.path\[97\] top.path\[98\] top.path\[99\] net527 top.translation.index\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04942_ sky130_fd_sc_hd__mux4_1
X_11770_ clknet_leaf_97_clk _02303_ _01125_ vssd1 vssd1 vccd1 vccd1 top.compVal\[28\]
+ sky130_fd_sc_hd__dfrtp_2
X_10721_ clknet_leaf_112_clk _01320_ _00140_ vssd1 vssd1 vccd1 vccd1 top.path\[97\]
+ sky130_fd_sc_hd__dfrtp_1
X_10652_ clknet_leaf_60_clk _01251_ _00071_ vssd1 vssd1 vccd1 vccd1 top.hist_addr\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10583_ net746 net586 vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__and2_1
XANTENNA__08452__S net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06761__A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11204_ clknet_leaf_4_clk _01752_ _00559_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[106\]
+ sky130_fd_sc_hd__dfrtp_2
X_11135_ clknet_leaf_13_clk _01683_ _00490_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[37\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_input34_X net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11066_ clknet_leaf_42_clk _01614_ _00421_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[96\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05586__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_695 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10017_ net819 net659 vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__and2_1
XFILLER_91_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11968_ net453 vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__clkbuf_1
X_10919_ clknet_leaf_28_clk _01474_ _00274_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.i\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__05510__A2 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11350__Q top.findLeastValue.sum\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06110_ _02947_ _02981_ _02851_ vssd1 vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__o21a_1
X_07090_ top.findLeastValue.val1\[2\] top.findLeastValue.val2\[2\] vssd1 vssd1 vccd1
+ vccd1 _03748_ sky130_fd_sc_hd__and2_1
X_06041_ top.cb_syn.wait_cycle net431 vssd1 vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__nor2_1
XFILLER_99_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07992_ _04488_ _04489_ _04494_ _04490_ vssd1 vssd1 vccd1 vccd1 _04495_ sky130_fd_sc_hd__or4b_1
XANTENNA__06223__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout207 net211 vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__buf_2
X_09800_ net775 net615 vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__and2_1
Xfanout229 net235 vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__clkbuf_4
Xfanout218 net219 vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__buf_2
XFILLER_99_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06774__B2 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06774__A1 top.findLeastValue.least1\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09731_ net769 net609 vssd1 vssd1 vccd1 vccd1 _00345_ sky130_fd_sc_hd__and2_1
X_06943_ top.findLeastValue.val2\[12\] net147 net120 _03613_ vssd1 vssd1 vccd1 vccd1
+ _01954_ sky130_fd_sc_hd__o22a_1
X_09662_ net782 net622 vssd1 vssd1 vccd1 vccd1 _00276_ sky130_fd_sc_hd__and2_1
X_06874_ _03567_ _03576_ _02482_ vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__mux2_1
XFILLER_67_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08613_ top.cb_syn.num_lefts\[5\] top.cb_syn.num_lefts\[4\] _04829_ vssd1 vssd1 vccd1
+ vccd1 _04832_ sky130_fd_sc_hd__and3_1
X_09593_ net853 net693 vssd1 vssd1 vccd1 vccd1 _00207_ sky130_fd_sc_hd__and2_1
X_05825_ top.sram_interface.write_counter_FLV\[2\] top.sram_interface.write_counter_FLV\[1\]
+ top.sram_interface.write_counter_FLV\[0\] _02536_ _02538_ vssd1 vssd1 vccd1 vccd1
+ _02839_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout266_A net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08544_ net1287 top.cb_syn.char_path_n\[32\] net233 vssd1 vssd1 vccd1 vccd1 _01550_
+ sky130_fd_sc_hd__mux2_1
X_05756_ top.compVal\[38\] net173 _02783_ top.WB.CPU_DAT_O\[6\] vssd1 vssd1 vccd1
+ vccd1 _02323_ sky130_fd_sc_hd__a22o_1
XFILLER_23_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05687_ net450 top.WB.prev_BUSY_O _02759_ vssd1 vssd1 vccd1 vccd1 _02761_ sky130_fd_sc_hd__and3_1
X_08475_ net1262 top.cb_syn.char_path_n\[101\] net228 vssd1 vssd1 vccd1 vccd1 _01619_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout433_A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07426_ net1394 net297 _03999_ _04021_ _04023_ vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__a221o_1
XANTENNA__05501__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout221_X net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07357_ top.findLeastValue.sum\[2\] net275 net270 _03971_ vssd1 vssd1 vccd1 vccd1
+ _01898_ sky130_fd_sc_hd__a22o_1
XFILLER_108_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06308_ net450 top.histogram.state\[3\] net366 vssd1 vssd1 vccd1 vccd1 _03171_ sky130_fd_sc_hd__and3_1
XFILLER_108_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09027_ net1065 top.WB.CPU_DAT_O\[30\] net291 vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__mux2_1
X_07288_ _03810_ _03923_ vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__or2_1
X_06239_ top.cb_syn.curr_index\[4\] _02558_ _03105_ net460 _03104_ vssd1 vssd1 vccd1
+ vccd1 _03107_ sky130_fd_sc_hd__a221o_1
XANTENNA__09400__B1 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold261 top.histogram.sram_out\[21\] vssd1 vssd1 vccd1 vccd1 net1214 sky130_fd_sc_hd__dlygate4sd3_1
Xhold250 top.cb_syn.char_path\[110\] vssd1 vssd1 vccd1 vccd1 net1203 sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 top.cb_syn.char_path\[88\] vssd1 vssd1 vccd1 vccd1 net1236 sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 top.cb_syn.char_path\[35\] vssd1 vssd1 vccd1 vccd1 net1225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 top.cb_syn.char_path\[106\] vssd1 vssd1 vccd1 vccd1 net1247 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06765__A1 top.findLeastValue.histo_index\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05568__A2 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout741 net744 vssd1 vssd1 vccd1 vccd1 net741 sky130_fd_sc_hd__clkbuf_2
Xfanout730 net731 vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__buf_1
Xfanout785 net786 vssd1 vssd1 vccd1 vccd1 net785 sky130_fd_sc_hd__clkbuf_2
X_09929_ net776 net616 vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__and2_1
Xfanout774 net776 vssd1 vssd1 vccd1 vccd1 net774 sky130_fd_sc_hd__clkbuf_2
Xfanout763 net767 vssd1 vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__clkbuf_2
Xfanout752 net754 vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__clkbuf_2
Xfanout796 net806 vssd1 vssd1 vccd1 vccd1 net796 sky130_fd_sc_hd__buf_1
XFILLER_46_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11822_ clknet_leaf_99_clk _02338_ _01177_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_103_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05740__A2 _02763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11753_ clknet_leaf_96_clk _02286_ _01108_ vssd1 vssd1 vccd1 vccd1 top.compVal\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11684_ clknet_leaf_63_clk _02217_ _01039_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_24_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ clknet_leaf_1_clk _01303_ _00123_ vssd1 vssd1 vccd1 vccd1 top.path\[80\]
+ sky130_fd_sc_hd__dfrtp_1
X_10635_ clknet_leaf_73_clk _00044_ _00054_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.word_cnt\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload109 clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 clkload109/Y sky130_fd_sc_hd__inv_12
X_10566_ net810 net650 vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__and2_1
X_10497_ net814 net654 vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_114_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08910__S _05072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11118_ clknet_leaf_24_clk _01666_ _00473_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06174__A1_N net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11049_ clknet_leaf_8_clk _01597_ _00404_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[79\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput7 DAT_I[14] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_91_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05610_ top.histogram.sram_out\[12\] net363 net419 top.hTree.node_reg\[12\] _02696_
+ vssd1 vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__a221o_2
X_06590_ _03370_ _03371_ _03373_ _03374_ _03378_ vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__o221ai_1
X_05541_ _02637_ _02638_ net476 vssd1 vssd1 vccd1 vccd1 _02639_ sky130_fd_sc_hd__o21a_1
X_05472_ _02575_ _02578_ _02579_ vssd1 vssd1 vccd1 vccd1 _02580_ sky130_fd_sc_hd__or3_1
X_08260_ top.cb_syn.char_path_n\[39\] net199 _04657_ vssd1 vssd1 vccd1 vccd1 _01685_
+ sky130_fd_sc_hd__o21a_1
X_08191_ top.cb_syn.char_path_n\[74\] net379 net338 top.cb_syn.char_path_n\[72\] net183
+ vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__a221o_1
X_07211_ _03837_ _03838_ _03846_ vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_89_Left_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_07142_ top.findLeastValue.val1\[23\] top.findLeastValue.val2\[23\] vssd1 vssd1 vccd1
+ vccd1 _03800_ sky130_fd_sc_hd__or2_1
XANTENNA__08433__A1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07073_ _03729_ _03730_ vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__nor2_1
XANTENNA__05448__C _02555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06024_ net1481 top.WB.CPU_DAT_O\[11\] net356 vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__mux2_1
XFILLER_101_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07975_ _04478_ vssd1 vssd1 vccd1 vccd1 _04479_ sky130_fd_sc_hd__inv_2
XANTENNA__09217__A top.controller.fin_reg\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_98_Left_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09714_ net792 net632 vssd1 vssd1 vccd1 vccd1 _00328_ sky130_fd_sc_hd__and2_1
X_06926_ top.compVal\[20\] top.findLeastValue.val1\[20\] net161 vssd1 vssd1 vccd1
+ vccd1 _03605_ sky130_fd_sc_hd__mux2_1
X_09645_ net803 net643 vssd1 vssd1 vccd1 vccd1 _00259_ sky130_fd_sc_hd__and2_1
X_06857_ net498 _03570_ vssd1 vssd1 vccd1 vccd1 _03571_ sky130_fd_sc_hd__and2_1
X_05808_ top.sram_interface.counter_HTREE\[1\] top.sram_interface.counter_HTREE\[0\]
+ _02826_ vssd1 vssd1 vccd1 vccd1 _02828_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout269_X net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_fanout171_X net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09576_ net766 net606 vssd1 vssd1 vccd1 vccd1 _00190_ sky130_fd_sc_hd__and2_1
X_06788_ top.findLeastValue.val1\[42\] net131 net115 top.compVal\[42\] vssd1 vssd1
+ vccd1 vccd1 _02050_ sky130_fd_sc_hd__o22a_1
X_05739_ net453 net423 vssd1 vssd1 vccd1 vccd1 _02774_ sky130_fd_sc_hd__nor2_1
X_08527_ net1227 top.cb_syn.char_path_n\[49\] net223 vssd1 vssd1 vccd1 vccd1 _01567_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout436_X net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08458_ net1284 top.cb_syn.char_path_n\[118\] net229 vssd1 vssd1 vccd1 vccd1 _01636_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09887__A net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07409_ top.dut.out\[7\] _04008_ top.dut.out_valid_next vssd1 vssd1 vccd1 vccd1 _04009_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09102__D _02763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10420_ net873 net713 vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__and2_1
X_08389_ _04733_ _04747_ top.cb_syn.end_cnt\[5\] vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__or3b_1
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_10351_ net866 net706 vssd1 vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__and2_1
XANTENNA__07694__X _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10282_ net726 net566 vssd1 vssd1 vccd1 vccd1 _00896_ sky130_fd_sc_hd__and2_1
XANTENNA__08727__A2 _04188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07935__A0 top.findLeastValue.sum\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xteam_05_887 vssd1 vssd1 vccd1 vccd1 team_05_887/HI gpio_out[2] sky130_fd_sc_hd__conb_1
Xfanout560 top.sram_interface.word_cnt\[0\] vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__buf_2
Xfanout582 net584 vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__clkbuf_2
Xteam_05_898 vssd1 vssd1 vccd1 vccd1 team_05_898/HI gpio_out[13] sky130_fd_sc_hd__conb_1
Xfanout593 net594 vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__buf_1
Xfanout571 net574 vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__buf_1
XFILLER_86_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05713__A2 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11805_ clknet_leaf_93_clk _02322_ _01160_ vssd1 vssd1 vccd1 vccd1 top.compVal\[37\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_33_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11736_ clknet_leaf_50_clk _02269_ _01091_ vssd1 vssd1 vccd1 vccd1 top.CB_read_complete
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05477__A1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11667_ clknet_leaf_45_clk _02200_ _01022_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10618_ net804 net644 vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__and2_1
X_11598_ clknet_leaf_43_clk _02146_ _00953_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08415__A1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06652__C net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10549_ net829 net669 vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__and2_1
XFILLER_111_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_111_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_71_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07760_ top.findLeastValue.sum\[36\] _04313_ net398 vssd1 vssd1 vccd1 vccd1 _04314_
+ sky130_fd_sc_hd__mux2_1
X_06711_ _03490_ _03493_ _03496_ _03498_ vssd1 vssd1 vccd1 vccd1 _03499_ sky130_fd_sc_hd__or4_1
X_09430_ net989 vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__clkbuf_1
X_07691_ net263 _04257_ _04258_ net1018 net446 vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__a32o_1
XFILLER_37_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06642_ top.compVal\[31\] top.compVal\[30\] top.compVal\[29\] top.compVal\[28\] vssd1
+ vssd1 vccd1 vccd1 _03431_ sky130_fd_sc_hd__or4_1
XANTENNA__06396__A net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09361_ net1517 net242 net219 _04342_ vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__a22o_1
X_06573_ _02444_ top.findLeastValue.val1\[5\] top.findLeastValue.val1\[4\] _02445_
+ vssd1 vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__o22a_1
X_09292_ _03991_ net298 vssd1 vssd1 vccd1 vccd1 top.dut.bit_buf_next\[8\] sky130_fd_sc_hd__and2_1
X_05524_ net456 top.hTree.node_reg\[58\] _02583_ net420 top.hTree.node_reg\[26\] vssd1
+ vssd1 vccd1 vccd1 _02625_ sky130_fd_sc_hd__a32o_1
XANTENNA__08103__B1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08312_ top.cb_syn.char_path_n\[13\] net195 _04683_ vssd1 vssd1 vccd1 vccd1 _01659_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__09300__C1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08243_ top.cb_syn.char_path_n\[48\] net376 net336 top.cb_syn.char_path_n\[46\] net181
+ vssd1 vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__a221o_1
XANTENNA__09500__A net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05455_ net541 _02562_ vssd1 vssd1 vccd1 vccd1 _02563_ sky130_fd_sc_hd__or2_2
XANTENNA_fanout229_A net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout131_A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07862__C1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08406__B2 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05386_ top.cw2\[0\] vssd1 vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__inv_2
X_08174_ top.cb_syn.char_path_n\[82\] net202 _04614_ vssd1 vssd1 vccd1 vccd1 _01728_
+ sky130_fd_sc_hd__o21a_1
XFILLER_106_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07125_ top.findLeastValue.val1\[17\] top.findLeastValue.val2\[17\] vssd1 vssd1 vccd1
+ vccd1 _03783_ sky130_fd_sc_hd__nor2_1
X_07056_ _03712_ _03713_ vssd1 vssd1 vccd1 vccd1 _03714_ sky130_fd_sc_hd__nand2_1
XANTENNA__08550__S net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06007_ net1594 top.WB.CPU_DAT_O\[28\] net358 vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_7_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_07958_ top.findLeastValue.least1\[0\] top.findLeastValue.least2\[0\] _04462_ vssd1
+ vssd1 vccd1 vccd1 _04469_ sky130_fd_sc_hd__mux2_1
XANTENNA__08786__A net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout553_X net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06909_ top.findLeastValue.val2\[29\] net148 net121 _03596_ vssd1 vssd1 vccd1 vccd1
+ _01971_ sky130_fd_sc_hd__o22a_1
X_07889_ top.findLeastValue.sum\[10\] top.hTree.tree_reg\[10\] net278 vssd1 vssd1
+ vccd1 vccd1 _04417_ sky130_fd_sc_hd__mux2_1
X_09628_ net757 net597 vssd1 vssd1 vccd1 vccd1 _00242_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_26_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09559_ net843 net683 vssd1 vssd1 vccd1 vccd1 _00173_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_54_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10556__A net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire213 _02587_ vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__clkbuf_1
X_11521_ clknet_leaf_63_clk _02069_ _00876_ vssd1 vssd1 vccd1 vccd1 top.cw1\[4\] sky130_fd_sc_hd__dfrtp_1
X_11452_ clknet_leaf_70_clk _02000_ _00807_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least2\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10403_ net793 net633 vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__and2_1
X_11383_ clknet_leaf_85_clk _01931_ _00738_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[35\]
+ sky130_fd_sc_hd__dfrtp_1
X_10334_ net792 net632 vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_111_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10265_ net868 net708 vssd1 vssd1 vccd1 vccd1 _00879_ sky130_fd_sc_hd__and2_1
X_10196_ net858 net698 vssd1 vssd1 vccd1 vccd1 _00810_ sky130_fd_sc_hd__and2_1
Xfanout390 _04564_ vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__buf_2
XFILLER_19_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07804__S net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload7_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08884__A1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05832__B net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05698__B2 top.WB.CPU_DAT_O\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11719_ clknet_leaf_122_clk _02252_ _01074_ vssd1 vssd1 vccd1 vccd1 top.path\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xinput21 DAT_I[27] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
Xinput10 DAT_I[17] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
Xinput43 gpio_in[9] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__buf_1
Xinput32 DAT_I[8] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_1
XFILLER_107_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08930_ top.WB.CPU_DAT_O\[24\] net1314 net372 vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__mux2_1
X_08861_ _02519_ _02785_ vssd1 vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__nor2_1
XFILLER_111_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_97_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07812_ net428 _04354_ _04355_ net259 vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_4_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08792_ _04969_ _04972_ _04973_ _04974_ _02520_ vssd1 vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__a221o_1
XANTENNA__07714__S net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07743_ net443 net1404 net254 top.findLeastValue.sum\[40\] _04300_ vssd1 vssd1 vccd1
+ vccd1 _01845_ sky130_fd_sc_hd__a221o_1
X_07674_ top.findLeastValue.least2\[6\] top.hTree.tree_reg\[52\] net280 vssd1 vssd1
+ vccd1 vccd1 _04244_ sky130_fd_sc_hd__mux2_1
XANTENNA__08875__A1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09413_ top.hTree.nulls\[58\] net407 net244 vssd1 vssd1 vccd1 vccd1 _05286_ sky130_fd_sc_hd__o21a_1
XANTENNA__05689__B2 top.WB.CPU_DAT_O\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06625_ _03397_ _03398_ vssd1 vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__nand2b_1
XANTENNA__08545__S net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06556_ _02430_ top.findLeastValue.val1\[19\] top.findLeastValue.val1\[18\] _02431_
+ vssd1 vssd1 vccd1 vccd1 _03345_ sky130_fd_sc_hd__o22a_1
X_09344_ net991 net237 net214 _04410_ vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__a22o_1
X_09275_ _05213_ _05225_ _05226_ _05214_ net1603 vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_zero_count\[5\]
+ sky130_fd_sc_hd__a32o_1
X_05507_ top.histogram.sram_out\[29\] net365 _02609_ _02610_ vssd1 vssd1 vccd1 vccd1
+ _02611_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout513_A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06487_ _03288_ _03300_ vssd1 vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__nor2_1
X_08226_ top.cb_syn.char_path_n\[56\] net205 _04640_ vssd1 vssd1 vccd1 vccd1 _01702_
+ sky130_fd_sc_hd__o21a_1
X_05438_ net503 net504 vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__or2_1
XFILLER_20_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08157_ top.cb_syn.char_path_n\[91\] net387 net348 top.cb_syn.char_path_n\[89\] net193
+ vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__a221o_1
XANTENNA__05861__B2 top.WB.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05369_ top.findLeastValue.least2\[3\] vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__inv_2
XANTENNA__09052__A1 top.WB.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07108_ _03765_ vssd1 vssd1 vccd1 vccd1 _03766_ sky130_fd_sc_hd__inv_2
X_08088_ top.cb_syn.char_path_n\[125\] net206 _04571_ vssd1 vssd1 vccd1 vccd1 _01771_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_95_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06810__B1 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07039_ top.findLeastValue.val1\[29\] top.findLeastValue.val2\[29\] vssd1 vssd1 vccd1
+ vccd1 _03697_ sky130_fd_sc_hd__nand2_1
X_10050_ net846 net686 vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__and2_1
XFILLER_87_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07624__S net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10952_ clknet_leaf_42_clk _01507_ _00307_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.end_check
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_90_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold725_A top.findLeastValue.sum\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08315__B1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06877__B1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10883_ clknet_leaf_47_clk _01460_ _00238_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.TRN_counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08455__S net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06764__A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11504_ clknet_leaf_89_clk _02052_ _00859_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[44\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_59_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05852__B2 top.WB.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09043__A1 top.WB.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11435_ clknet_leaf_90_clk _01983_ _00790_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[41\]
+ sky130_fd_sc_hd__dfstp_1
X_11366_ clknet_leaf_106_clk _01914_ _00721_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_112_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11297_ clknet_leaf_85_clk net1405 _00652_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06801__B1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10317_ net764 net604 vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__and2_1
X_10248_ net860 net700 vssd1 vssd1 vccd1 vccd1 _00862_ sky130_fd_sc_hd__and2_1
XANTENNA__09346__A2 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07357__A1 top.findLeastValue.sum\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10179_ net838 net678 vssd1 vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__and2_1
X_06410_ top.histogram.sram_out\[2\] _03243_ net301 vssd1 vssd1 vccd1 vccd1 _02117_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__11353__Q top.findLeastValue.sum\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07390_ top.dut.bit_buf\[7\] top.dut.bit_buf\[0\] net721 vssd1 vssd1 vccd1 vccd1
+ _03992_ sky130_fd_sc_hd__mux2_1
XANTENNA__08365__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05540__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06341_ net1183 _03201_ net302 vssd1 vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__mux2_1
XANTENNA__07817__C1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09060_ top.histogram.eof_n _05089_ _05090_ vssd1 vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__o21ba_2
XANTENNA__06096__A1 top.cb_syn.char_index\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06272_ _03134_ _03136_ _03137_ net470 vssd1 vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__o31a_1
XFILLER_30_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08011_ _04513_ vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__inv_2
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold602 top.hTree.tree_reg\[27\] vssd1 vssd1 vccd1 vccd1 net1555 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09034__A1 top.WB.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05843__B2 top.WB.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold624 top.cw1\[6\] vssd1 vssd1 vccd1 vccd1 net1577 sky130_fd_sc_hd__dlygate4sd3_1
Xhold635 top.hTree.tree_reg\[22\] vssd1 vssd1 vccd1 vccd1 net1588 sky130_fd_sc_hd__dlygate4sd3_1
Xhold613 top.findLeastValue.sum\[16\] vssd1 vssd1 vccd1 vccd1 net1566 sky130_fd_sc_hd__dlygate4sd3_1
Xhold679 top.cb_syn.zero_count\[3\] vssd1 vssd1 vccd1 vccd1 net1632 sky130_fd_sc_hd__dlygate4sd3_1
Xhold646 top.header_synthesis.start vssd1 vssd1 vccd1 vccd1 net1599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 top.cw2\[6\] vssd1 vssd1 vccd1 vccd1 net1610 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09962_ net777 net617 vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__and2_1
Xhold668 top.histogram.total\[0\] vssd1 vssd1 vccd1 vccd1 net1621 sky130_fd_sc_hd__dlygate4sd3_1
X_08913_ _04168_ _04187_ _05079_ vssd1 vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__a21bo_1
X_09893_ net774 net614 vssd1 vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__and2_1
XFILLER_111_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08844_ top.path\[45\] net328 _05011_ net434 top.translation.index\[2\] vssd1 vssd1
+ vccd1 vccd1 _05027_ sky130_fd_sc_hd__o221a_1
X_05987_ _02908_ _02918_ vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__nor2_1
X_08775_ top.path\[112\] net410 net328 top.path\[113\] _02522_ vssd1 vssd1 vccd1 vccd1
+ _04958_ sky130_fd_sc_hd__o221a_1
XANTENNA__06020__A1 top.WB.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout463_A net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07726_ net482 _04285_ vssd1 vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__or2_1
XFILLER_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout349_X net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout630_A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07657_ top.findLeastValue.least1\[1\] net250 _04229_ vssd1 vssd1 vccd1 vccd1 _04231_
+ sky130_fd_sc_hd__a21oi_1
X_07588_ net537 _04171_ _04174_ net531 vssd1 vssd1 vccd1 vccd1 _04175_ sky130_fd_sc_hd__a22o_1
XANTENNA__05531__B1 _02629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06608_ _02461_ top.compVal\[42\] _02408_ top.findLeastValue.val1\[43\] vssd1 vssd1
+ vccd1 vccd1 _03397_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_40_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09327_ _02543_ _05200_ _04922_ vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_write_zeroes
+ sky130_fd_sc_hd__o21ai_1
X_06539_ _02419_ top.findLeastValue.val1\[31\] top.findLeastValue.val1\[30\] _02420_
+ vssd1 vssd1 vccd1 vccd1 _03328_ sky130_fd_sc_hd__o22a_1
XFILLER_40_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09258_ _05213_ _05214_ top.cb_syn.zero_count\[0\] vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_zero_count\[0\]
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05834__A1 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08209_ top.cb_syn.char_path_n\[65\] net388 net347 top.cb_syn.char_path_n\[63\] net191
+ vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__a221o_1
X_09189_ _03324_ _04188_ vssd1 vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__nand2_1
XANTENNA__05487__X _02595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_11220_ clknet_leaf_29_clk _01768_ _00575_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[122\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_5_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_11151_ clknet_leaf_22_clk _01699_ _00506_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[53\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__05598__B1 _02686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10102_ net827 net667 vssd1 vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__and2_1
X_11082_ clknet_leaf_7_clk _01630_ _00437_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[112\]
+ sky130_fd_sc_hd__dfrtp_1
X_10033_ net837 net677 vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__and2_1
XANTENNA__06011__A1 top.WB.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input24_A DAT_I[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10935_ clknet_leaf_36_clk _01490_ _00290_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.state8
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05522__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10866_ clknet_leaf_46_clk _01452_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_14_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10797_ clknet_leaf_51_clk _00037_ _00216_ vssd1 vssd1 vccd1 vccd1 top.histogram.wr_r_en\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06781__X _03553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11418_ clknet_leaf_104_clk _01966_ _00773_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[24\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_117_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05589__B1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11349_ clknet_leaf_93_clk _01897_ _00704_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_67_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11348__Q top.findLeastValue.sum\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05910_ _02562_ _02880_ _02882_ _02881_ top.sram_interface.CB_write_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__a32o_1
X_06890_ top.compVal\[38\] top.findLeastValue.val1\[38\] net165 vssd1 vssd1 vccd1
+ vccd1 _03587_ sky130_fd_sc_hd__mux2_1
XFILLER_94_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06002__A1 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05841_ top.compVal\[26\] net169 net155 top.WB.CPU_DAT_O\[26\] vssd1 vssd1 vccd1
+ vccd1 _02301_ sky130_fd_sc_hd__a22o_1
X_08560_ net1159 top.cb_syn.char_path_n\[16\] net222 vssd1 vssd1 vccd1 vccd1 _01534_
+ sky130_fd_sc_hd__mux2_1
X_05772_ _02792_ _02787_ net1633 vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__mux2_1
X_07511_ _04098_ _04099_ _04100_ _04101_ _04072_ _04071_ vssd1 vssd1 vccd1 vccd1 _04102_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_81_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08491_ net1294 top.cb_syn.char_path_n\[85\] net233 vssd1 vssd1 vccd1 vccd1 _01603_
+ sky130_fd_sc_hd__mux2_1
X_07442_ _04001_ _04017_ _04036_ _03999_ _04033_ vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__a221o_1
XANTENNA__05513__B1 _02614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07373_ top.cw1\[2\] net167 vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__and2_1
X_09112_ net451 net423 vssd1 vssd1 vccd1 vccd1 _05130_ sky130_fd_sc_hd__nor2_1
X_06324_ top.hist_data_o\[18\] top.hist_data_o\[17\] _03185_ vssd1 vssd1 vccd1 vccd1
+ _03187_ sky130_fd_sc_hd__and3_1
XFILLER_30_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06255_ top.cb_syn.max_index\[3\] _03025_ _03027_ top.hTree.nullSumIndex\[2\] vssd1
+ vssd1 vccd1 vccd1 _03122_ sky130_fd_sc_hd__a22o_1
X_09043_ net1150 top.WB.CPU_DAT_O\[14\] net292 vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_111_Right_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06186_ _02565_ _02972_ _03055_ vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__or3_1
Xhold410 net59 vssd1 vssd1 vccd1 vccd1 net1363 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06343__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08215__C1 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05748__A _02539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold454 net69 vssd1 vssd1 vccd1 vccd1 net1407 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_6_0_clk_X clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold443 top.path\[57\] vssd1 vssd1 vccd1 vccd1 net1396 sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 top.path\[117\] vssd1 vssd1 vccd1 vccd1 net1385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold421 top.cb_syn.char_path\[105\] vssd1 vssd1 vccd1 vccd1 net1374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 net67 vssd1 vssd1 vccd1 vccd1 net1429 sky130_fd_sc_hd__dlygate4sd3_1
Xhold465 net96 vssd1 vssd1 vccd1 vccd1 net1418 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold487 top.hTree.tree_reg\[21\] vssd1 vssd1 vccd1 vccd1 net1440 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06241__B2 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold498 top.cb_syn.curr_index\[2\] vssd1 vssd1 vccd1 vccd1 net1451 sky130_fd_sc_hd__dlygate4sd3_1
X_09945_ net741 net581 vssd1 vssd1 vccd1 vccd1 _00559_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout580_A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout678_A net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09876_ net761 net601 vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__and2_1
XANTENNA__06792__A2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout299_X net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08827_ top.path\[12\] top.path\[13\] top.path\[14\] top.path\[15\] net527 top.translation.index\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05010_ sky130_fd_sc_hd__mux4_1
XFILLER_38_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout466_X net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout845_A net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08758_ net522 _04940_ vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__and2_1
X_08689_ _02511_ _04880_ vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__nand2_1
X_07709_ net263 _04272_ _04273_ net1015 net446 vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__a32o_1
XFILLER_54_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05504__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10720_ clknet_leaf_112_clk _01319_ _00139_ vssd1 vssd1 vccd1 vccd1 top.path\[96\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_109_Left_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10651_ clknet_leaf_60_clk _01250_ _00070_ vssd1 vssd1 vccd1 vccd1 top.hist_addr\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout800_X net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09246__A1 top.cb_syn.char_index\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10582_ net746 net586 vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__and2_1
X_11203_ clknet_leaf_10_clk _01751_ _00558_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[105\]
+ sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_118_Left_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_61_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11134_ clknet_leaf_13_clk _01682_ _00489_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[36\]
+ sky130_fd_sc_hd__dfrtp_2
X_11065_ clknet_leaf_43_clk _01613_ _00420_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[95\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_76_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10016_ net819 net659 vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__and2_1
XFILLER_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05680__X _02755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11967_ net63 vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_47_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10918_ clknet_leaf_32_clk _01473_ _00273_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.i\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_44_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10849_ clknet_leaf_108_clk _01435_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_119_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_14_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08996__A0 top.WB.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06040_ _02457_ _02930_ vssd1 vssd1 vccd1 vccd1 _02931_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_29_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07991_ top.cb_syn.zeroes\[0\] _02531_ _04484_ vssd1 vssd1 vccd1 vccd1 _04494_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06223__B2 top.findLeastValue.histo_index\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xfanout208 net210 vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__clkbuf_4
Xfanout219 _05262_ vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_4_7_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_7_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__06774__A2 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09730_ net769 net609 vssd1 vssd1 vccd1 vccd1 _00344_ sky130_fd_sc_hd__and2_1
X_06942_ top.compVal\[12\] top.findLeastValue.val1\[12\] net162 vssd1 vssd1 vccd1
+ vccd1 _03613_ sky130_fd_sc_hd__mux2_1
X_09661_ net785 net625 vssd1 vssd1 vccd1 vccd1 _00275_ sky130_fd_sc_hd__and2_1
X_06873_ _02546_ _03011_ _03576_ _03567_ net1501 vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__a32o_1
X_08612_ top.cb_syn.num_lefts\[4\] _04829_ vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__nand2_1
X_05824_ top.sram_interface.write_counter_FLV\[1\] top.sram_interface.write_counter_FLV\[0\]
+ net289 vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__and3_1
X_09592_ net847 net687 vssd1 vssd1 vccd1 vccd1 _00206_ sky130_fd_sc_hd__and2_1
XANTENNA__08818__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08543_ net1253 top.cb_syn.char_path_n\[33\] net233 vssd1 vssd1 vccd1 vccd1 _01551_
+ sky130_fd_sc_hd__mux2_1
X_05755_ top.compVal\[39\] net173 _02783_ top.WB.CPU_DAT_O\[7\] vssd1 vssd1 vccd1
+ vccd1 _02324_ sky130_fd_sc_hd__a22o_1
XANTENNA__07487__A0 top.cb_syn.char_path_n\[32\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout259_A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05686_ net450 top.WB.prev_BUSY_O vssd1 vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__and2_2
X_08474_ net1204 top.cb_syn.char_path_n\[102\] net226 vssd1 vssd1 vccd1 vccd1 _01620_
+ sky130_fd_sc_hd__mux2_1
X_07425_ net354 _04005_ _04022_ _04001_ vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__o211a_1
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08436__C1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07356_ _03754_ _03756_ vssd1 vssd1 vccd1 vccd1 _03971_ sky130_fd_sc_hd__xnor2_1
X_06307_ net1398 net142 _03170_ net160 vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__a22o_1
X_07287_ _03813_ _03922_ _03794_ vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08987__A0 top.WB.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06238_ top.cb_syn.char_index\[0\] _03095_ _03097_ net478 vssd1 vssd1 vccd1 vccd1
+ _03106_ sky130_fd_sc_hd__o211a_1
X_09026_ net1081 top.WB.CPU_DAT_O\[31\] net291 vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__mux2_1
XFILLER_117_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06169_ net497 net412 _03013_ net498 vssd1 vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__a22o_1
Xhold262 top.cb_syn.char_path\[86\] vssd1 vssd1 vccd1 vccd1 net1215 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 top.cb_syn.char_path\[102\] vssd1 vssd1 vccd1 vccd1 net1204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold240 top.cb_syn.char_path\[9\] vssd1 vssd1 vccd1 vccd1 net1193 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 top.cb_syn.char_path\[20\] vssd1 vssd1 vccd1 vccd1 net1248 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07693__A net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold284 top.path\[63\] vssd1 vssd1 vccd1 vccd1 net1237 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 top.path\[28\] vssd1 vssd1 vccd1 vccd1 net1226 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout720 net722 vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__clkbuf_4
X_09928_ net775 net615 vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__and2_1
Xfanout742 net744 vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__clkbuf_2
Xfanout731 net734 vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__buf_1
Xfanout775 net776 vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__clkbuf_2
Xfanout753 net754 vssd1 vssd1 vccd1 vccd1 net753 sky130_fd_sc_hd__buf_1
Xfanout764 net767 vssd1 vssd1 vccd1 vccd1 net764 sky130_fd_sc_hd__buf_1
Xfanout786 net807 vssd1 vssd1 vccd1 vccd1 net786 sky130_fd_sc_hd__clkbuf_2
XFILLER_105_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout797 net800 vssd1 vssd1 vccd1 vccd1 net797 sky130_fd_sc_hd__clkbuf_2
XFILLER_92_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09859_ net771 net611 vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__and2_1
XFILLER_73_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11821_ clknet_leaf_56_clk _02337_ _01176_ vssd1 vssd1 vccd1 vccd1 top.TRN_char_index\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ clknet_leaf_95_clk _02285_ _01107_ vssd1 vssd1 vccd1 vccd1 top.compVal\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11683_ clknet_leaf_61_clk _02216_ _01038_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10703_ clknet_leaf_11_clk _01302_ _00122_ vssd1 vssd1 vccd1 vccd1 top.path\[79\]
+ sky130_fd_sc_hd__dfrtp_1
X_10634_ clknet_leaf_49_clk _00038_ _00053_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.word_cnt\[0\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_62_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08978__A0 top.WB.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07650__A0 top.findLeastValue.least1\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10565_ net808 net648 vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__and2_1
XFILLER_5_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10496_ net815 net655 vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_114_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11117_ clknet_leaf_22_clk _01665_ _00472_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05835__B _02843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11048_ clknet_leaf_10_clk _01596_ _00403_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[78\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput8 DAT_I[15] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XANTENNA__05716__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06781__A_N net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05540_ top.cb_syn.char_path\[23\] net559 net314 top.cb_syn.char_path\[119\] vssd1
+ vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__a22o_1
XFILLER_32_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_05471_ net478 net561 vssd1 vssd1 vccd1 vccd1 _02579_ sky130_fd_sc_hd__and2_1
XANTENNA__06141__B1 top.findLeastValue.histo_index\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11361__Q top.findLeastValue.sum\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05495__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08190_ top.cb_syn.char_path_n\[74\] net199 _04622_ vssd1 vssd1 vccd1 vccd1 _01720_
+ sky130_fd_sc_hd__o21a_1
X_07210_ _03865_ _03866_ top.findLeastValue.sum\[44\] net276 vssd1 vssd1 vccd1 vccd1
+ _01940_ sky130_fd_sc_hd__a2bb2o_1
X_07141_ top.findLeastValue.val1\[16\] top.findLeastValue.val2\[16\] vssd1 vssd1 vccd1
+ vccd1 _03799_ sky130_fd_sc_hd__xnor2_2
XANTENNA__08969__A0 top.WB.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07072_ top.findLeastValue.val1\[11\] top.findLeastValue.val2\[11\] vssd1 vssd1 vccd1
+ vccd1 _03730_ sky130_fd_sc_hd__xnor2_1
XFILLER_114_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08816__S0 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06023_ net1591 top.WB.CPU_DAT_O\[12\] net356 vssd1 vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__mux2_1
XFILLER_114_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09394__B1 _05272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05585__X _02676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07974_ top.cb_syn.h_element\[63\] _02553_ vssd1 vssd1 vccd1 vccd1 _04478_ sky130_fd_sc_hd__nor2_2
XANTENNA__09217__B top.controller.fin_reg\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05955__A0 top.WB.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05464__C net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09713_ net792 net632 vssd1 vssd1 vccd1 vccd1 _00327_ sky130_fd_sc_hd__and2_1
X_06925_ top.findLeastValue.val2\[21\] net146 net120 _03604_ vssd1 vssd1 vccd1 vccd1
+ _01963_ sky130_fd_sc_hd__o22a_1
X_09644_ net803 net643 vssd1 vssd1 vccd1 vccd1 _00258_ sky130_fd_sc_hd__and2_1
XANTENNA__08548__S net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06856_ _03567_ _03569_ vssd1 vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout376_A net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06857__A net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05807_ top.sram_interface.counter_HTREE\[0\] _02826_ vssd1 vssd1 vccd1 vccd1 _02827_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_2_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10379__A net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout543_A net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09575_ net819 net659 vssd1 vssd1 vccd1 vccd1 _00189_ sky130_fd_sc_hd__and2_1
X_06787_ top.findLeastValue.val1\[43\] net131 net115 top.compVal\[43\] vssd1 vssd1
+ vccd1 vccd1 _02051_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout164_X net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05738_ top.findLeastValue.startup _02772_ net470 vssd1 vssd1 vccd1 vccd1 _02773_
+ sky130_fd_sc_hd__o21ai_4
X_08526_ net1268 top.cb_syn.char_path_n\[50\] net223 vssd1 vssd1 vccd1 vccd1 _01568_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout710_A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout331_X net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08457_ net1140 top.cb_syn.char_path_n\[119\] net229 vssd1 vssd1 vccd1 vccd1 _01637_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09887__B net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05669_ top.hTree.node_reg\[34\] net311 _02745_ net480 vssd1 vssd1 vccd1 vccd1 _02746_
+ sky130_fd_sc_hd__a22o_1
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07408_ _03994_ _03996_ _04006_ _04007_ vssd1 vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__a22o_1
XANTENNA__08409__C1 _02504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_109_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_08388_ net505 _04742_ _04745_ _04746_ _02503_ vssd1 vssd1 vccd1 vccd1 _04747_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_21_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07339_ _03733_ _03734_ _03954_ vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__nand3_1
X_10350_ net870 net710 vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__and2_1
XANTENNA__06435__A1 top.header_synthesis.enable vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10281_ net725 net565 vssd1 vssd1 vccd1 vccd1 _00895_ sky130_fd_sc_hd__and2_1
X_09009_ top.WB.CPU_DAT_O\[16\] net1344 net317 vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__mux2_1
XFILLER_105_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05495__X _02601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07627__S net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_05_888 vssd1 vssd1 vccd1 vccd1 team_05_888/HI gpio_out[3] sky130_fd_sc_hd__conb_1
Xfanout550 top.sram_interface.word_cnt\[5\] vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__buf_2
XANTENNA__05946__A0 top.WB.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_05_899 vssd1 vssd1 vccd1 vccd1 team_05_899/HI gpio_out[14] sky130_fd_sc_hd__conb_1
Xfanout561 net562 vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__buf_2
Xfanout583 net584 vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__buf_1
XFILLER_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout572 net574 vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__clkbuf_2
Xfanout594 net597 vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__buf_1
XFILLER_100_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08360__A1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ clknet_leaf_91_clk _02321_ _01159_ vssd1 vssd1 vccd1 vccd1 top.compVal\[36\]
+ sky130_fd_sc_hd__dfrtp_4
X_11735_ clknet_leaf_50_clk _02268_ _01090_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.CB_write_counter\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_42_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_14_0_clk_X clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11666_ clknet_leaf_45_clk _02199_ _01021_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_11597_ clknet_leaf_43_clk _02145_ _00952_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10617_ net810 net650 vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__and2_1
XANTENNA__06652__D _03440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07623__A0 top.findLeastValue.least1\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10548_ net834 net674 vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__and2_1
X_10479_ net861 net701 vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__and2_1
XANTENNA__05937__A0 top.WB.CPU_DAT_O\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11356__Q top.findLeastValue.sum\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06710_ _02432_ top.findLeastValue.val2\[17\] top.findLeastValue.val2\[16\] _02433_
+ _03497_ vssd1 vssd1 vccd1 vccd1 _03498_ sky130_fd_sc_hd__o221ai_2
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07690_ net490 _04254_ vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__or2_1
X_06641_ net494 top.compVal\[26\] top.compVal\[25\] top.compVal\[24\] vssd1 vssd1
+ vccd1 vccd1 _03430_ sky130_fd_sc_hd__or4_1
X_09360_ net1056 net239 net218 _04346_ vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__a22o_1
X_06572_ _03358_ _03359_ _03360_ vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__a21o_1
X_09291_ _03992_ net298 vssd1 vssd1 vccd1 vccd1 top.dut.bit_buf_next\[7\] sky130_fd_sc_hd__and2_1
X_05523_ _02622_ _02623_ net476 vssd1 vssd1 vccd1 vccd1 _02624_ sky130_fd_sc_hd__o21a_1
X_08311_ top.cb_syn.char_path_n\[14\] net373 net333 top.cb_syn.char_path_n\[12\] net178
+ vssd1 vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__a221o_1
XANTENNA__09300__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05454_ net555 net547 vssd1 vssd1 vccd1 vccd1 _02562_ sky130_fd_sc_hd__or2_2
X_08242_ top.cb_syn.char_path_n\[48\] net197 _04648_ vssd1 vssd1 vccd1 vccd1 _01694_
+ sky130_fd_sc_hd__o21a_1
XFILLER_119_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__08406__A2 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08173_ top.cb_syn.char_path_n\[83\] net382 net341 top.cb_syn.char_path_n\[81\] net186
+ vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__a221o_1
X_05385_ top.findLeastValue.val2\[15\] vssd1 vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout124_A net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08811__C1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07124_ _03723_ _03776_ _03781_ vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__o21a_2
X_07055_ top.findLeastValue.val1\[14\] top.findLeastValue.val2\[14\] vssd1 vssd1 vccd1
+ vccd1 _03713_ sky130_fd_sc_hd__or2_1
X_06006_ net1614 top.WB.CPU_DAT_O\[29\] net358 vssd1 vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__mux2_1
XANTENNA__06351__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_7_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05928__A0 top.WB.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07957_ net1484 _04468_ _04461_ vssd1 vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__mux2_1
XFILLER_87_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06908_ top.compVal\[29\] top.findLeastValue.val1\[29\] net163 vssd1 vssd1 vccd1
+ vccd1 _03596_ sky130_fd_sc_hd__mux2_1
X_07888_ net440 net1569 net251 top.findLeastValue.sum\[11\] _04416_ vssd1 vssd1 vccd1
+ vccd1 _01816_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout546_X net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06839_ top.findLeastValue.least1\[5\] net498 _03424_ vssd1 vssd1 vccd1 vccd1 _03559_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09627_ net755 net595 vssd1 vssd1 vccd1 vccd1 _00241_ sky130_fd_sc_hd__and2_1
X_09558_ net843 net683 vssd1 vssd1 vccd1 vccd1 _00172_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_54_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08509_ net1128 top.cb_syn.char_path_n\[67\] net227 vssd1 vssd1 vccd1 vccd1 _01585_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11520_ clknet_leaf_64_clk _02068_ _00875_ vssd1 vssd1 vccd1 vccd1 top.cw1\[3\] sky130_fd_sc_hd__dfrtp_1
X_09489_ net733 net573 vssd1 vssd1 vccd1 vccd1 _00103_ sky130_fd_sc_hd__and2_1
XANTENNA__10556__B net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07853__B1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11451_ clknet_leaf_70_clk _01999_ _00806_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least2\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10402_ net792 net632 vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__and2_1
X_11382_ clknet_leaf_86_clk _01930_ _00737_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_109_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10333_ net845 net685 vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__and2_1
XANTENNA__06959__A2 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09358__B1 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10264_ net867 net707 vssd1 vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__and2_1
XANTENNA__08042__A net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05631__A2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10195_ net858 net698 vssd1 vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__and2_1
XANTENNA__07908__B2 top.findLeastValue.sum\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08581__A1 top.cb_syn.char_index\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout391 net393 vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__clkbuf_4
Xfanout380 net382 vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_109_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08333__B2 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09601__A net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08097__B1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07519__S0 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07820__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__07844__A0 top.findLeastValue.sum\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11718_ clknet_leaf_122_clk _02251_ _01073_ vssd1 vssd1 vccd1 vccd1 top.path\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput11 DAT_I[18] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
Xinput22 DAT_I[28] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
X_11649_ clknet_leaf_113_clk _02182_ _01004_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput44 nrst vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_2
Xinput33 DAT_I[9] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
XFILLER_116_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09349__B1 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08860_ top.translation.resEn _05040_ vssd1 vssd1 vccd1 vccd1 _05042_ sky130_fd_sc_hd__or2_1
X_07811_ net484 _04353_ vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_4_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07791__A net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08791_ _02522_ _04939_ _04941_ _02521_ vssd1 vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__o31a_1
X_07742_ net429 _04298_ _04299_ net260 vssd1 vssd1 vccd1 vccd1 _04300_ sky130_fd_sc_hd__o211a_1
X_07673_ net457 net1064 net257 _04243_ vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_84_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09412_ net406 _04221_ vssd1 vssd1 vccd1 vccd1 _05285_ sky130_fd_sc_hd__nand2_1
XFILLER_52_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06624_ _03410_ _03411_ _03412_ vssd1 vssd1 vccd1 vccd1 _03413_ sky130_fd_sc_hd__and3b_1
XANTENNA__05461__D net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07730__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09343_ net1071 net237 net214 _04414_ vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__a22o_1
XFILLER_80_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout241_A net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout339_A net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06555_ _03341_ _03342_ _03343_ _03340_ vssd1 vssd1 vccd1 vccd1 _03344_ sky130_fd_sc_hd__or4b_1
X_09274_ _02533_ _05222_ vssd1 vssd1 vccd1 vccd1 _05226_ sky130_fd_sc_hd__nand2_1
X_05506_ net456 top.hTree.node_reg\[61\] net362 net422 top.hTree.node_reg\[29\] vssd1
+ vssd1 vccd1 vccd1 _02610_ sky130_fd_sc_hd__a32o_1
XANTENNA__07835__A0 top.findLeastValue.sum\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06486_ net1534 _03287_ vssd1 vssd1 vccd1 vccd1 _03300_ sky130_fd_sc_hd__nor2_1
XFILLER_21_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05437_ net499 net500 top.findLeastValue.histo_index\[3\] net502 vssd1 vssd1 vccd1
+ vccd1 _02545_ sky130_fd_sc_hd__or4_1
X_08225_ top.cb_syn.char_path_n\[57\] net384 net343 top.cb_syn.char_path_n\[55\] net188
+ vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_31_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08156_ top.cb_syn.char_path_n\[91\] net210 _04605_ vssd1 vssd1 vccd1 vccd1 _01737_
+ sky130_fd_sc_hd__o21a_1
X_05368_ top.findLeastValue.least2\[4\] vssd1 vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__inv_2
XANTENNA__05861__A2 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08561__S net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07107_ _03742_ _03743_ vssd1 vssd1 vccd1 vccd1 _03765_ sky130_fd_sc_hd__nand2b_1
X_08087_ top.cb_syn.char_path_n\[126\] net385 net344 top.cb_syn.char_path_n\[124\]
+ net189 vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__a221o_1
XANTENNA__10392__A net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05299_ top.compVal\[44\] vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_95_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05613__A2 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07038_ top.findLeastValue.val1\[29\] top.findLeastValue.val2\[29\] vssd1 vssd1 vccd1
+ vccd1 _03696_ sky130_fd_sc_hd__and2_1
XANTENNA__07366__A2 _03553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08989_ top.WB.CPU_DAT_O\[3\] net1197 net324 vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__mux2_1
X_10951_ clknet_leaf_33_clk _01506_ _00306_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.num_lefts\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10882_ clknet_leaf_47_clk _01459_ _00237_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.TRN_counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11503_ clknet_leaf_90_clk _02051_ _00858_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[43\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_8_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__05852__A2 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11434_ clknet_leaf_89_clk _01982_ _00789_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[40\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_59_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_100_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_100_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11365_ clknet_leaf_101_clk _01913_ _00720_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05396__A net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11296_ clknet_leaf_83_clk _01844_ _00651_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[39\]
+ sky130_fd_sc_hd__dfrtp_1
X_10316_ net764 net604 vssd1 vssd1 vccd1 vccd1 _00930_ sky130_fd_sc_hd__and2_1
XFILLER_98_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10247_ net841 net681 vssd1 vssd1 vccd1 vccd1 _00861_ sky130_fd_sc_hd__and2_1
XANTENNA__07815__S net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10178_ net828 net668 vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__and2_1
XANTENNA__06868__A1 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__10477__A net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06340_ top.hist_data_o\[29\] _03193_ _03199_ vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__o21ba_1
X_06271_ net549 _02573_ _03132_ net368 net503 vssd1 vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__a32o_1
X_08010_ _02502_ _04512_ vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__nor2_1
XANTENNA__05843__A2 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08381__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold603 _01832_ vssd1 vssd1 vccd1 vccd1 net1556 sky130_fd_sc_hd__dlygate4sd3_1
Xhold636 top.controller.fin_reg\[7\] vssd1 vssd1 vccd1 vccd1 net1589 sky130_fd_sc_hd__dlygate4sd3_1
Xhold614 top.histogram.total\[19\] vssd1 vssd1 vccd1 vccd1 net1567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold625 top.hTree.tree_reg\[6\] vssd1 vssd1 vccd1 vccd1 net1578 sky130_fd_sc_hd__dlygate4sd3_1
Xhold647 top.histogram.state\[3\] vssd1 vssd1 vccd1 vccd1 net1600 sky130_fd_sc_hd__dlygate4sd3_1
X_09961_ net777 net617 vssd1 vssd1 vccd1 vccd1 _00575_ sky130_fd_sc_hd__and2_1
Xhold669 top.sram_interface.counter_HTREE\[3\] vssd1 vssd1 vccd1 vccd1 net1622 sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 top.findLeastValue.sum\[31\] vssd1 vssd1 vccd1 vccd1 net1611 sky130_fd_sc_hd__dlygate4sd3_1
X_08912_ _04187_ _05065_ _05078_ vssd1 vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__or3b_1
X_09892_ net774 net614 vssd1 vssd1 vccd1 vccd1 _00506_ sky130_fd_sc_hd__and2_1
XANTENNA__07348__A2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout191_A net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08843_ net434 _05012_ _05025_ vssd1 vssd1 vccd1 vccd1 _05026_ sky130_fd_sc_hd__o21a_1
X_05986_ top.sram_interface.init_counter\[7\] _02914_ vssd1 vssd1 vccd1 vccd1 _02918_
+ sky130_fd_sc_hd__nor2_1
X_08774_ top.path\[114\] top.path\[115\] net528 vssd1 vssd1 vccd1 vccd1 _04957_ sky130_fd_sc_hd__mux2_1
X_11892__919 vssd1 vssd1 vccd1 vccd1 _11892__919/HI net919 sky130_fd_sc_hd__conb_1
X_07725_ top.hTree.tree_reg\[43\] top.findLeastValue.sum\[43\] net247 vssd1 vssd1
+ vccd1 vccd1 _04286_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout456_A net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_2_0_clk_X clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07656_ top.findLeastValue.least1\[1\] top.hTree.tree_reg\[56\] net280 vssd1 vssd1
+ vccd1 vccd1 _04230_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout623_A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07587_ _04148_ _04173_ vssd1 vssd1 vccd1 vccd1 _04174_ sky130_fd_sc_hd__nand2_1
XANTENNA__10387__A net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06607_ top.compVal\[40\] _02462_ vssd1 vssd1 vccd1 vccd1 _03396_ sky130_fd_sc_hd__or2_1
X_09326_ _02786_ net431 net36 net325 vssd1 vssd1 vccd1 vccd1 top.controller.fin_TRN
+ sky130_fd_sc_hd__and4b_1
X_06538_ _02419_ top.findLeastValue.val1\[31\] vssd1 vssd1 vccd1 vccd1 _03327_ sky130_fd_sc_hd__and2_1
XANTENNA__07808__B1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09257_ top.header_synthesis.write_zeroes _04922_ net519 vssd1 vssd1 vccd1 vccd1
+ _05214_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_97_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08208_ top.cb_syn.char_path_n\[65\] net209 _04631_ vssd1 vssd1 vccd1 vccd1 _01711_
+ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout509_X net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06469_ top.histogram.total\[29\] top.histogram.total\[28\] _03291_ vssd1 vssd1 vccd1
+ vccd1 _03292_ sky130_fd_sc_hd__and3_1
X_09188_ _02541_ _02544_ _02591_ vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08616__A_N _04826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05834__A2 _02843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08139_ top.cb_syn.char_path_n\[100\] net380 net340 top.cb_syn.char_path_n\[98\]
+ net184 vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__a221o_1
X_11150_ clknet_leaf_22_clk _01698_ _00505_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[52\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout878_X net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__05598__B2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10101_ net816 net656 vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__and2_1
XANTENNA__06795__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11081_ clknet_leaf_6_clk _01629_ _00436_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[111\]
+ sky130_fd_sc_hd__dfrtp_1
X_10032_ net839 net679 vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__and2_1
XFILLER_102_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06759__B _03546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input17_A DAT_I[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10934_ clknet_leaf_35_clk _01489_ _00289_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.cb_enable
+ sky130_fd_sc_hd__dfrtp_1
X_10865_ clknet_leaf_47_clk _01451_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_14_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10796_ clknet_leaf_57_clk _00036_ _00215_ vssd1 vssd1 vccd1 vccd1 top.histogram.wr_r_en\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__06078__A2 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05397__Y _02505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11417_ clknet_leaf_98_clk _01965_ _00772_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[23\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_117_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11348_ clknet_leaf_92_clk _01896_ _00703_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__06786__B1 net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06250__A2 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11279_ clknet_leaf_78_clk _01827_ _00634_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_79_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06002__A2 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05840_ net494 net169 net155 top.WB.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1 _02302_
+ sky130_fd_sc_hd__a22o_1
X_07510_ top.cb_syn.char_path_n\[96\] top.cb_syn.char_path_n\[95\] top.cb_syn.char_path_n\[94\]
+ top.cb_syn.char_path_n\[93\] net402 net353 vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__mux4_1
X_05771_ _02787_ _02791_ vssd1 vssd1 vccd1 vccd1 _02792_ sky130_fd_sc_hd__nor2_1
XANTENNA__05761__A1 top.compVal\[33\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05761__B2 top.WB.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08490_ net1215 top.cb_syn.char_path_n\[86\] net233 vssd1 vssd1 vccd1 vccd1 _01604_
+ sky130_fd_sc_hd__mux2_1
X_07441_ _04027_ _04035_ net354 vssd1 vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07502__A2 top.cb_syn.char_path_n\[42\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07372_ net1572 net135 _03547_ net127 _03979_ vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__a32o_1
XFILLER_50_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09111_ _05126_ _05129_ vssd1 vssd1 vccd1 vccd1 _00045_ sky130_fd_sc_hd__nand2_1
X_06323_ top.hist_data_o\[17\] _03185_ vssd1 vssd1 vccd1 vccd1 _03186_ sky130_fd_sc_hd__and2_1
X_06254_ _02418_ _03120_ vssd1 vssd1 vccd1 vccd1 _03121_ sky130_fd_sc_hd__nor2_1
X_09042_ net1067 top.WB.CPU_DAT_O\[15\] net292 vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__mux2_1
X_06185_ top.TRN_char_index\[4\] _02971_ vssd1 vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__nor2_1
Xhold411 top.path\[56\] vssd1 vssd1 vccd1 vccd1 net1364 sky130_fd_sc_hd__dlygate4sd3_1
Xhold400 _01847_ vssd1 vssd1 vccd1 vccd1 net1353 sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 top.cb_syn.char_path\[121\] vssd1 vssd1 vccd1 vccd1 net1375 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout204_A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold433 top.path\[112\] vssd1 vssd1 vccd1 vccd1 net1386 sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 top.path\[104\] vssd1 vssd1 vccd1 vccd1 net1397 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06777__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold455 top.hTree.tree_reg\[31\] vssd1 vssd1 vccd1 vccd1 net1408 sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 top.cb_syn.char_path\[46\] vssd1 vssd1 vccd1 vccd1 net1419 sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 top.path\[118\] vssd1 vssd1 vccd1 vccd1 net1430 sky130_fd_sc_hd__dlygate4sd3_1
Xhold488 top.hTree.tree_reg\[34\] vssd1 vssd1 vccd1 vccd1 net1441 sky130_fd_sc_hd__dlygate4sd3_1
X_09944_ net741 net581 vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__and2_1
Xhold499 top.hTree.tree_reg\[4\] vssd1 vssd1 vccd1 vccd1 net1452 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09875_ net761 net601 vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__and2_1
XANTENNA_input9_A DAT_I[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout194_X net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_08826_ net434 _05007_ _05008_ vssd1 vssd1 vccd1 vccd1 _05009_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout573_A net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05969_ top.sram_interface.init_counter\[2\] top.sram_interface.init_counter\[1\]
+ _02903_ vssd1 vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout838_A net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout361_X net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05752__B2 top.WB.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08757_ top.path\[108\] top.path\[109\] top.path\[110\] top.path\[111\] net527 net523
+ vssd1 vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout740_A net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08688_ top.cb_syn.zeroes\[6\] _04887_ _04884_ vssd1 vssd1 vccd1 vccd1 _01487_ sky130_fd_sc_hd__o21a_1
X_07708_ net490 _04269_ vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__or2_1
XFILLER_26_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08151__C1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07639_ top.findLeastValue.least1\[4\] net248 _04214_ vssd1 vssd1 vccd1 vccd1 _04216_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_14_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout626_X net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10650_ clknet_leaf_60_clk _01249_ _00069_ vssd1 vssd1 vccd1 vccd1 top.hist_addr\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09309_ _05239_ _05240_ _05242_ _05243_ vssd1 vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_101_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10581_ net746 net586 vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__and2_1
XANTENNA__05498__X _02603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11202_ clknet_leaf_10_clk _01750_ _00557_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[104\]
+ sky130_fd_sc_hd__dfrtp_2
X_11133_ clknet_leaf_13_clk _01681_ _00488_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_110_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06783__A3 _03547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11064_ clknet_leaf_42_clk _01612_ _00419_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[94\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09182__B2 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10015_ net819 net659 vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__and2_1
XFILLER_48_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05961__X _02899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07732__A2 _04290_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10917_ clknet_leaf_38_clk top.header_synthesis.next_char_added _00272_ vssd1 vssd1
+ vccd1 vccd1 top.header_synthesis.char_added sky130_fd_sc_hd__dfrtp_1
XFILLER_44_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08924__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10848_ clknet_leaf_107_clk _01434_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10779_ clknet_leaf_46_clk _01378_ _00198_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11359__Q top.findLeastValue.sum\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07990_ _04485_ _04486_ _04487_ vssd1 vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__or3_1
XFILLER_99_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout209 net210 vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__buf_2
X_06941_ top.findLeastValue.val2\[13\] net147 net121 _03612_ vssd1 vssd1 vccd1 vccd1
+ _01955_ sky130_fd_sc_hd__o22a_1
X_09660_ net782 net622 vssd1 vssd1 vccd1 vccd1 _00274_ sky130_fd_sc_hd__and2_1
X_08611_ _04829_ vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__inv_2
X_06872_ net502 _03567_ _03576_ _03131_ vssd1 vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__a22o_1
X_05823_ net556 _02778_ _02836_ net423 _02549_ vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__a2111oi_1
X_09591_ net846 net686 vssd1 vssd1 vccd1 vccd1 _00205_ sky130_fd_sc_hd__and2_1
XFILLER_54_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08542_ net1322 top.cb_syn.char_path_n\[34\] net228 vssd1 vssd1 vccd1 vccd1 _01552_
+ sky130_fd_sc_hd__mux2_1
X_05754_ top.compVal\[40\] net172 net158 top.WB.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1
+ _02325_ sky130_fd_sc_hd__a22o_1
XFILLER_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08133__C1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08473_ net1285 top.cb_syn.char_path_n\[103\] net225 vssd1 vssd1 vccd1 vccd1 _01621_
+ sky130_fd_sc_hd__mux2_1
X_07424_ top.dut.bits_in_buf_next\[1\] _03990_ vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__or2_1
X_05685_ top.WB.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__nand2_2
XANTENNA__05498__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout154_A net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11822__Q top.WB.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07239__A1 _03817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07355_ _03760_ net270 _03970_ net275 top.findLeastValue.sum\[3\] vssd1 vssd1 vccd1
+ vccd1 _01899_ sky130_fd_sc_hd__a32o_1
X_06306_ net471 _03163_ _03169_ vssd1 vssd1 vccd1 vccd1 _03170_ sky130_fd_sc_hd__a21o_1
X_07286_ _03782_ _03807_ vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout419_A net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06237_ top.cb_syn.max_index\[4\] _03025_ _03027_ top.hTree.nullSumIndex\[3\] vssd1
+ vssd1 vccd1 vccd1 _03105_ sky130_fd_sc_hd__a22o_1
X_09025_ top.WB.CPU_DAT_O\[0\] net1130 net320 vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__mux2_1
XANTENNA__07974__A top.cb_syn.h_element\[63\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05670__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout690_A net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06168_ net1324 net141 _03038_ net159 vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__a22o_1
Xhold230 top.histogram.sram_out\[29\] vssd1 vssd1 vccd1 vccd1 net1183 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09400__A2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold252 top.cb_syn.char_path\[15\] vssd1 vssd1 vccd1 vccd1 net1205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 net104 vssd1 vssd1 vccd1 vccd1 net1194 sky130_fd_sc_hd__dlygate4sd3_1
X_06099_ top.TRN_char_index\[4\] _02971_ vssd1 vssd1 vccd1 vccd1 _02972_ sky130_fd_sc_hd__and2_1
Xhold296 top.cb_syn.char_path\[58\] vssd1 vssd1 vccd1 vccd1 net1249 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout788_A net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold274 top.cb_syn.char_path\[49\] vssd1 vssd1 vccd1 vccd1 net1227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 top.cb_syn.char_path\[11\] vssd1 vssd1 vccd1 vccd1 net1216 sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 top.cb_syn.char_path\[40\] vssd1 vssd1 vccd1 vccd1 net1238 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout721 net722 vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__clkbuf_2
Xfanout710 net717 vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06765__A3 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09927_ net776 net616 vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__and2_1
Xfanout732 net734 vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09164__A1 _03270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout776 net807 vssd1 vssd1 vccd1 vccd1 net776 sky130_fd_sc_hd__clkbuf_2
Xfanout743 net744 vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__buf_1
Xfanout765 net766 vssd1 vssd1 vccd1 vccd1 net765 sky130_fd_sc_hd__clkbuf_2
Xfanout754 net757 vssd1 vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__buf_1
Xfanout798 net799 vssd1 vssd1 vccd1 vccd1 net798 sky130_fd_sc_hd__clkbuf_2
Xfanout787 net791 vssd1 vssd1 vccd1 vccd1 net787 sky130_fd_sc_hd__clkbuf_2
X_09858_ net772 net612 vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__and2_1
XFILLER_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09789_ net742 net582 vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__and2_1
X_08809_ top.path\[58\] top.path\[59\] net525 vssd1 vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__mux2_1
X_11820_ clknet_leaf_56_clk _02336_ _01175_ vssd1 vssd1 vccd1 vccd1 top.TRN_char_index\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_44_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ clknet_leaf_95_clk _02284_ _01106_ vssd1 vssd1 vccd1 vccd1 top.compVal\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05489__B1 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_80_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_clk sky130_fd_sc_hd__clkbuf_8
X_10702_ clknet_leaf_3_clk _01301_ _00121_ vssd1 vssd1 vccd1 vccd1 top.path\[78\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_41_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11682_ clknet_leaf_61_clk _02215_ _01037_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_10633_ net852 net692 vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_62_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10564_ net808 net648 vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__and2_1
XANTENNA__05661__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10495_ net815 net655 vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_114_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11116_ clknet_leaf_22_clk _01664_ _00471_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[18\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__09155__A1 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_10_0_clk_X clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11047_ clknet_leaf_4_clk _01595_ _00402_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[77\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_92_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05716__B2 top.WB.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput9 DAT_I[16] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06913__B1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_71_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_60_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05470_ net478 _02577_ vssd1 vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__and2_2
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07140_ _03794_ _03797_ vssd1 vssd1 vccd1 vccd1 _03798_ sky130_fd_sc_hd__or2_1
X_07071_ _03727_ _03728_ vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__nand2_1
XANTENNA__06902__S net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06022_ net1666 top.WB.CPU_DAT_O\[13\] net356 vssd1 vssd1 vccd1 vccd1 _02188_ sky130_fd_sc_hd__mux2_1
XANTENNA__08816__S1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09712_ net787 net627 vssd1 vssd1 vccd1 vccd1 _00326_ sky130_fd_sc_hd__and2_1
X_07973_ net446 net286 net1278 vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__o21bai_1
XANTENNA__08354__C1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08829__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06924_ top.compVal\[21\] top.findLeastValue.val1\[21\] net161 vssd1 vssd1 vccd1
+ vccd1 _03604_ sky130_fd_sc_hd__mux2_1
X_09643_ net804 net644 vssd1 vssd1 vccd1 vccd1 _00257_ sky130_fd_sc_hd__and2_1
X_06855_ net500 _03109_ vssd1 vssd1 vccd1 vccd1 _03569_ sky130_fd_sc_hd__nand2_1
XFILLER_67_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout271_A net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05806_ _02822_ _02825_ _02818_ _02820_ vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__and4bb_1
X_09574_ net794 net634 vssd1 vssd1 vccd1 vccd1 _00188_ sky130_fd_sc_hd__and2_1
XANTENNA__05707__B2 top.WB.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10379__B net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06349__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08525_ net1230 top.cb_syn.char_path_n\[51\] net223 vssd1 vssd1 vccd1 vccd1 _01569_
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06786_ top.findLeastValue.val1\[44\] net132 net116 top.compVal\[44\] vssd1 vssd1
+ vccd1 vccd1 _02052_ sky130_fd_sc_hd__o22a_1
XANTENNA_clkbuf_leaf_60_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_62_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout536_A top.cb_syn.curr_state\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05737_ top.findLeastValue.histo_index\[7\] _02769_ _02771_ _02480_ vssd1 vssd1 vccd1
+ vccd1 _02772_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout157_X net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08456_ net1360 top.cb_syn.char_path_n\[120\] net229 vssd1 vssd1 vccd1 vccd1 _01638_
+ sky130_fd_sc_hd__mux2_1
X_05668_ _02743_ _02744_ vssd1 vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__or2_1
X_07407_ top.dut.bit_buf\[13\] top.dut.bit_buf\[6\] net720 vssd1 vssd1 vccd1 vccd1
+ _04007_ sky130_fd_sc_hd__mux2_1
X_08387_ _02504_ _04736_ _04739_ vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__or3_1
XANTENNA__07880__A1 top.findLeastValue.sum\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout703_A net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07338_ _03733_ _03734_ _03954_ vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_21_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05599_ top.cb_syn.char_path\[77\] net551 net542 top.cb_syn.char_path\[45\] vssd1
+ vssd1 vccd1 vccd1 _02687_ sky130_fd_sc_hd__a22o_1
XANTENNA__09082__B1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_75_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07269_ net268 _03900_ _03909_ net273 net1593 vssd1 vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__a32o_1
XANTENNA__05643__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10280_ net725 net565 vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__and2_1
X_09008_ top.WB.CPU_DAT_O\[17\] net1391 net317 vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__mux2_1
Xfanout540 top.cb_syn.curr_state\[1\] vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09137__A1 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout551 net555 vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__clkbuf_4
Xfanout562 top.sram_interface.word_cnt\[0\] vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__clkbuf_2
Xfanout584 net585 vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_13_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_05_889 vssd1 vssd1 vccd1 vccd1 team_05_889/HI gpio_out[4] sky130_fd_sc_hd__conb_1
Xfanout573 net574 vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__clkbuf_2
Xfanout595 net596 vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__clkbuf_2
XFILLER_92_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_53_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_28_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11803_ clknet_leaf_92_clk _02320_ _01158_ vssd1 vssd1 vccd1 vccd1 top.compVal\[35\]
+ sky130_fd_sc_hd__dfrtp_2
X_11734_ clknet_leaf_49_clk _02267_ _01089_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.CB_write_counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05477__A3 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11665_ clknet_leaf_45_clk _02198_ _01020_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[23\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_4_6_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_6_0_clk sky130_fd_sc_hd__clkbuf_8
X_10616_ net862 net702 vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__and2_1
X_11596_ clknet_leaf_43_clk _02144_ _00951_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10547_ net833 net673 vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__and2_1
X_10478_ net856 net696 vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__and2_1
XANTENNA__05686__X _02760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06640_ _03425_ _03426_ _03428_ vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_86_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_44_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_clk sky130_fd_sc_hd__clkbuf_8
X_06571_ _02445_ top.findLeastValue.val1\[4\] top.findLeastValue.val1\[3\] _02446_
+ vssd1 vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__a22o_1
X_09290_ _04015_ _05232_ vssd1 vssd1 vccd1 vccd1 top.dut.bit_buf_next\[6\] sky130_fd_sc_hd__and2_1
X_05522_ top.cb_syn.char_path\[26\] net559 net314 top.cb_syn.char_path\[122\] vssd1
+ vssd1 vccd1 vccd1 _02623_ sky130_fd_sc_hd__a22o_1
XANTENNA__08384__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08310_ top.cb_syn.char_path_n\[14\] net195 _04682_ vssd1 vssd1 vccd1 vccd1 _01660_
+ sky130_fd_sc_hd__o21a_1
X_05453_ net555 net546 vssd1 vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__nor2_1
X_08241_ top.cb_syn.char_path_n\[49\] net376 net336 top.cb_syn.char_path_n\[47\] net181
+ vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__a221o_1
XFILLER_119_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_08172_ top.cb_syn.char_path_n\[83\] net202 _04613_ vssd1 vssd1 vccd1 vccd1 _01729_
+ sky130_fd_sc_hd__o21a_1
X_05384_ top.findLeastValue.val2\[20\] vssd1 vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__inv_2
XFILLER_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08811__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07123_ _03723_ _03780_ _03726_ _03724_ vssd1 vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__o211a_1
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 WE_O sky130_fd_sc_hd__buf_2
X_07054_ top.findLeastValue.val1\[14\] top.findLeastValue.val2\[14\] vssd1 vssd1 vccd1
+ vccd1 _03712_ sky130_fd_sc_hd__nand2_1
XANTENNA__05625__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06005_ net1498 top.WB.CPU_DAT_O\[30\] net357 vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__mux2_1
XANTENNA__07378__B1 _03553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07029__A top.findLeastValue.val1\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06050__B1 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07956_ top.findLeastValue.least1\[1\] top.findLeastValue.least2\[1\] _04462_ vssd1
+ vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__mux2_1
X_06907_ top.findLeastValue.val2\[30\] net148 net121 _03595_ vssd1 vssd1 vccd1 vccd1
+ _01972_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_106_Right_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout274_X net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout653_A net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07887_ net425 _04414_ _04415_ net259 vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__o211a_1
XFILLER_102_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06838_ _02474_ net152 net126 _03558_ vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_16_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_26_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09626_ net759 net599 vssd1 vssd1 vccd1 vccd1 _00240_ sky130_fd_sc_hd__and2_1
X_06769_ net502 net412 net119 net134 top.cw1\[2\] vssd1 vssd1 vccd1 vccd1 _02067_
+ sky130_fd_sc_hd__a32o_1
X_09557_ net795 net635 vssd1 vssd1 vccd1 vccd1 _00171_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_54_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout441_X net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout820_A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_35_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07699__A net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08508_ net1090 top.cb_syn.char_path_n\[68\] net227 vssd1 vssd1 vccd1 vccd1 _01586_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09488_ net732 net572 vssd1 vssd1 vccd1 vccd1 _00102_ sky130_fd_sc_hd__and2_1
X_08439_ _02503_ _04789_ _04791_ _04792_ _04797_ vssd1 vssd1 vccd1 vccd1 _04798_ sky130_fd_sc_hd__o32a_1
XFILLER_24_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout706_X net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07853__A1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11450_ clknet_leaf_71_clk _01998_ _00805_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least2\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_12_Left_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11381_ clknet_leaf_86_clk _01929_ _00736_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[33\]
+ sky130_fd_sc_hd__dfrtp_1
X_10401_ net767 net607 vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__and2_1
XANTENNA__06408__A2 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10332_ net795 net635 vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__and2_1
XANTENNA__05616__B1 _02700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10263_ net873 net713 vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__and2_1
XFILLER_78_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11457__Q top.findLeastValue.least2\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10194_ net863 net703 vssd1 vssd1 vccd1 vccd1 _00808_ sky130_fd_sc_hd__and2_1
XANTENNA__09154__A net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout370 _05086_ vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__buf_2
Xfanout392 net393 vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout381 net382 vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Left_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06895__A2 net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09601__B net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_26_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07519__S1 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11717_ clknet_leaf_122_clk _02250_ _01072_ vssd1 vssd1 vccd1 vccd1 top.path\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_30_Left_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05855__B1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput12 DAT_I[19] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
X_11648_ clknet_leaf_113_clk _02181_ _01003_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput34 en vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_2
Xinput23 DAT_I[29] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
X_11579_ clknet_leaf_108_clk _02127_ _00934_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05607__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11367__Q top.findLeastValue.sum\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07375__A3 _03547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07810_ top.findLeastValue.sum\[26\] _04353_ net395 vssd1 vssd1 vccd1 vccd1 _04354_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08790_ net437 _04942_ _04944_ _04945_ net520 vssd1 vssd1 vccd1 vccd1 _04973_ sky130_fd_sc_hd__a221o_1
XFILLER_111_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07741_ net488 _04297_ vssd1 vssd1 vccd1 vccd1 _04299_ sky130_fd_sc_hd__or2_1
X_07672_ _04241_ _04242_ net486 vssd1 vssd1 vccd1 vccd1 _04243_ sky130_fd_sc_hd__mux2_1
XFILLER_37_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09411_ net1001 net241 _05283_ _05284_ vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__a22o_1
X_06623_ top.compVal\[44\] _02460_ _03391_ _03403_ vssd1 vssd1 vccd1 vccd1 _03412_
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_17_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_8
X_06554_ _02427_ top.findLeastValue.val1\[22\] top.findLeastValue.val1\[21\] _02428_
+ vssd1 vssd1 vccd1 vccd1 _03343_ sky130_fd_sc_hd__a22o_1
X_09342_ net1053 net236 net214 _04418_ vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__a22o_1
X_05505_ _02607_ _02608_ net474 vssd1 vssd1 vccd1 vccd1 _02609_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_51_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09273_ _05224_ vssd1 vssd1 vccd1 vccd1 _05225_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout234_A net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06485_ net1487 _03288_ vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__xor2_1
XANTENNA__11830__Q top.WB.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05436_ top.WB.curr_state\[2\] top.WB.curr_state\[1\] vssd1 vssd1 vccd1 vccd1 _02544_
+ sky130_fd_sc_hd__nor2_1
X_08224_ top.cb_syn.char_path_n\[57\] net205 _04639_ vssd1 vssd1 vccd1 vccd1 _01703_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__05846__B1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout401_A net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08155_ top.cb_syn.char_path_n\[92\] net389 net348 top.cb_syn.char_path_n\[90\] net193
+ vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__a221o_1
X_05367_ top.findLeastValue.least2\[5\] vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__inv_2
XFILLER_119_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07106_ top.findLeastValue.val1\[4\] top.findLeastValue.val2\[4\] _03743_ _03742_
+ vssd1 vssd1 vccd1 vccd1 _03764_ sky130_fd_sc_hd__a31o_1
XANTENNA__05767__A net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08086_ top.cb_syn.char_path_n\[126\] net207 _04570_ vssd1 vssd1 vccd1 vccd1 _01772_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__06362__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05298_ top.compVal\[45\] vssd1 vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__inv_2
XANTENNA__06271__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06810__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07037_ _03689_ _03693_ vssd1 vssd1 vccd1 vccd1 _03695_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout391_X net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout868_A net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08988_ top.WB.CPU_DAT_O\[4\] net1410 net323 vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__mux2_1
X_07939_ top.findLeastValue.sum\[0\] top.hTree.tree_reg\[0\] net284 vssd1 vssd1 vccd1
+ vccd1 _04457_ sky130_fd_sc_hd__mux2_1
X_10950_ clknet_leaf_36_clk _01505_ _00305_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.num_lefts\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_90_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07206__B _03657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_09609_ net844 net684 vssd1 vssd1 vccd1 vccd1 _00223_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout823_X net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10881_ clknet_leaf_110_clk _01458_ _00236_ vssd1 vssd1 vccd1 vccd1 top.translation.totalEn
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__06877__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11502_ clknet_leaf_90_clk _02050_ _00857_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[42\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__05837__B1 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11433_ clknet_leaf_91_clk _01981_ _00788_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[39\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_59_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08053__A net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11364_ clknet_leaf_106_clk _01912_ _00719_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08251__B2 top.cb_syn.char_path_n\[42\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11295_ clknet_leaf_83_clk _01843_ _00650_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06801__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10315_ net764 net604 vssd1 vssd1 vccd1 vccd1 _00929_ sky130_fd_sc_hd__and2_1
XFILLER_98_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10246_ net842 net682 vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__and2_1
XFILLER_105_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10177_ net836 net676 vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__and2_1
XANTENNA__08927__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10477__B net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05540__A2 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06270_ _02574_ _02992_ _03135_ vssd1 vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__and3_1
XANTENNA__09019__A0 top.WB.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08778__C1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold615 top.cb_syn.state8 vssd1 vssd1 vccd1 vccd1 net1568 sky130_fd_sc_hd__dlygate4sd3_1
Xhold604 top.histogram.state\[6\] vssd1 vssd1 vccd1 vccd1 net1557 sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 top.hTree.tree_reg\[7\] vssd1 vssd1 vccd1 vccd1 net1579 sky130_fd_sc_hd__dlygate4sd3_1
Xhold659 top.cw1\[5\] vssd1 vssd1 vccd1 vccd1 net1612 sky130_fd_sc_hd__dlygate4sd3_1
Xhold637 _00013_ vssd1 vssd1 vccd1 vccd1 net1590 sky130_fd_sc_hd__dlygate4sd3_1
X_09960_ net771 net611 vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_6_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_8
Xhold648 top.histogram.total\[12\] vssd1 vssd1 vccd1 vccd1 net1601 sky130_fd_sc_hd__dlygate4sd3_1
X_08911_ top.cb_syn.max_index\[3\] top.cb_syn.max_index\[2\] top.cb_syn.max_index\[1\]
+ top.cb_syn.max_index\[4\] vssd1 vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__a31o_1
XANTENNA__06910__S net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09891_ net773 net613 vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__and2_1
XFILLER_69_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07753__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08842_ top.path\[40\] net410 net328 top.path\[41\] net437 vssd1 vssd1 vccd1 vccd1
+ _05025_ sky130_fd_sc_hd__o221a_1
XFILLER_111_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05985_ _02915_ _02917_ vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__nor2_1
XANTENNA__11825__Q top.WB.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08773_ net521 _04949_ _04948_ _02522_ vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout184_A net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07724_ top.findLeastValue.sum\[43\] top.hTree.tree_reg\[43\] net283 vssd1 vssd1
+ vccd1 vccd1 _04285_ sky130_fd_sc_hd__mux2_1
XFILLER_38_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07655_ top.hTree.tree_reg\[56\] net397 net286 vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout351_A net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06606_ _02410_ top.findLeastValue.val1\[39\] vssd1 vssd1 vccd1 vccd1 _03395_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_36_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07586_ top.cb_syn.max_index\[2\] top.cb_syn.max_index\[1\] top.cb_syn.max_index\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04173_ sky130_fd_sc_hd__o21ai_1
XFILLER_80_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__05531__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06537_ top.FLV_done _02548_ _03326_ net287 net958 vssd1 vssd1 vccd1 vccd1 _02073_
+ sky130_fd_sc_hd__a32o_1
X_09325_ net36 _05258_ _05259_ vssd1 vssd1 vccd1 vccd1 top.translation.writeBin sky130_fd_sc_hd__and3_1
XANTENNA__07808__A1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09256_ _02543_ _04921_ _05200_ vssd1 vssd1 vccd1 vccd1 _05213_ sky130_fd_sc_hd__nor3_4
XANTENNA_fanout616_A net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06468_ top.histogram.total\[27\] top.histogram.total\[26\] _03290_ vssd1 vssd1 vccd1
+ vccd1 _03291_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_97_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05419_ net529 vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__inv_2
X_08207_ top.cb_syn.char_path_n\[66\] net388 net347 top.cb_syn.char_path_n\[64\] net191
+ vssd1 vssd1 vccd1 vccd1 _04631_ sky130_fd_sc_hd__a221o_1
X_09187_ net1686 _02541_ _02593_ vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__a21o_1
X_06399_ net1114 _03236_ net300 vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__mux2_1
X_08138_ top.cb_syn.char_path_n\[100\] net203 _04596_ vssd1 vssd1 vccd1 vccd1 _01746_
+ sky130_fd_sc_hd__o21a_1
XFILLER_108_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_08069_ _04131_ _04478_ vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__nor2_1
X_11080_ clknet_leaf_6_clk _01628_ _00435_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[110\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05598__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10100_ net827 net667 vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__and2_1
X_10031_ net839 net679 vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__and2_1
XFILLER_102_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10933_ clknet_leaf_32_clk _01488_ _00288_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.zeroes\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_106_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05507__C1 _02610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05522__A2 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10864_ clknet_leaf_79_clk _01450_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[56\]
+ sky130_fd_sc_hd__dfxtp_1
X_10795_ clknet_leaf_52_clk net1473 _00214_ vssd1 vssd1 vccd1 vccd1 top.histogram.state\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08482__S net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11416_ clknet_leaf_103_clk _01964_ _00771_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[22\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_117_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11347_ clknet_leaf_59_clk net1695 _00702_ vssd1 vssd1 vccd1 vccd1 top.cw2\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_4_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08775__A2 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11278_ clknet_leaf_77_clk _01826_ _00633_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09326__B net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10229_ net827 net667 vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__and2_1
Xhold1 top.controller.fin_FINISHED vssd1 vssd1 vccd1 vccd1 net954 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_67_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05770_ top.translation.index\[6\] top.translation.index\[5\] _02789_ vssd1 vssd1
+ vccd1 vccd1 _02791_ sky130_fd_sc_hd__or3_1
X_07440_ _04030_ _04034_ net404 vssd1 vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__mux2_1
XANTENNA__05513__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07502__A3 top.cb_syn.char_path_n\[41\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07371_ top.findLeastValue.histo_index\[3\] _03553_ _03978_ vssd1 vssd1 vccd1 vccd1
+ _03979_ sky130_fd_sc_hd__a21o_1
X_09110_ net447 _02820_ _05127_ net455 _05128_ vssd1 vssd1 vccd1 vccd1 _05129_ sky130_fd_sc_hd__o221a_1
X_06322_ top.hist_data_o\[16\] top.hist_data_o\[15\] top.hist_data_o\[14\] _03184_
+ vssd1 vssd1 vccd1 vccd1 _03185_ sky130_fd_sc_hd__and4_1
X_09041_ net1229 top.WB.CPU_DAT_O\[16\] net291 vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__mux2_1
X_06253_ _02912_ _02942_ _02944_ _03021_ _03119_ vssd1 vssd1 vccd1 vccd1 _03120_ sky130_fd_sc_hd__a32o_1
Xhold401 net88 vssd1 vssd1 vccd1 vccd1 net1354 sky130_fd_sc_hd__dlygate4sd3_1
X_06184_ top.TRN_char_index\[4\] _02975_ vssd1 vssd1 vccd1 vccd1 _03054_ sky130_fd_sc_hd__nor2_1
Xhold445 net64 vssd1 vssd1 vccd1 vccd1 net1398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold412 top.path\[45\] vssd1 vssd1 vccd1 vccd1 net1365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 top.path\[59\] vssd1 vssd1 vccd1 vccd1 net1376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 top.hTree.tree_reg\[3\] vssd1 vssd1 vccd1 vccd1 net1387 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold467 top.histogram.sram_out\[30\] vssd1 vssd1 vccd1 vccd1 net1420 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06777__B2 top.findLeastValue.histo_index\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold456 _01836_ vssd1 vssd1 vccd1 vccd1 net1409 sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 top.histogram.sram_out\[7\] vssd1 vssd1 vccd1 vccd1 net1431 sky130_fd_sc_hd__dlygate4sd3_1
X_09943_ net744 net584 vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__and2_1
Xhold489 top.cb_syn.char_path\[76\] vssd1 vssd1 vccd1 vccd1 net1442 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09874_ net788 net628 vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout399_A net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08825_ top.path\[8\] net410 net328 top.path\[9\] net437 vssd1 vssd1 vccd1 vccd1
+ _05008_ sky130_fd_sc_hd__o221a_1
X_05968_ top.sram_interface.init_counter\[1\] _02903_ vssd1 vssd1 vccd1 vccd1 _02904_
+ sky130_fd_sc_hd__and2_1
X_08756_ net434 _04937_ _04938_ vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__o21a_1
X_08687_ _04875_ _04882_ vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__nor2_1
X_05899_ net536 _02868_ _02873_ vssd1 vssd1 vccd1 vccd1 _02874_ sky130_fd_sc_hd__a21o_1
X_07707_ net490 _04271_ vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout733_A net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05504__A2 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07638_ top.findLeastValue.least1\[4\] top.hTree.tree_reg\[59\] net279 vssd1 vssd1
+ vccd1 vccd1 _04215_ sky130_fd_sc_hd__mux2_1
XFILLER_14_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07569_ top.cb_syn.max_index\[6\] _04136_ _04155_ _04158_ vssd1 vssd1 vccd1 vccd1
+ _04159_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout521_X net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09398__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09308_ top.histogram.total\[8\] net409 net327 top.histogram.total\[9\] net436 vssd1
+ vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_101_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10580_ net746 net586 vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_11_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09239_ net296 _05204_ vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_header\[0\]
+ sky130_fd_sc_hd__and2_1
XFILLER_119_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10634__Q top.sram_interface.word_cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11201_ clknet_leaf_9_clk _01749_ _00556_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[103\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06768__A1 top.findLeastValue.histo_index\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11132_ clknet_leaf_17_clk _01680_ _00487_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[34\]
+ sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11063_ clknet_leaf_42_clk _01611_ _00418_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[93\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10014_ net819 net659 vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__and2_1
XFILLER_63_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06153__C1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10916_ clknet_leaf_75_clk _01472_ _00271_ vssd1 vssd1 vccd1 vccd1 top.hTree.finish_check
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10847_ clknet_leaf_106_clk _01433_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_4_Left_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10778_ clknet_leaf_45_clk _01377_ _00197_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08940__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06940_ top.compVal\[13\] top.findLeastValue.val1\[13\] net162 vssd1 vssd1 vccd1
+ vccd1 _03612_ sky130_fd_sc_hd__mux2_1
X_06871_ _03012_ _03110_ _03576_ _03567_ top.findLeastValue.histo_index\[3\] vssd1
+ vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__a32o_1
X_08610_ top.cb_syn.num_lefts\[3\] top.cb_syn.num_lefts\[2\] top.cb_syn.num_lefts\[1\]
+ top.cb_syn.num_lefts\[0\] vssd1 vssd1 vccd1 vccd1 _04829_ sky130_fd_sc_hd__and4_1
X_05822_ net556 _02835_ net546 net454 vssd1 vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__a2bb2o_1
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09590_ net844 net684 vssd1 vssd1 vccd1 vccd1 _00204_ sky130_fd_sc_hd__and2_1
X_08541_ net1225 top.cb_syn.char_path_n\[35\] net228 vssd1 vssd1 vccd1 vccd1 _01553_
+ sky130_fd_sc_hd__mux2_1
X_05753_ top.compVal\[41\] net172 net158 top.WB.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1
+ _02326_ sky130_fd_sc_hd__a22o_1
X_05684_ top.WB.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__and2_1
XANTENNA__08133__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08472_ net1379 top.cb_syn.char_path_n\[104\] net225 vssd1 vssd1 vccd1 vccd1 _01622_
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07423_ _03993_ _04020_ _03986_ vssd1 vssd1 vccd1 vccd1 _04021_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_59_Left_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08436__B2 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07354_ _03747_ _03758_ _03757_ vssd1 vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__a21o_1
XFILLER_109_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout314_A net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06305_ _03168_ _03165_ _03164_ vssd1 vssd1 vccd1 vccd1 _03169_ sky130_fd_sc_hd__or3b_1
X_07285_ _03782_ _03799_ vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__or2_1
X_06236_ top.TRN_char_index\[0\] _03102_ _03103_ net464 vssd1 vssd1 vccd1 vccd1 _03104_
+ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09024_ top.WB.CPU_DAT_O\[1\] net1145 net320 vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__mux2_1
XANTENNA__05670__A1 top.histogram.sram_out\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold220 top.path\[62\] vssd1 vssd1 vccd1 vccd1 net1173 sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 top.header_synthesis.header\[4\] vssd1 vssd1 vccd1 vccd1 net1206 sky130_fd_sc_hd__dlygate4sd3_1
X_06167_ net471 _03018_ _03037_ vssd1 vssd1 vccd1 vccd1 _03038_ sky130_fd_sc_hd__a21bo_1
Xhold242 top.hTree.nulls\[61\] vssd1 vssd1 vccd1 vccd1 net1195 sky130_fd_sc_hd__dlygate4sd3_1
Xhold231 top.hTree.tree_reg\[57\] vssd1 vssd1 vccd1 vccd1 net1184 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06098_ top.TRN_char_index\[3\] top.TRN_char_index\[2\] top.TRN_char_index\[1\] vssd1
+ vssd1 vccd1 vccd1 _02971_ sky130_fd_sc_hd__and3_1
Xfanout700 net717 vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout683_A net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold264 top.cb_syn.char_path\[21\] vssd1 vssd1 vccd1 vccd1 net1217 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_68_Left_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold286 top.histogram.sram_out\[19\] vssd1 vssd1 vccd1 vccd1 net1239 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold275 top.path\[24\] vssd1 vssd1 vccd1 vccd1 net1228 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout722 net37 vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__buf_4
Xfanout711 net712 vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__clkbuf_2
X_09926_ net790 net630 vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__and2_1
Xhold297 top.path\[39\] vssd1 vssd1 vccd1 vccd1 net1250 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout733 net734 vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__clkbuf_2
Xfanout766 net767 vssd1 vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__clkbuf_2
Xfanout744 net745 vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__clkbuf_2
Xfanout755 net756 vssd1 vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__clkbuf_2
Xfanout799 net800 vssd1 vssd1 vccd1 vccd1 net799 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout850_A net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout777 net779 vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__clkbuf_2
Xfanout788 net791 vssd1 vssd1 vccd1 vccd1 net788 sky130_fd_sc_hd__clkbuf_2
X_09857_ net772 net612 vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__and2_1
X_08808_ top.path\[61\] net326 _04990_ vssd1 vssd1 vccd1 vccd1 _04991_ sky130_fd_sc_hd__o21a_1
X_09788_ net741 net581 vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__and2_1
X_08739_ _03245_ _04921_ vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_77_Left_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ clknet_leaf_95_clk _02283_ _01105_ vssd1 vssd1 vccd1 vccd1 top.compVal\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05489__A1 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10701_ clknet_leaf_11_clk _01300_ _00120_ vssd1 vssd1 vccd1 vccd1 top.path\[77\]
+ sky130_fd_sc_hd__dfrtp_1
X_11681_ clknet_leaf_61_clk _02214_ _01036_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10632_ net857 net697 vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_62_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10563_ net814 net654 vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__and2_1
XFILLER_10_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08045__B net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_10494_ net825 net665 vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__and2_1
XANTENNA__08760__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11115_ clknet_leaf_22_clk _01663_ _00470_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[17\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_96_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11046_ clknet_leaf_4_clk _01594_ _00401_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[76\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_103_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08902__A2 _04188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05716__A2 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09312__C1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11879_ clknet_leaf_70_clk _02395_ _01234_ vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__dfrtp_1
XFILLER_44_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07070_ top.findLeastValue.val1\[10\] top.findLeastValue.val2\[10\] vssd1 vssd1 vccd1
+ vccd1 _03728_ sky130_fd_sc_hd__or2_1
X_06021_ net1715 top.WB.CPU_DAT_O\[14\] net356 vssd1 vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__mux2_1
XFILLER_99_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07929__A0 top.findLeastValue.sum\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09217__D top.controller.fin_reg\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09711_ net789 net629 vssd1 vssd1 vccd1 vccd1 _00325_ sky130_fd_sc_hd__and2_1
X_07972_ top.findLeastValue.alternator_timer\[0\] _03565_ _04477_ _03326_ vssd1 vssd1
+ vccd1 vccd1 _01793_ sky130_fd_sc_hd__a22o_1
XANTENNA__08354__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06923_ top.findLeastValue.val2\[22\] net146 net120 _03603_ vssd1 vssd1 vccd1 vccd1
+ _01964_ sky130_fd_sc_hd__o22a_1
X_09642_ net804 net644 vssd1 vssd1 vccd1 vccd1 _00256_ sky130_fd_sc_hd__and2_1
X_06854_ top.findLeastValue.startup net470 net288 vssd1 vssd1 vccd1 vccd1 _03568_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__06904__A1 top.findLeastValue.val1\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09573_ net796 net636 vssd1 vssd1 vccd1 vccd1 _00187_ sky130_fd_sc_hd__and2_1
X_05805_ _02816_ _02824_ vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__and2_1
XANTENNA__11833__Q top.WB.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06785_ top.findLeastValue.val1\[45\] net133 net117 top.compVal\[45\] vssd1 vssd1
+ vccd1 vccd1 _02053_ sky130_fd_sc_hd__o22a_1
X_05736_ _02769_ _02770_ _02765_ vssd1 vssd1 vccd1 vccd1 _02771_ sky130_fd_sc_hd__o21ba_1
XANTENNA_fanout264_A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08524_ net1417 top.cb_syn.char_path_n\[52\] net222 vssd1 vssd1 vccd1 vccd1 _01570_
+ sky130_fd_sc_hd__mux2_1
X_08455_ net1375 top.cb_syn.char_path_n\[121\] net231 vssd1 vssd1 vccd1 vccd1 _01639_
+ sky130_fd_sc_hd__mux2_1
X_05667_ top.cb_syn.char_path\[2\] net558 net316 top.cb_syn.char_path\[98\] vssd1
+ vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout431_A _02530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07406_ top.dut.bits_in_buf\[1\] top.dut.bits_in_buf\[2\] net404 vssd1 vssd1 vccd1
+ vccd1 _04006_ sky130_fd_sc_hd__and3_1
XANTENNA__08409__B2 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08386_ top.cb_syn.char_path_n\[97\] net391 _04744_ vssd1 vssd1 vccd1 vccd1 _04745_
+ sky130_fd_sc_hd__a21oi_1
X_05598_ net1270 net138 _02686_ net174 vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__a22o_1
XFILLER_11_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_07337_ net270 _03956_ _03959_ net275 net1685 vssd1 vssd1 vccd1 vccd1 _01906_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_21_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07268_ _03702_ _03708_ _03899_ vssd1 vssd1 vccd1 vccd1 _03909_ sky130_fd_sc_hd__nand3_1
X_06219_ net1407 _02595_ _03087_ net160 vssd1 vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__a22o_1
XFILLER_117_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06840__B1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09007_ top.WB.CPU_DAT_O\[18\] net1097 net317 vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__mux2_1
X_07199_ _03848_ _03851_ _03854_ _03856_ _03847_ vssd1 vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__o221a_1
XFILLER_104_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xfanout530 top.cb_syn.curr_state\[7\] vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__buf_2
Xfanout541 top.sram_interface.word_cnt\[12\] vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__buf_2
XANTENNA__07491__S1 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07924__S net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout552 net555 vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__buf_2
XFILLER_58_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09909_ net760 net600 vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__and2_1
Xfanout563 net567 vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__clkbuf_2
Xfanout574 net585 vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__clkbuf_2
Xfanout585 net647 vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__clkbuf_2
Xfanout596 net597 vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_85_Left_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11970__A net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ clknet_leaf_92_clk _02319_ _01157_ vssd1 vssd1 vccd1 vccd1 top.compVal\[34\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_61_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ clknet_leaf_61_clk _02266_ _01088_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.check
+ sky130_fd_sc_hd__dfrtp_1
X_11664_ clknet_leaf_16_clk _02197_ _01019_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08056__A net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10615_ net768 net608 vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_94_Left_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11595_ clknet_leaf_40_clk _02143_ _00950_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08490__S net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08820__A1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10546_ net832 net672 vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__and2_1
X_10477_ net856 net696 vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__and2_1
XFILLER_108_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__07834__S net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11029_ clknet_leaf_27_clk _01577_ _00384_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05570__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06570_ _02446_ top.findLeastValue.val1\[3\] top.findLeastValue.val1\[2\] _02447_
+ vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__o22a_1
X_05521_ top.cb_syn.char_path\[90\] net553 net544 top.cb_syn.char_path\[58\] vssd1
+ vssd1 vccd1 vccd1 _02622_ sky130_fd_sc_hd__a22o_1
XANTENNA__07847__C1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05452_ net463 net561 vssd1 vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__nand2_1
X_08240_ top.cb_syn.char_path_n\[49\] net198 _04647_ vssd1 vssd1 vccd1 vccd1 _01695_
+ sky130_fd_sc_hd__o21a_1
X_08171_ top.cb_syn.char_path_n\[84\] net382 net341 top.cb_syn.char_path_n\[82\] net186
+ vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__a221o_1
X_07122_ _03779_ vssd1 vssd1 vccd1 vccd1 _03780_ sky130_fd_sc_hd__inv_2
X_05383_ top.findLeastValue.val2\[21\] vssd1 vssd1 vccd1 vccd1 _02491_ sky130_fd_sc_hd__inv_2
Xoutput100 net100 vssd1 vssd1 vccd1 vccd1 DAT_O[5] sky130_fd_sc_hd__buf_2
X_07053_ _03709_ _03710_ vssd1 vssd1 vccd1 vccd1 _03711_ sky130_fd_sc_hd__and2b_1
X_06004_ net1491 top.WB.CPU_DAT_O\[31\] net357 vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__mux2_1
Xoutput111 net111 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
XANTENNA__11828__Q top.WB.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07029__B top.findLeastValue.val2\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07955_ net1456 _04467_ _04461_ vssd1 vssd1 vccd1 vccd1 _01800_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout381_A net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07744__S net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout479_A net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06906_ top.compVal\[30\] top.findLeastValue.val1\[30\] net163 vssd1 vssd1 vccd1
+ vccd1 _03595_ sky130_fd_sc_hd__mux2_1
X_09625_ net844 net684 vssd1 vssd1 vccd1 vccd1 _00239_ sky130_fd_sc_hd__and2_1
XANTENNA__08422__S0 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07886_ net482 _04413_ vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout646_A net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout267_X net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06837_ top.findLeastValue.least1\[6\] net497 _03424_ vssd1 vssd1 vccd1 vccd1 _03558_
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06768_ top.findLeastValue.histo_index\[3\] net412 net119 net135 net1561 vssd1 vssd1
+ vccd1 vccd1 _02068_ sky130_fd_sc_hd__a32o_1
XANTENNA__08575__S net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09556_ net733 net573 vssd1 vssd1 vccd1 vccd1 _00170_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_54_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08507_ net1125 top.cb_syn.char_path_n\[69\] net227 vssd1 vssd1 vccd1 vccd1 _01587_
+ sky130_fd_sc_hd__mux2_1
X_05719_ net13 net418 net360 top.WB.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1 _02339_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout434_X net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06699_ top.compVal\[20\] _02492_ top.findLeastValue.val2\[16\] _02433_ vssd1 vssd1
+ vccd1 vccd1 _03487_ sky130_fd_sc_hd__a22o_1
X_09487_ net729 net569 vssd1 vssd1 vccd1 vccd1 _00101_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout813_A net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08438_ _02504_ _04794_ _04796_ top.cb_syn.end_cnt\[4\] vssd1 vssd1 vccd1 vccd1 _04797_
+ sky130_fd_sc_hd__a31o_1
XFILLER_11_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08369_ _02506_ top.cb_syn.char_path_n\[120\] _04727_ net511 vssd1 vssd1 vccd1 vccd1
+ _04728_ sky130_fd_sc_hd__o211a_1
XANTENNA__09055__A1 top.WB.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05864__B2 top.WB.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11380_ clknet_leaf_86_clk _01928_ _00735_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[32\]
+ sky130_fd_sc_hd__dfrtp_1
X_10400_ net766 net606 vssd1 vssd1 vccd1 vccd1 _01014_ sky130_fd_sc_hd__and2_1
XANTENNA__07919__S net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10331_ net793 net633 vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__and2_1
XANTENNA__06813__B1 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10262_ net872 net712 vssd1 vssd1 vccd1 vccd1 _00876_ sky130_fd_sc_hd__and2_1
XFILLER_3_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09358__A2 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10193_ net863 net703 vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__and2_1
XANTENNA__05963__A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09154__B net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout371 net372 vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__clkbuf_4
Xfanout393 _04539_ vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__buf_2
Xfanout360 _02761_ vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout382 net390 vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__buf_2
XFILLER_19_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_109_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05552__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_11716_ clknet_leaf_121_clk _02249_ _01071_ vssd1 vssd1 vccd1 vccd1 top.path\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__05855__B2 top.WB.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09046__A1 top.WB.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput13 DAT_I[1] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
X_11647_ clknet_leaf_113_clk _02180_ _01002_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput35 gpio_in[10] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__buf_1
XANTENNA__07829__S net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput24 DAT_I[2] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
X_11578_ clknet_leaf_109_clk _02126_ _00933_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10529_ net848 net688 vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__and2_1
XANTENNA__06804__B1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08006__C1 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05873__A _02760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06032__A1 top.WB.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07740_ top.findLeastValue.sum\[40\] _04297_ net398 vssd1 vssd1 vccd1 vccd1 _04298_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__08309__B1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_74_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07671_ top.findLeastValue.least2\[7\] _04241_ net395 vssd1 vssd1 vccd1 vccd1 _04242_
+ sky130_fd_sc_hd__mux2_1
X_09410_ top.hTree.nulls\[57\] net406 net245 vssd1 vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__o21a_1
XANTENNA__05543__B1 _02639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06622_ _03401_ _03399_ _03396_ _03400_ vssd1 vssd1 vccd1 vccd1 _03411_ sky130_fd_sc_hd__and4b_1
XFILLER_80_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06553_ _02426_ top.findLeastValue.val1\[23\] vssd1 vssd1 vccd1 vccd1 _03342_ sky130_fd_sc_hd__and2_1
X_09341_ net995 net236 net214 _04422_ vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__a22o_1
X_05504_ top.cb_syn.char_path\[29\] net559 net314 top.cb_syn.char_path\[125\] vssd1
+ vssd1 vccd1 vccd1 _02608_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_51_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_89_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09272_ _02533_ _05222_ vssd1 vssd1 vccd1 vccd1 _05224_ sky130_fd_sc_hd__nor2_1
XFILLER_60_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06484_ _03289_ _03299_ vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__nor2_1
X_05435_ top.header_synthesis.write_zeroes vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__inv_2
X_08223_ top.cb_syn.char_path_n\[58\] net384 net342 top.cb_syn.char_path_n\[56\] net188
+ vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__a221o_1
XANTENNA__09037__A1 top.WB.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05846__B2 top.WB.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08154_ top.cb_syn.char_path_n\[92\] net208 _04604_ vssd1 vssd1 vccd1 vccd1 _01738_
+ sky130_fd_sc_hd__o21a_1
X_05366_ top.findLeastValue.least2\[6\] vssd1 vssd1 vccd1 vccd1 _02474_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout227_A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_12_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07739__S net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08085_ top.cb_syn.char_path_n\[127\] net386 net345 top.cb_syn.char_path_n\[125\]
+ net190 vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__a221o_1
XANTENNA__08424__A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07105_ _03744_ _03762_ vssd1 vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__and2_1
XANTENNA__05767__B net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05297_ net722 vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__inv_2
XANTENNA__06271__A1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07036_ _03693_ vssd1 vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout596_A net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_27_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06023__A1 top.WB.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_5_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_5_0_clk sky130_fd_sc_hd__clkbuf_8
X_08987_ top.WB.CPU_DAT_O\[5\] net1512 net323 vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout763_A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07938_ net440 net1463 net251 top.findLeastValue.sum\[1\] _04456_ vssd1 vssd1 vccd1
+ vccd1 _01806_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout551_X net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07869_ top.findLeastValue.sum\[14\] top.hTree.tree_reg\[14\] net284 vssd1 vssd1
+ vccd1 vccd1 _04401_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10880_ clknet_leaf_41_clk _00011_ _00235_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.curr_state\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_09608_ net843 net683 vssd1 vssd1 vccd1 vccd1 _00222_ sky130_fd_sc_hd__and2_1
XANTENNA__05534__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09539_ net732 net572 vssd1 vssd1 vccd1 vccd1 _00153_ sky130_fd_sc_hd__and2_1
XFILLER_12_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09028__A1 top.WB.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11501_ clknet_leaf_91_clk _02049_ _00856_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[41\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__05837__B2 top.WB.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11432_ clknet_leaf_88_clk _01980_ _00787_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[38\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_59_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11363_ clknet_leaf_98_clk _01911_ _00718_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[15\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11294_ clknet_leaf_84_clk net1544 _00649_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[37\]
+ sky130_fd_sc_hd__dfrtp_1
X_10314_ net763 net603 vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__and2_1
X_10245_ net838 net678 vssd1 vssd1 vccd1 vccd1 _00859_ sky130_fd_sc_hd__and2_1
XANTENNA__06014__A1 top.WB.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10176_ net828 net668 vssd1 vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__and2_1
XANTENNA__07762__A1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout190 net194 vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__buf_2
XFILLER_78_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload5_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05525__B1 _02624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07700__X _04266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold605 top.histogram.wr_r_en\[0\] vssd1 vssd1 vccd1 vccd1 net1558 sky130_fd_sc_hd__dlygate4sd3_1
Xhold627 top.findLeastValue.sum\[37\] vssd1 vssd1 vccd1 vccd1 net1580 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold616 top.hTree.tree_reg\[11\] vssd1 vssd1 vccd1 vccd1 net1569 sky130_fd_sc_hd__dlygate4sd3_1
Xhold649 top.FLV_done vssd1 vssd1 vccd1 vccd1 net1602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 top.hist_data_o\[12\] vssd1 vssd1 vccd1 vccd1 net1591 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_94_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08910_ top.cb_syn.max_index\[5\] _05077_ _05072_ vssd1 vssd1 vccd1 vccd1 _01391_
+ sky130_fd_sc_hd__mux2_1
X_09890_ net773 net613 vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__and2_1
XANTENNA__06005__A1 top.WB.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08841_ _02521_ _05021_ _05023_ vssd1 vssd1 vccd1 vccd1 _05024_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08950__A0 top.WB.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05984_ top.sram_interface.init_counter\[8\] _02908_ vssd1 vssd1 vccd1 vccd1 _02917_
+ sky130_fd_sc_hd__nor2_1
XFILLER_97_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_08772_ top.path\[84\] net409 _04954_ vssd1 vssd1 vccd1 vccd1 _04955_ sky130_fd_sc_hd__o21a_1
X_07723_ net440 net1537 net251 top.findLeastValue.sum\[44\] _04284_ vssd1 vssd1 vccd1
+ vccd1 _01849_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout177_A _02589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05516__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07654_ net262 _04227_ _04228_ net1184 net445 vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_36_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06605_ _02414_ top.findLeastValue.val1\[34\] vssd1 vssd1 vccd1 vccd1 _03394_ sky130_fd_sc_hd__nor2_1
X_07585_ net533 top.cb_syn.h_element\[48\] net539 top.cb_syn.h_element\[57\] _04135_
+ vssd1 vssd1 vccd1 vccd1 _04172_ sky130_fd_sc_hd__a221o_1
XFILLER_43_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11841__Q top.WB.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06536_ net424 net288 vssd1 vssd1 vccd1 vccd1 _03326_ sky130_fd_sc_hd__nor2_1
X_09324_ top.header_synthesis.bit1 top.header_synthesis.enable net431 vssd1 vssd1
+ vccd1 vccd1 _05259_ sky130_fd_sc_hd__a21o_1
X_09255_ net1185 _05212_ net296 vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_header\[8\]
+ sky130_fd_sc_hd__mux2_1
X_06467_ top.histogram.total\[25\] _03289_ vssd1 vssd1 vccd1 vccd1 _03290_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout132_X net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05418_ net539 vssd1 vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout609_A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08206_ top.cb_syn.char_path_n\[66\] net202 _04630_ vssd1 vssd1 vccd1 vccd1 _01712_
+ sky130_fd_sc_hd__o21a_1
XFILLER_21_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09186_ net1061 _02541_ _02588_ vssd1 vssd1 vccd1 vccd1 _00002_ sky130_fd_sc_hd__a21o_1
XFILLER_107_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06398_ top.hist_data_o\[6\] _03177_ vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__xor2_1
X_05349_ net530 vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__inv_2
X_08137_ top.cb_syn.char_path_n\[101\] net381 net340 top.cb_syn.char_path_n\[99\]
+ net185 vssd1 vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__a221o_1
XFILLER_107_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08068_ net538 _04554_ vssd1 vssd1 vccd1 vccd1 _04555_ sky130_fd_sc_hd__and2_1
XANTENNA__06795__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07019_ top.findLeastValue.val1\[27\] top.findLeastValue.val2\[27\] vssd1 vssd1 vccd1
+ vccd1 _03677_ sky130_fd_sc_hd__nand2_1
XFILLER_108_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10030_ net837 net677 vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__and2_1
XFILLER_76_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10932_ clknet_leaf_33_clk _01487_ _00287_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.zeroes\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_84_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10863_ clknet_leaf_46_clk _01449_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_71_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10794_ clknet_leaf_51_clk _00034_ _00213_ vssd1 vssd1 vccd1 vccd1 top.histogram.state\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08763__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08209__C1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05688__A net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11415_ clknet_leaf_101_clk _01963_ _00770_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[21\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_117_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11346_ clknet_leaf_59_clk _01894_ _00701_ vssd1 vssd1 vccd1 vccd1 top.cw2\[6\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__06786__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11277_ clknet_leaf_79_clk _01825_ _00632_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08932__A0 top.WB.CPU_DAT_O\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09326__C net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10228_ net817 net657 vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__and2_1
XFILLER_39_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xhold2 top.HT_fin_reg vssd1 vssd1 vccd1 vccd1 net955 sky130_fd_sc_hd__dlygate4sd3_1
X_10159_ net820 net660 vssd1 vssd1 vccd1 vccd1 _00773_ sky130_fd_sc_hd__and2_1
XFILLER_90_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07370_ top.cw1\[3\] net167 vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__and2_1
XANTENNA__08999__A0 top.WB.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06321_ top.hist_data_o\[13\] top.hist_data_o\[12\] _03178_ _03181_ vssd1 vssd1 vccd1
+ vccd1 _03184_ sky130_fd_sc_hd__and4_1
X_06252_ top.hist_addr\[3\] top.hist_addr\[2\] top.hist_addr\[1\] top.hist_addr\[0\]
+ net495 vssd1 vssd1 vccd1 vccd1 _03119_ sky130_fd_sc_hd__a41oi_1
XANTENNA__07671__A0 top.findLeastValue.least2\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09040_ net1178 top.WB.CPU_DAT_O\[17\] net291 vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_41_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06183_ net460 _03052_ vssd1 vssd1 vccd1 vccd1 _03053_ sky130_fd_sc_hd__nand2_1
Xhold402 top.path\[106\] vssd1 vssd1 vccd1 vccd1 net1355 sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 top.cb_syn.char_path\[116\] vssd1 vssd1 vccd1 vccd1 net1366 sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 top.histogram.total\[31\] vssd1 vssd1 vccd1 vccd1 net1388 sky130_fd_sc_hd__dlygate4sd3_1
Xhold424 top.path\[113\] vssd1 vssd1 vccd1 vccd1 net1377 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06777__A2 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold446 top.hTree.tree_reg\[19\] vssd1 vssd1 vccd1 vccd1 net1399 sky130_fd_sc_hd__dlygate4sd3_1
X_09942_ net743 net583 vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__and2_1
Xhold468 top.path\[33\] vssd1 vssd1 vccd1 vccd1 net1421 sky130_fd_sc_hd__dlygate4sd3_1
Xhold457 top.path\[100\] vssd1 vssd1 vccd1 vccd1 net1410 sky130_fd_sc_hd__dlygate4sd3_1
Xhold479 net87 vssd1 vssd1 vccd1 vccd1 net1432 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08923__A0 top.WB.CPU_DAT_O\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09873_ net788 net628 vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__and2_1
XANTENNA__11836__Q top.WB.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08824_ top.path\[10\] top.path\[11\] net528 vssd1 vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__mux2_1
XFILLER_85_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08755_ top.path\[104\] net411 net329 top.path\[105\] net437 vssd1 vssd1 vccd1 vccd1
+ _04938_ sky130_fd_sc_hd__o221a_1
X_05967_ top.sram_interface.init_counter\[0\] _02581_ _02760_ _02851_ vssd1 vssd1
+ vccd1 vccd1 _02903_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout461_A net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout559_A net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07706_ _02479_ net396 _04270_ vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__o21a_1
X_08686_ top.cb_syn.zeroes\[7\] _04884_ _04885_ _04886_ vssd1 vssd1 vccd1 vccd1 _01488_
+ sky130_fd_sc_hd__a22o_1
X_05898_ top.cb_syn.end_check top.cb_syn.curr_state\[5\] vssd1 vssd1 vccd1 vccd1 _02873_
+ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_49_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07637_ top.hTree.tree_reg\[59\] net394 net286 vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__and3_1
X_07568_ net537 _04154_ _04157_ net531 vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__a22o_1
X_09307_ net433 _05241_ vssd1 vssd1 vccd1 vccd1 _05242_ sky130_fd_sc_hd__or2_1
X_06519_ _03275_ _03313_ vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_101_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07499_ _04086_ _04087_ _04088_ _04089_ _04072_ _04071_ vssd1 vssd1 vccd1 vccd1 _04090_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout514_X net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07662__A0 top.findLeastValue.least1\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_09238_ top.header_synthesis.header\[0\] top.cb_syn.char_index\[0\] net518 vssd1
+ vssd1 vccd1 vccd1 _05204_ sky130_fd_sc_hd__mux2_1
X_09169_ net449 net1557 _02581_ _05109_ vssd1 vssd1 vccd1 vccd1 _00034_ sky130_fd_sc_hd__a211o_1
XANTENNA__08206__A2 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11200_ clknet_leaf_9_clk _01748_ _00555_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[102\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_119_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_107_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_102_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_11131_ clknet_leaf_17_clk _01679_ _00486_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[33\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_95_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11062_ clknet_leaf_27_clk _01610_ _00417_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[92\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10013_ net822 net662 vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__and2_1
XANTENNA__11973__A top.translation.writeBin vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09443__A net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input22_A DAT_I[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10915_ clknet_leaf_33_clk top.header_synthesis.next_write_zeroes _00270_ vssd1 vssd1
+ vccd1 vccd1 top.header_synthesis.write_zeroes sky130_fd_sc_hd__dfrtp_2
X_10846_ clknet_leaf_107_clk _01432_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_119_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10777_ clknet_leaf_45_clk _01376_ _00196_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11329_ clknet_leaf_51_clk _01877_ _00684_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.curr_index\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_105_Left_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06870_ _03569_ _03576_ _03579_ _03567_ net500 vssd1 vssd1 vccd1 vccd1 _01993_ sky130_fd_sc_hd__a32o_1
XANTENNA__05719__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05821_ top.sram_interface.word_cnt\[8\] net546 vssd1 vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__or2_1
XFILLER_94_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08540_ net1242 top.cb_syn.char_path_n\[36\] net227 vssd1 vssd1 vccd1 vccd1 _01554_
+ sky130_fd_sc_hd__mux2_1
X_05752_ top.compVal\[42\] net172 net158 top.WB.CPU_DAT_O\[10\] vssd1 vssd1 vccd1
+ vccd1 _02327_ sky130_fd_sc_hd__a22o_1
XANTENNA__09330__B1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05683_ net1066 net145 _02757_ net177 vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__a22o_1
XANTENNA__08133__B2 top.cb_syn.char_path_n\[101\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08471_ net1374 top.cb_syn.char_path_n\[105\] net225 vssd1 vssd1 vccd1 vccd1 _01623_
+ sky130_fd_sc_hd__mux2_1
X_07422_ _04015_ _04019_ _03987_ vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__mux2_1
XANTENNA__05498__A2 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_114_Left_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08436__A2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07353_ _03762_ net272 _03969_ net277 top.findLeastValue.sum\[4\] vssd1 vssd1 vccd1
+ vccd1 _01900_ sky130_fd_sc_hd__a32o_1
X_06304_ _02482_ top.sram_interface.word_cnt\[8\] net470 net413 _03167_ vssd1 vssd1
+ vccd1 vccd1 _03168_ sky130_fd_sc_hd__a41o_1
X_07284_ _03782_ _03799_ vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__nor2_1
X_06235_ _02563_ _02970_ _03102_ _03101_ vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__a31o_1
X_09023_ top.WB.CPU_DAT_O\[2\] net1166 net320 vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__mux2_1
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold210 top.hTree.tree_reg\[55\] vssd1 vssd1 vccd1 vccd1 net1163 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05670__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout307_A _02892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold232 top.header_synthesis.header\[7\] vssd1 vssd1 vccd1 vccd1 net1185 sky130_fd_sc_hd__dlygate4sd3_1
X_06166_ _02961_ _03031_ _03036_ _03024_ vssd1 vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__o211a_1
Xhold243 top.cb_syn.char_path\[83\] vssd1 vssd1 vccd1 vccd1 net1196 sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 top.cb_syn.char_path\[70\] vssd1 vssd1 vccd1 vccd1 net1174 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06097_ top.TRN_char_index\[2\] top.TRN_char_index\[1\] vssd1 vssd1 vccd1 vccd1 _02970_
+ sky130_fd_sc_hd__nand2_1
Xhold265 top.path\[42\] vssd1 vssd1 vccd1 vccd1 net1218 sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 top.path\[16\] vssd1 vssd1 vccd1 vccd1 net1229 sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 top.path\[102\] vssd1 vssd1 vccd1 vccd1 net1240 sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 top.path\[67\] vssd1 vssd1 vccd1 vccd1 net1207 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout712 net716 vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__clkbuf_2
Xfanout701 net717 vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__buf_1
X_09925_ net776 net616 vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__and2_1
Xfanout723 net727 vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__clkbuf_2
Xhold298 top.path\[25\] vssd1 vssd1 vccd1 vccd1 net1251 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_86_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09856_ net769 net609 vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__and2_1
Xfanout745 net807 vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__clkbuf_2
Xfanout767 net807 vssd1 vssd1 vccd1 vccd1 net767 sky130_fd_sc_hd__clkbuf_2
Xfanout756 net757 vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__clkbuf_2
Xfanout734 net745 vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__clkbuf_2
XFILLER_105_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xfanout778 net779 vssd1 vssd1 vccd1 vccd1 net778 sky130_fd_sc_hd__clkbuf_2
Xfanout789 net790 vssd1 vssd1 vccd1 vccd1 net789 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08372__A1 _02505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05791__A net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08807_ top.path\[60\] net408 _04989_ net432 net521 vssd1 vssd1 vccd1 vccd1 _04990_
+ sky130_fd_sc_hd__o221a_1
XFILLER_105_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_fanout843_A net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06999_ _03646_ _03651_ _03656_ _03641_ vssd1 vssd1 vccd1 vccd1 _03657_ sky130_fd_sc_hd__a31o_1
X_09787_ net736 net576 vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__and2_1
X_08738_ _04921_ vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__inv_2
X_08669_ _02933_ _04870_ _04871_ vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout631_X net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10700_ clknet_leaf_111_clk _01299_ _00119_ vssd1 vssd1 vccd1 vccd1 top.path\[76\]
+ sky130_fd_sc_hd__dfrtp_1
X_11680_ clknet_leaf_62_clk _02213_ _01035_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10631_ net853 net693 vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_62_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10562_ net854 net694 vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__and2_1
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11968__A net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05966__A _02581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05661__A2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10493_ net825 net665 vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_114_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08060__B1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05949__A0 top.WB.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07938__B2 top.findLeastValue.sum\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11114_ clknet_leaf_7_clk _01662_ _00469_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11045_ clknet_leaf_3_clk _01593_ _00400_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[75\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input25_X net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09312__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07874__A0 top.findLeastValue.sum\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11878_ clknet_leaf_39_clk _02394_ _01233_ vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__dfrtp_1
XFILLER_32_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10829_ clknet_leaf_77_clk _01415_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07626__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06020_ net1720 top.WB.CPU_DAT_O\[15\] net356 vssd1 vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__mux2_1
XANTENNA__05652__A2 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07971_ top.findLeastValue.alternator_timer\[0\] _02771_ vssd1 vssd1 vccd1 vccd1
+ _04477_ sky130_fd_sc_hd__nor2_1
XFILLER_113_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09710_ net802 net642 vssd1 vssd1 vccd1 vccd1 _00324_ sky130_fd_sc_hd__and2_1
XFILLER_101_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06922_ top.compVal\[22\] top.findLeastValue.val1\[22\] net161 vssd1 vssd1 vccd1
+ vccd1 _03603_ sky130_fd_sc_hd__mux2_1
X_09641_ net804 net644 vssd1 vssd1 vccd1 vccd1 _00255_ sky130_fd_sc_hd__and2_1
X_06853_ _02773_ _03325_ vssd1 vssd1 vccd1 vccd1 _03567_ sky130_fd_sc_hd__and2_1
X_09572_ net796 net636 vssd1 vssd1 vccd1 vccd1 _00186_ sky130_fd_sc_hd__and2_1
X_05804_ _02796_ _02800_ _02823_ vssd1 vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__and3_1
X_06784_ top.findLeastValue.val1\[46\] net288 net117 vssd1 vssd1 vccd1 vccd1 _02054_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__10022__A net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05735_ top.findLeastValue.alternator_timer\[2\] _02764_ top.findLeastValue.alternator_timer\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02770_ sky130_fd_sc_hd__o21a_1
X_08523_ net1339 top.cb_syn.char_path_n\[53\] net230 vssd1 vssd1 vccd1 vccd1 _01571_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout257_A _04190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08454_ net1299 top.cb_syn.char_path_n\[122\] net231 vssd1 vssd1 vccd1 vccd1 _01640_
+ sky130_fd_sc_hd__mux2_1
X_05666_ top.cb_syn.char_path\[66\] net553 net545 top.cb_syn.char_path\[34\] vssd1
+ vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__a22o_1
XANTENNA__09022__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07405_ _04003_ _04004_ net404 vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__mux2_1
XANTENNA__08409__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08385_ top.cb_syn.char_path_n\[98\] net332 _04743_ net509 net508 vssd1 vssd1 vccd1
+ vccd1 _04744_ sky130_fd_sc_hd__a221o_1
X_05597_ top.histogram.sram_out\[14\] net363 _02684_ _02685_ vssd1 vssd1 vccd1 vccd1
+ _02686_ sky130_fd_sc_hd__a211o_1
XFILLER_23_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08814__C1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07336_ _03729_ _03955_ vssd1 vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_21_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07267_ net268 _03907_ _03908_ net273 net1640 vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__a32o_1
X_09006_ top.WB.CPU_DAT_O\[19\] net1220 net317 vssd1 vssd1 vccd1 vccd1 _01306_ sky130_fd_sc_hd__mux2_1
X_06218_ _03076_ _03085_ _03086_ vssd1 vssd1 vccd1 vccd1 _03087_ sky130_fd_sc_hd__or3b_1
XANTENNA_fanout793_A net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05643__A2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07198_ _03841_ _03844_ _03843_ vssd1 vssd1 vccd1 vccd1 _03856_ sky130_fd_sc_hd__a21o_1
XFILLER_117_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06149_ top.hist_addr\[1\] top.hist_addr\[0\] vssd1 vssd1 vccd1 vccd1 _03020_ sky130_fd_sc_hd__nand2_1
XFILLER_2_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08593__A1 top.cb_syn.char_index\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout531 top.cb_syn.curr_state\[7\] vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__clkbuf_2
Xfanout542 net543 vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__clkbuf_4
Xfanout520 top.translation.index\[3\] vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__clkbuf_4
Xfanout553 net555 vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__clkbuf_4
X_09908_ net761 net601 vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__and2_1
Xfanout575 net577 vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__clkbuf_2
Xfanout564 net567 vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__clkbuf_2
XFILLER_100_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09839_ net797 net637 vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__and2_1
XFILLER_86_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout586 net588 vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__clkbuf_2
Xfanout597 net647 vssd1 vssd1 vccd1 vccd1 net597 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_29_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ clknet_leaf_92_clk _02318_ _01156_ vssd1 vssd1 vccd1 vccd1 top.compVal\[33\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07940__S net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11732_ clknet_leaf_122_clk _02265_ _01087_ vssd1 vssd1 vccd1 vccd1 top.path\[63\]
+ sky130_fd_sc_hd__dfrtp_1
X_11663_ clknet_leaf_15_clk _02196_ _01018_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_25_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07608__B1 _04190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08056__B net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10614_ net768 net608 vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__and2_1
X_11594_ clknet_leaf_40_clk _02142_ _00949_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08805__C1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10545_ net832 net672 vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__and2_1
X_10476_ net844 net684 vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__and2_1
XFILLER_108_494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_75_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07792__C1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08336__A1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11028_ clknet_leaf_27_clk _01576_ _00383_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_49_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__07850__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05520_ net1200 net139 _02621_ net176 vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__a22o_1
X_05451_ net464 net561 vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__and2_1
XFILLER_82_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07151__A _03782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08170_ top.cb_syn.char_path_n\[84\] net202 _04612_ vssd1 vssd1 vccd1 vccd1 _01730_
+ sky130_fd_sc_hd__o21a_1
XFILLER_32_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07121_ top.findLeastValue.val1\[11\] top.findLeastValue.val2\[11\] _03731_ _03777_
+ _03778_ vssd1 vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__a221o_1
X_05382_ top.findLeastValue.val2\[22\] vssd1 vssd1 vccd1 vccd1 _02490_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_121_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_121_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08811__A2 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput101 net101 vssd1 vssd1 vccd1 vccd1 DAT_O[6] sky130_fd_sc_hd__buf_2
X_07052_ top.findLeastValue.val1\[15\] top.findLeastValue.val2\[15\] vssd1 vssd1 vccd1
+ vccd1 _03710_ sky130_fd_sc_hd__nand2_1
XANTENNA__05625__A2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06003_ net450 net466 top.histogram.state\[2\] vssd1 vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__and3_2
XANTENNA__07378__A2 _03423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08575__A1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_87_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07954_ top.findLeastValue.least1\[2\] top.findLeastValue.least2\[2\] _04462_ vssd1
+ vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__mux2_1
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__11844__Q top.WB.CPU_DAT_O\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06905_ top.findLeastValue.val2\[31\] net148 net124 _03594_ vssd1 vssd1 vccd1 vccd1
+ _01973_ sky130_fd_sc_hd__o22a_1
X_07885_ top.hTree.tree_reg\[11\] top.findLeastValue.sum\[11\] net247 vssd1 vssd1
+ vccd1 vccd1 _04414_ sky130_fd_sc_hd__mux2_1
X_09624_ net844 net684 vssd1 vssd1 vccd1 vccd1 _00238_ sky130_fd_sc_hd__and2_1
X_06836_ top.findLeastValue.least2\[7\] net152 net125 _03557_ vssd1 vssd1 vccd1 vccd1
+ _02005_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout374_A net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08422__S1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07760__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout639_A net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06767_ net501 net412 net118 net134 top.cw1\[4\] vssd1 vssd1 vccd1 vccd1 _02069_
+ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout162_X net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09555_ net733 net573 vssd1 vssd1 vccd1 vccd1 _00169_ sky130_fd_sc_hd__and2_1
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07838__B1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08506_ net1174 top.cb_syn.char_path_n\[70\] net226 vssd1 vssd1 vccd1 vccd1 _01588_
+ sky130_fd_sc_hd__mux2_1
X_09486_ net728 net568 vssd1 vssd1 vccd1 vccd1 _00100_ sky130_fd_sc_hd__and2_1
X_06698_ _02434_ top.findLeastValue.val2\[15\] _03477_ _03484_ vssd1 vssd1 vccd1 vccd1
+ _03486_ sky130_fd_sc_hd__o22a_1
X_05718_ net24 net418 net360 top.WB.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 _02340_
+ sky130_fd_sc_hd__a22o_1
XFILLER_24_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08437_ top.cb_syn.char_path_n\[38\] net330 _04795_ vssd1 vssd1 vccd1 vccd1 _04796_
+ sky130_fd_sc_hd__a21o_1
X_05649_ top.cb_syn.char_path\[5\] top.sram_interface.word_cnt\[0\] net316 top.cb_syn.char_path\[101\]
+ vssd1 vssd1 vccd1 vccd1 _02729_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout806_A net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08368_ net515 top.cb_syn.char_path_n\[119\] vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__or2_1
X_08299_ top.cb_syn.char_path_n\[20\] net376 net343 top.cb_syn.char_path_n\[18\] net188
+ vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__a221o_1
X_07319_ _03711_ _03946_ vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__or2_1
XANTENNA__08802__A2 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_112_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_112_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10330_ net793 net633 vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__and2_1
X_10261_ net871 net711 vssd1 vssd1 vccd1 vccd1 _00875_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_111_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07935__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10192_ net839 net679 vssd1 vssd1 vccd1 vccd1 _00806_ sky130_fd_sc_hd__and2_1
Xfanout350 net351 vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout383 net384 vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__buf_2
Xfanout372 _05085_ vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout361 net362 vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__clkbuf_4
Xfanout394 net395 vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07670__S net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11715_ clknet_leaf_121_clk _02248_ _01070_ vssd1 vssd1 vccd1 vccd1 top.path\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05855__A2 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11646_ clknet_leaf_113_clk _02179_ _01001_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput25 DAT_I[30] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__buf_1
Xinput36 gpio_in[2] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_2
Xinput14 DAT_I[20] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_103_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_103_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11577_ clknet_leaf_109_clk _02125_ _00932_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_116_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10528_ net849 net689 vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__and2_1
XANTENNA__05607__A2 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07845__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10459_ net723 net563 vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__and2_1
XFILLER_42_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07670_ top.findLeastValue.least2\[7\] top.hTree.tree_reg\[53\] net285 vssd1 vssd1
+ vccd1 vccd1 _04241_ sky130_fd_sc_hd__mux2_1
XFILLER_65_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06621_ _03389_ _03404_ _03407_ _03409_ vssd1 vssd1 vccd1 vccd1 _03410_ sky130_fd_sc_hd__or4_1
X_06552_ _02429_ top.findLeastValue.val1\[20\] vssd1 vssd1 vccd1 vccd1 _03341_ sky130_fd_sc_hd__and2_1
X_09340_ net994 net236 net214 _04426_ vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__a22o_1
X_09271_ _05213_ _05222_ _05223_ _05214_ net1642 vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_zero_count\[4\]
+ sky130_fd_sc_hd__a32o_1
X_05503_ top.cb_syn.char_path\[93\] net554 net545 top.cb_syn.char_path\[61\] vssd1
+ vssd1 vccd1 vccd1 _02607_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_51_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08222_ top.cb_syn.char_path_n\[58\] net207 _04638_ vssd1 vssd1 vccd1 vccd1 _01704_
+ sky130_fd_sc_hd__o21a_1
XFILLER_60_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06483_ net1723 _03288_ net1462 vssd1 vssd1 vccd1 vccd1 _03299_ sky130_fd_sc_hd__a21oi_1
X_05434_ top.header_synthesis.header\[8\] vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__inv_2
XANTENNA__06924__S net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05846__A2 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08153_ top.cb_syn.char_path_n\[93\] net387 net348 top.cb_syn.char_path_n\[91\] net193
+ vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__a221o_1
X_05365_ top.findLeastValue.least2\[8\] vssd1 vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout122_A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08084_ top.cb_syn.char_path_n\[127\] net207 _04569_ vssd1 vssd1 vccd1 vccd1 _01773_
+ sky130_fd_sc_hd__o21a_1
X_07104_ _03761_ vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__inv_2
X_05296_ net453 vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__inv_2
XANTENNA__11839__Q top.WB.CPU_DAT_O\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07035_ _03690_ _03692_ vssd1 vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__nor2_1
XANTENNA__07755__S net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05783__B net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08986_ top.WB.CPU_DAT_O\[6\] net1240 net324 vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__mux2_1
XFILLER_88_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07937_ net425 _04454_ _04455_ net258 vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout377_X net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout756_A net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07868_ net441 net1574 net253 top.findLeastValue.sum\[15\] _04400_ vssd1 vssd1 vccd1
+ vccd1 _01820_ sky130_fd_sc_hd__a221o_1
X_09607_ net844 net684 vssd1 vssd1 vccd1 vccd1 _00221_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout544_X net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07799_ top.findLeastValue.sum\[28\] top.hTree.tree_reg\[28\] net284 vssd1 vssd1
+ vccd1 vccd1 _04345_ sky130_fd_sc_hd__mux2_1
X_06819_ top.findLeastValue.val1\[11\] net128 net112 top.compVal\[11\] vssd1 vssd1
+ vccd1 vccd1 _02019_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_39_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09538_ net732 net572 vssd1 vssd1 vccd1 vccd1 _00152_ sky130_fd_sc_hd__and2_1
X_09469_ net749 net589 vssd1 vssd1 vccd1 vccd1 _00083_ sky130_fd_sc_hd__and2_1
X_11500_ clknet_leaf_90_clk _02048_ _00855_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[40\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__06834__S _03424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05837__A2 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11431_ clknet_leaf_88_clk _01979_ _00786_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[37\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_59_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11362_ clknet_leaf_101_clk _01910_ _00717_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08902__X _05072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10313_ net812 net652 vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__and2_1
XANTENNA__06798__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06262__A2 top.cb_syn.char_index\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11293_ clknet_leaf_84_clk net1402 _00648_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[36\]
+ sky130_fd_sc_hd__dfrtp_1
X_10244_ net828 net668 vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__and2_1
XANTENNA__07747__C1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10175_ net828 net668 vssd1 vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__and2_1
XFILLER_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07762__A2 _04314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout191 net193 vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__buf_2
Xfanout180 net181 vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__buf_2
XFILLER_74_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11629_ clknet_leaf_54_clk top.dut.bit_buf_next\[1\] _00984_ vssd1 vssd1 vccd1 vccd1
+ top.dut.bit_buf\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__08778__B2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold606 top.cb_syn.num_lefts\[7\] vssd1 vssd1 vccd1 vccd1 net1559 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06045__A net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold617 top.findLeastValue.sum\[41\] vssd1 vssd1 vccd1 vccd1 net1570 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06789__B1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold639 top.hTree.node_reg\[25\] vssd1 vssd1 vccd1 vccd1 net1592 sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 top.findLeastValue.sum\[25\] vssd1 vssd1 vccd1 vccd1 net1581 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_94_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08840_ _02522_ _04979_ _04982_ _05022_ top.translation.index\[4\] vssd1 vssd1 vccd1
+ vccd1 _05023_ sky130_fd_sc_hd__o311a_1
XFILLER_69_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05983_ _02909_ _02916_ vssd1 vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__nor2_1
XFILLER_85_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06961__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08771_ top.path\[85\] net327 _04953_ net433 net522 vssd1 vssd1 vccd1 vccd1 _04954_
+ sky130_fd_sc_hd__o221a_1
XANTENNA_clkbuf_4_7_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07722_ net426 _04282_ _04283_ net258 vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__o211a_1
XANTENNA__08163__C1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07653_ net486 _04225_ vssd1 vssd1 vccd1 vccd1 _04228_ sky130_fd_sc_hd__or2_1
XFILLER_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06604_ _02410_ top.findLeastValue.val1\[39\] vssd1 vssd1 vccd1 vccd1 _03393_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_36_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07584_ top.cb_syn.h_element\[57\] top.cb_syn.h_element\[48\] _04145_ vssd1 vssd1
+ vccd1 vccd1 _04171_ sky130_fd_sc_hd__mux2_1
X_09323_ top.translation.resEn _05257_ net431 vssd1 vssd1 vccd1 vccd1 _05258_ sky130_fd_sc_hd__o21ai_1
X_06535_ _02824_ _03323_ vssd1 vssd1 vccd1 vccd1 _03325_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout337_A net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_09254_ net518 top.header_synthesis.header\[8\] vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__or2_1
X_06466_ top.histogram.total\[24\] top.histogram.total\[23\] _03288_ vssd1 vssd1 vccd1
+ vccd1 _03289_ sky130_fd_sc_hd__and3_1
X_09185_ top.cb_syn.curr_state\[2\] net476 _04125_ _04868_ _05174_ vssd1 vssd1 vccd1
+ vccd1 _00004_ sky130_fd_sc_hd__a41o_1
X_05417_ top.cb_syn.max_index\[1\] vssd1 vssd1 vccd1 vccd1 _02525_ sky130_fd_sc_hd__inv_2
X_08205_ top.cb_syn.char_path_n\[67\] net381 net339 top.cb_syn.char_path_n\[65\] net185
+ vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__a221o_1
X_08136_ top.cb_syn.char_path_n\[101\] net201 _04595_ vssd1 vssd1 vccd1 vccd1 _01747_
+ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout125_X net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06397_ net1431 net299 _03234_ _03235_ vssd1 vssd1 vccd1 vccd1 _02122_ sky130_fd_sc_hd__a22o_1
XANTENNA__11569__Q top.histogram.sram_out\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05348_ top.hist_data_o\[0\] vssd1 vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__inv_2
X_08067_ _04125_ _04507_ vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__or2_1
X_07018_ top.findLeastValue.val1\[27\] top.findLeastValue.val2\[27\] vssd1 vssd1 vccd1
+ vccd1 _03676_ sky130_fd_sc_hd__or2_1
X_08969_ top.WB.CPU_DAT_O\[23\] net1199 net321 vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__mux2_1
XANTENNA__05755__B2 top.WB.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10931_ clknet_leaf_32_clk _01486_ _00286_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.zeroes\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10862_ clknet_leaf_77_clk _01448_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10793_ clknet_leaf_52_clk net1598 _00212_ vssd1 vssd1 vccd1 vccd1 top.histogram.state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_14_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05688__B _02760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11414_ clknet_leaf_101_clk _01962_ _00769_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[20\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__07968__C1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_73_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11345_ clknet_leaf_62_clk _01893_ _00700_ vssd1 vssd1 vccd1 vccd1 top.cw2\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_4_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08080__A net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11276_ clknet_leaf_78_clk _01824_ _00631_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_106_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10227_ net816 net656 vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__and2_1
XFILLER_94_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09326__D net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10115__A net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_88_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold3 top.cb_syn.curr_state\[3\] vssd1 vssd1 vccd1 vccd1 net956 sky130_fd_sc_hd__dlygate4sd3_1
X_10158_ net816 net656 vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__and2_1
X_10089_ net832 net672 vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_11_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08696__B1 _04875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08160__A2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_clkbuf_leaf_26_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06320_ top.hist_data_o\[14\] top.hist_data_o\[13\] _03182_ vssd1 vssd1 vccd1 vccd1
+ _03183_ sky130_fd_sc_hd__and3_1
X_06251_ _03116_ _03117_ net470 vssd1 vssd1 vccd1 vccd1 _03118_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_96_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_4_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_4_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__05682__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06182_ top.cb_syn.max_index\[6\] _03025_ _03027_ top.hTree.nullSumIndex\[5\] vssd1
+ vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__a22o_1
Xhold436 top.cb_syn.char_path\[115\] vssd1 vssd1 vccd1 vccd1 net1389 sky130_fd_sc_hd__dlygate4sd3_1
Xhold414 top.hTree.tree_reg\[59\] vssd1 vssd1 vccd1 vccd1 net1367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold403 top.hTree.nulls\[47\] vssd1 vssd1 vccd1 vccd1 net1356 sky130_fd_sc_hd__dlygate4sd3_1
Xhold425 top.path\[85\] vssd1 vssd1 vccd1 vccd1 net1378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold447 top.cb_syn.char_path\[61\] vssd1 vssd1 vccd1 vccd1 net1400 sky130_fd_sc_hd__dlygate4sd3_1
Xhold469 top.hTree.tree_reg\[33\] vssd1 vssd1 vccd1 vccd1 net1422 sky130_fd_sc_hd__dlygate4sd3_1
X_09941_ net743 net583 vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__and2_1
Xhold458 net102 vssd1 vssd1 vccd1 vccd1 net1411 sky130_fd_sc_hd__dlygate4sd3_1
X_09872_ net790 net630 vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__and2_1
XANTENNA__10025__A net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08823_ top.path\[0\] net410 _05005_ vssd1 vssd1 vccd1 vccd1 _05006_ sky130_fd_sc_hd__o21a_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05966_ _02581_ _02760_ _02851_ vssd1 vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout287_A _03325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08754_ top.path\[106\] top.path\[107\] net527 vssd1 vssd1 vccd1 vccd1 _04937_ sky130_fd_sc_hd__mux2_1
XFILLER_66_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07705_ net396 _04269_ vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__nand2_1
XANTENNA__09025__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08685_ top.cb_syn.zeroes\[7\] _04883_ vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout454_A net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05897_ net536 _02868_ vssd1 vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__nand2_1
XANTENNA__11852__Q top.WB.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_92_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_92_clk sky130_fd_sc_hd__clkbuf_8
X_07636_ net263 _04212_ _04213_ net1222 net446 vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__a32o_1
XFILLER_26_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout621_A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07567_ _04150_ _04156_ vssd1 vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__nand2_1
XFILLER_53_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout719_A net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09306_ top.histogram.total\[10\] top.histogram.total\[11\] top.translation.index\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05241_ sky130_fd_sc_hd__mux2_1
X_06518_ net1550 _03273_ vssd1 vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__nor2_1
X_09237_ _04917_ _05203_ net296 vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_char_added
+ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_101_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07498_ top.cb_syn.char_path_n\[64\] top.cb_syn.char_path_n\[63\] top.cb_syn.char_path_n\[62\]
+ top.cb_syn.char_path_n\[61\] net401 net352 vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__mux4_1
XFILLER_70_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout507_X net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06449_ top.histogram.total\[0\] _03271_ vssd1 vssd1 vccd1 vccd1 _03272_ sky130_fd_sc_hd__and2_1
X_09168_ net1597 net295 _05165_ vssd1 vssd1 vccd1 vccd1 _00033_ sky130_fd_sc_hd__a21o_1
XANTENNA__05673__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09099_ _02774_ _02843_ _03166_ _02559_ vssd1 vssd1 vccd1 vccd1 _05119_ sky130_fd_sc_hd__a211o_1
X_08119_ top.cb_syn.char_path_n\[110\] net373 net333 top.cb_syn.char_path_n\[108\]
+ net178 vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__a221o_1
XANTENNA__07965__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11130_ clknet_leaf_18_clk _01678_ _00485_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[32\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09167__A1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11061_ clknet_leaf_27_clk _01609_ _00416_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[91\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_76_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07717__A2 _04278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10012_ net818 net658 vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__and2_1
XANTENNA__09443__B net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input15_A DAT_I[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_83_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_clk sky130_fd_sc_hd__clkbuf_8
X_10914_ clknet_leaf_36_clk top.header_synthesis.next_enable _00269_ vssd1 vssd1 vccd1
+ vccd1 top.header_synthesis.enable sky130_fd_sc_hd__dfrtp_4
XFILLER_71_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08774__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10845_ clknet_leaf_106_clk _01431_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_119_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10776_ clknet_leaf_45_clk _01375_ _00195_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[52\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_119_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05664__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11328_ clknet_leaf_52_clk _01876_ _00683_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.curr_index\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07500__S1 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11259_ clknet_leaf_83_clk _01807_ _00614_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08366__C1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07706__X _04271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05820_ net1036 net449 _02581_ vssd1 vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__a21o_1
XANTENNA__05719__B2 top.WB.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_74_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_clk sky130_fd_sc_hd__clkbuf_8
X_05751_ top.compVal\[43\] net172 net158 top.WB.CPU_DAT_O\[11\] vssd1 vssd1 vccd1
+ vccd1 _02328_ sky130_fd_sc_hd__a22o_1
XANTENNA__09330__A1 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08133__A2 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05682_ top.histogram.sram_out\[0\] net367 net422 top.hTree.node_reg\[0\] _02756_
+ vssd1 vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_46_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_08470_ net1247 top.cb_syn.char_path_n\[106\] net221 vssd1 vssd1 vccd1 vccd1 _01624_
+ sky130_fd_sc_hd__mux2_1
X_07421_ top.dut.bit_buf\[5\] net43 net722 vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__mux2_1
XFILLER_90_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07352_ _03744_ _03745_ _03746_ _03759_ vssd1 vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__a211o_1
X_06303_ top.sram_interface.word_cnt\[12\] net463 net546 _02937_ _03166_ vssd1 vssd1
+ vccd1 vccd1 _03167_ sky130_fd_sc_hd__a221o_1
X_07283_ net1643 _03658_ net268 _03919_ vssd1 vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__a22o_1
X_06234_ top.TRN_char_index\[2\] top.TRN_char_index\[1\] vssd1 vssd1 vccd1 vccd1 _03102_
+ sky130_fd_sc_hd__or2_1
XANTENNA__05655__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06932__S net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09022_ top.WB.CPU_DAT_O\[3\] net1207 net320 vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__mux2_1
XFILLER_116_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold211 top.cb_syn.char_path\[28\] vssd1 vssd1 vccd1 vccd1 net1164 sky130_fd_sc_hd__dlygate4sd3_1
X_06165_ _02560_ _02977_ _03029_ _03033_ _03035_ vssd1 vssd1 vccd1 vccd1 _03036_ sky130_fd_sc_hd__o311a_1
Xhold200 top.cb_syn.char_path\[2\] vssd1 vssd1 vccd1 vccd1 net1153 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 top.path\[99\] vssd1 vssd1 vccd1 vccd1 net1197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold222 top.path\[77\] vssd1 vssd1 vccd1 vccd1 net1175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 top.cb_syn.char_path\[77\] vssd1 vssd1 vccd1 vccd1 net1186 sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 net93 vssd1 vssd1 vccd1 vccd1 net1219 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06096_ top.cb_syn.char_index\[6\] _02579_ _02961_ _02968_ vssd1 vssd1 vccd1 vccd1
+ _02969_ sky130_fd_sc_hd__a31o_1
XANTENNA__09149__A1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold277 top.cb_syn.char_path\[51\] vssd1 vssd1 vccd1 vccd1 net1230 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 net80 vssd1 vssd1 vccd1 vccd1 net1208 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11847__Q top.WB.CPU_DAT_O\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout713 net716 vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__clkbuf_2
Xfanout702 net703 vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__clkbuf_2
X_09924_ net788 net628 vssd1 vssd1 vccd1 vccd1 _00538_ sky130_fd_sc_hd__and2_1
Xhold288 top.path\[18\] vssd1 vssd1 vccd1 vccd1 net1241 sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 top.path\[1\] vssd1 vssd1 vccd1 vccd1 net1252 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout724 net727 vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07616__X _04197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09855_ net739 net579 vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__and2_1
XANTENNA_input7_A DAT_I[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout746 net748 vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__clkbuf_2
Xfanout757 net807 vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__clkbuf_2
Xfanout735 net737 vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__clkbuf_2
Xfanout779 net786 vssd1 vssd1 vccd1 vccd1 net779 sky130_fd_sc_hd__buf_1
XFILLER_100_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout768 net769 vssd1 vssd1 vccd1 vccd1 net768 sky130_fd_sc_hd__clkbuf_2
X_08806_ top.path\[62\] top.path\[63\] net525 vssd1 vssd1 vccd1 vccd1 _04989_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout571_A net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout669_A net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06907__B1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06998_ _03652_ _03653_ _03654_ _03655_ vssd1 vssd1 vccd1 vccd1 _03656_ sky130_fd_sc_hd__and4_1
X_09786_ net741 net581 vssd1 vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__and2_1
XANTENNA__06383__A1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08737_ top.cb_syn.zeroes\[7\] top.cb_syn.zeroes\[6\] _04892_ _04920_ top.cb_syn.state8
+ vssd1 vssd1 vccd1 vccd1 _04921_ sky130_fd_sc_hd__o41a_2
Xclkbuf_leaf_65_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_clk sky130_fd_sc_hd__clkbuf_8
X_05949_ top.WB.CPU_DAT_O\[6\] net1448 net307 vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__mux2_1
XFILLER_39_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout836_A net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08668_ net536 net538 vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__nor2_1
XFILLER_53_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08124__A2 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07619_ top.findLeastValue.least1\[8\] net394 net248 top.hTree.tree_reg\[63\] vssd1
+ vssd1 vccd1 vccd1 _04200_ sky130_fd_sc_hd__o22ai_1
XFILLER_53_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07883__A1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10630_ net853 net693 vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__and2_1
X_08599_ top.CB_write_complete top.CB_read_complete top.cb_syn.curr_state\[8\] vssd1
+ vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__and3b_1
XANTENNA__07883__B2 top.findLeastValue.sum\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10561_ net854 net694 vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__and2_1
X_10492_ net826 net666 vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__and2_1
XANTENNA__05966__B _02760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11113_ clknet_leaf_6_clk _01661_ _00468_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[15\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_clkbuf_4_15_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08348__C1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11044_ clknet_leaf_11_clk _01592_ _00399_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[74\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_36_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_56_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07323__B1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11877_ clknet_leaf_39_clk _02393_ _01232_ vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__dfrtp_1
XFILLER_60_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10828_ clknet_leaf_79_clk _01414_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_10759_ clknet_leaf_43_clk _01358_ _00178_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07626__A1 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05637__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06053__A _02767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07485__S0 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06062__B1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07970_ _02764_ _03326_ _04476_ _03565_ top.findLeastValue.alternator_timer\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__a32o_1
XANTENNA__05892__A top.cb_syn.h_element\[63\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07583__S _04144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06921_ top.findLeastValue.val2\[23\] net146 net120 _03602_ vssd1 vssd1 vccd1 vccd1
+ _01965_ sky130_fd_sc_hd__o22a_1
XANTENNA__09000__A0 top.WB.CPU_DAT_O\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08354__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09640_ net804 net644 vssd1 vssd1 vccd1 vccd1 _00254_ sky130_fd_sc_hd__and2_1
X_06852_ net423 net287 vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__nand2_1
X_06783_ net1393 net134 _03547_ net126 _03554_ vssd1 vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__a32o_1
X_09571_ net796 net636 vssd1 vssd1 vccd1 vccd1 _00185_ sky130_fd_sc_hd__and2_1
X_05803_ top.hTree.state\[8\] _02811_ _02813_ vssd1 vssd1 vccd1 vccd1 _02823_ sky130_fd_sc_hd__and3_1
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10022__B net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05734_ _02763_ _02768_ vssd1 vssd1 vccd1 vccd1 _02769_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_47_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_clk sky130_fd_sc_hd__clkbuf_8
X_08522_ net1300 top.cb_syn.char_path_n\[54\] net230 vssd1 vssd1 vccd1 vccd1 _01572_
+ sky130_fd_sc_hd__mux2_1
X_08453_ net1381 top.cb_syn.char_path_n\[123\] net231 vssd1 vssd1 vccd1 vccd1 _01641_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09303__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07404_ top.dut.bit_buf\[11\] top.dut.bit_buf\[4\] net720 vssd1 vssd1 vccd1 vccd1
+ _04004_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout152_A net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05665_ net1106 net145 _02742_ net177 vssd1 vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__a22o_1
XANTENNA__07865__A1 top.findLeastValue.sum\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08384_ top.cb_syn.char_path_n\[99\] top.cb_syn.char_path_n\[100\] net513 vssd1 vssd1
+ vccd1 vccd1 _04743_ sky130_fd_sc_hd__mux2_1
X_05596_ net457 top.hTree.node_reg\[46\] net361 net421 top.hTree.node_reg\[14\] vssd1
+ vssd1 vccd1 vccd1 _02685_ sky130_fd_sc_hd__a32o_1
XANTENNA__08814__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07335_ net270 _03957_ _03958_ net275 net1714 vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_21_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07266_ _03699_ _03906_ vssd1 vssd1 vccd1 vccd1 _03908_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout417_A net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06217_ _02560_ _02975_ _03082_ _03081_ _03071_ vssd1 vssd1 vccd1 vccd1 _03086_ sky130_fd_sc_hd__o311a_1
X_09005_ top.WB.CPU_DAT_O\[20\] net1274 net318 vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__mux2_1
X_07197_ _03837_ _03838_ _03846_ _03854_ vssd1 vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__a211o_1
X_06148_ top.sram_interface.init_counter\[7\] _02946_ vssd1 vssd1 vccd1 vccd1 _03019_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout786_A net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06079_ _02566_ _02580_ _02951_ _02952_ vssd1 vssd1 vccd1 vccd1 _02953_ sky130_fd_sc_hd__or4_1
Xfanout532 net533 vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__buf_2
Xfanout510 top.cb_syn.end_cnt\[1\] vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__clkbuf_4
X_09907_ net787 net627 vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__and2_1
Xfanout521 net522 vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__clkbuf_4
XFILLER_116_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xfanout554 net555 vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__clkbuf_2
Xfanout543 net547 vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__buf_2
XANTENNA_fanout574_X net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout565 net567 vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__clkbuf_2
X_09838_ net782 net622 vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__and2_1
XFILLER_74_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout598 net599 vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__clkbuf_2
Xfanout576 net577 vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__clkbuf_2
Xfanout587 net588 vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__clkbuf_2
X_09769_ net782 net622 vssd1 vssd1 vccd1 vccd1 _00383_ sky130_fd_sc_hd__and2_1
XFILLER_18_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08750__C1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05307__A top.compVal\[33\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_38_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_8
X_11800_ clknet_leaf_92_clk _02317_ _01155_ vssd1 vssd1 vccd1 vccd1 top.compVal\[32\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__06108__B2 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06837__S _03424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ clknet_leaf_122_clk _02264_ _01086_ vssd1 vssd1 vccd1 vccd1 top.path\[62\]
+ sky130_fd_sc_hd__dfrtp_1
X_11662_ clknet_leaf_15_clk _02195_ _01017_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11593_ clknet_leaf_16_clk _02141_ _00948_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10613_ net768 net608 vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__and2_1
XANTENNA__08805__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10544_ net833 net673 vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__and2_1
XANTENNA__05619__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08072__B top.cb_syn.h_element\[54\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10475_ net856 net696 vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__and2_1
XFILLER_108_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08499__S net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08336__A2 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11027_ clknet_leaf_26_clk _01575_ _00382_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[57\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_29_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_86_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05570__A2 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_05450_ net481 _02557_ vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__and2_2
XFILLER_20_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05381_ top.findLeastValue.val2\[24\] vssd1 vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__inv_2
X_07120_ top.findLeastValue.val1\[11\] top.findLeastValue.val2\[11\] top.findLeastValue.val2\[10\]
+ top.findLeastValue.val1\[10\] vssd1 vssd1 vccd1 vccd1 _03778_ sky130_fd_sc_hd__o211a_1
XANTENNA__09078__B net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07051_ top.findLeastValue.val1\[15\] top.findLeastValue.val2\[15\] vssd1 vssd1 vccd1
+ vccd1 _03709_ sky130_fd_sc_hd__nor2_1
X_06002_ net458 net423 net422 top.hTree.write_HT_fin vssd1 vssd1 vccd1 vccd1 _02207_
+ sky130_fd_sc_hd__o22a_1
Xoutput102 net102 vssd1 vssd1 vccd1 vccd1 DAT_O[7] sky130_fd_sc_hd__buf_2
XFILLER_114_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07953_ net1497 _04466_ _04461_ vssd1 vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__mux2_1
XANTENNA__07607__A net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_06904_ top.compVal\[31\] top.findLeastValue.val1\[31\] net162 vssd1 vssd1 vccd1
+ vccd1 _03594_ sky130_fd_sc_hd__mux2_1
X_07884_ top.findLeastValue.sum\[11\] top.hTree.tree_reg\[11\] net283 vssd1 vssd1
+ vccd1 vccd1 _04413_ sky130_fd_sc_hd__mux2_1
X_09623_ net844 net684 vssd1 vssd1 vccd1 vccd1 _00237_ sky130_fd_sc_hd__and2_1
X_06835_ _03553_ _03556_ vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__and2b_1
XANTENNA__06889__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06766_ net499 net413 net118 net134 net1612 vssd1 vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__a32o_1
XANTENNA__05561__A2 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09554_ net734 net574 vssd1 vssd1 vccd1 vccd1 _00168_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout534_A net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07838__A1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07838__B2 top.findLeastValue.sum\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08505_ net1104 top.cb_syn.char_path_n\[71\] net226 vssd1 vssd1 vccd1 vccd1 _01589_
+ sky130_fd_sc_hd__mux2_1
X_06697_ _02435_ top.findLeastValue.val2\[14\] _03476_ vssd1 vssd1 vccd1 vccd1 _03485_
+ sky130_fd_sc_hd__or3_1
X_05717_ net27 net418 net360 top.WB.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 _02341_
+ sky130_fd_sc_hd__a22o_1
X_09485_ net732 net572 vssd1 vssd1 vccd1 vccd1 _00099_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout155_X net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08436_ top.cb_syn.char_path_n\[37\] net393 _04776_ net509 net438 vssd1 vssd1 vccd1
+ vccd1 _04795_ sky130_fd_sc_hd__a221o_1
X_05648_ top.cb_syn.char_path\[69\] net552 net543 top.cb_syn.char_path\[37\] vssd1
+ vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__a22o_1
XANTENNA__05849__B1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08367_ net511 _04724_ _04725_ vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout701_A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05579_ top.histogram.sram_out\[17\] net364 _02669_ _02670_ vssd1 vssd1 vccd1 vccd1
+ _02671_ sky130_fd_sc_hd__a211o_1
X_07318_ _03713_ _03945_ _03712_ vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__a21bo_1
XFILLER_109_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_08298_ top.cb_syn.char_path_n\[20\] net204 _04676_ vssd1 vssd1 vccd1 vccd1 _01666_
+ sky130_fd_sc_hd__o21a_1
X_07249_ _03830_ _03893_ vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__or2_1
XANTENNA__06813__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10260_ net872 net712 vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__and2_1
XFILLER_117_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07369__A3 _03547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10191_ net863 net703 vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__and2_1
XANTENNA__11100__Q top.cb_syn.char_path_n\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout340 net341 vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_6_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout384 net390 vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__buf_2
Xfanout362 _02583_ vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout351 net353 vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__clkbuf_4
Xfanout373 net374 vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__buf_2
XANTENNA__08318__A2 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09154__D _02767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout395 _04195_ vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__buf_4
XANTENNA__05537__C1 _02635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05552__A2 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11714_ clknet_leaf_121_clk _02247_ _01069_ vssd1 vssd1 vccd1 vccd1 top.path\[45\]
+ sky130_fd_sc_hd__dfrtp_1
X_11645_ clknet_leaf_113_clk _02178_ _01000_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput37 gpio_in[3] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_1
Xinput26 DAT_I[31] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
Xinput15 DAT_I[21] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
X_11576_ clknet_leaf_109_clk _02124_ _00931_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08254__A1 top.cb_syn.char_path_n\[42\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10527_ net849 net689 vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__and2_1
XANTENNA__06804__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10118__A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10458_ net728 net568 vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__and2_1
X_10389_ net756 net596 vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__and2_1
XFILLER_96_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06620_ _02412_ top.findLeastValue.val1\[36\] _03394_ _03408_ vssd1 vssd1 vccd1 vccd1
+ _03409_ sky130_fd_sc_hd__a211o_1
XFILLER_92_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__05543__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06551_ _02428_ top.findLeastValue.val1\[21\] top.findLeastValue.val1\[20\] _02429_
+ _03339_ vssd1 vssd1 vccd1 vccd1 _03340_ sky130_fd_sc_hd__o221a_1
X_09270_ top.cb_syn.zero_count\[4\] _05219_ vssd1 vssd1 vccd1 vccd1 _05223_ sky130_fd_sc_hd__or2_1
X_05502_ net1418 net139 _02606_ net175 vssd1 vssd1 vccd1 vccd1 _02400_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_51_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06482_ _03290_ _03298_ vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__nor2_1
X_05433_ net1 vssd1 vssd1 vccd1 vccd1 _02541_ sky130_fd_sc_hd__inv_2
X_08221_ top.cb_syn.char_path_n\[59\] net384 net345 top.cb_syn.char_path_n\[57\] net190
+ vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_99_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08152_ top.cb_syn.char_path_n\[93\] net208 _04603_ vssd1 vssd1 vccd1 vccd1 _01739_
+ sky130_fd_sc_hd__o21a_1
X_05364_ top.findLeastValue.val1\[26\] vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08083_ top.cb_syn.curr_path\[127\] net385 net344 top.cb_syn.char_path_n\[126\] net189
+ vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_9_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_8
X_07103_ _03746_ _03759_ _03744_ _03745_ vssd1 vssd1 vccd1 vccd1 _03761_ sky130_fd_sc_hd__o211a_1
XANTENNA__08796__A2 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_3_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10028__A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__06835__A_N _03553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout115_A net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07034_ top.findLeastValue.val1\[30\] top.findLeastValue.val2\[30\] vssd1 vssd1 vccd1
+ vccd1 _03692_ sky130_fd_sc_hd__nor2_1
XANTENNA__06940__S net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05783__C net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08985_ top.WB.CPU_DAT_O\[7\] net1318 net324 vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout484_A net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07936_ net482 _04453_ vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__or2_1
XFILLER_113_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05519__C1 _02620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08181__B1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07867_ net426 _04398_ _04399_ net261 vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout272_X net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout651_A net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09606_ net843 net683 vssd1 vssd1 vccd1 vccd1 _00220_ sky130_fd_sc_hd__and2_1
XANTENNA__05534__A2 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07798_ net446 net1403 net254 net1730 _04344_ vssd1 vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__a221o_1
X_06818_ top.findLeastValue.val1\[12\] net129 net113 top.compVal\[12\] vssd1 vssd1
+ vccd1 vccd1 _02020_ sky130_fd_sc_hd__o22a_1
XFILLER_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09537_ net750 net590 vssd1 vssd1 vccd1 vccd1 _00151_ sky130_fd_sc_hd__and2_1
X_06749_ _03534_ _03536_ _03531_ vssd1 vssd1 vccd1 vccd1 _03537_ sky130_fd_sc_hd__or3b_1
X_09468_ net753 net593 vssd1 vssd1 vccd1 vccd1 _00082_ sky130_fd_sc_hd__and2_1
X_09399_ net969 _05276_ net244 vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__mux2_1
X_08419_ top.cb_syn.char_path_n\[43\] top.cb_syn.char_path_n\[44\] net514 vssd1 vssd1
+ vccd1 vccd1 _04778_ sky130_fd_sc_hd__mux2_1
X_11430_ clknet_leaf_88_clk _01978_ _00785_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[36\]
+ sky130_fd_sc_hd__dfstp_1
X_11361_ clknet_leaf_97_clk _01909_ _00716_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_20_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10312_ net763 net603 vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__and2_1
X_11292_ clknet_leaf_84_clk net1428 _00647_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[35\]
+ sky130_fd_sc_hd__dfrtp_1
X_10243_ net828 net668 vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__and2_1
X_10174_ net832 net672 vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__and2_1
XFILLER_93_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout192 net193 vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__clkbuf_2
Xfanout181 net194 vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__clkbuf_2
Xfanout170 net171 vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__buf_2
XFILLER_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05525__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10401__A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08475__A1 top.cb_syn.char_path_n\[101\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11628_ clknet_leaf_55_clk top.dut.bit_buf_next\[0\] _00983_ vssd1 vssd1 vccd1 vccd1
+ top.dut.bit_buf\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_7_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08778__A2 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11559_ clknet_leaf_37_clk _02107_ _00914_ vssd1 vssd1 vccd1 vccd1 top.header_synthesis.count\[0\]
+ sky130_fd_sc_hd__dfrtp_2
Xhold607 top.histogram.total\[1\] vssd1 vssd1 vccd1 vccd1 net1560 sky130_fd_sc_hd__dlygate4sd3_1
Xhold618 top.hTree.tree_reg\[12\] vssd1 vssd1 vccd1 vccd1 net1571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold629 top.hTree.tree_reg\[14\] vssd1 vssd1 vccd1 vccd1 net1582 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_94_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07738__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06410__A0 top.histogram.sram_out\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05982_ top.sram_interface.init_counter\[9\] _02915_ vssd1 vssd1 vccd1 vccd1 _02916_
+ sky130_fd_sc_hd__nor2_1
X_08770_ top.path\[86\] top.path\[87\] net526 vssd1 vssd1 vccd1 vccd1 _04953_ sky130_fd_sc_hd__mux2_1
X_07721_ net483 _04281_ vssd1 vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__or2_1
XANTENNA__05516__A2 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07652_ net486 _04226_ vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__nand2_1
X_07583_ net1596 _04170_ _04144_ vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__mux2_1
XFILLER_25_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06603_ _02413_ top.findLeastValue.val1\[35\] vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__nand2_1
X_06534_ _02824_ _03323_ vssd1 vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__nor2_1
X_09322_ top.translation.totalEn _05255_ _05256_ vssd1 vssd1 vccd1 vccd1 _05257_ sky130_fd_sc_hd__a21oi_1
XFILLER_80_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_09253_ net1077 _05211_ _04918_ vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_header\[7\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout232_A net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07620__A net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06465_ top.histogram.total\[22\] _03287_ vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__and2_1
X_09184_ net475 _02863_ _02932_ _04139_ _05173_ vssd1 vssd1 vccd1 vccd1 _05174_ sky130_fd_sc_hd__a221o_1
X_08204_ top.cb_syn.char_path_n\[67\] net201 _04629_ vssd1 vssd1 vccd1 vccd1 _01713_
+ sky130_fd_sc_hd__o21a_1
X_05416_ net523 vssd1 vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__inv_2
X_06396_ net299 _03178_ vssd1 vssd1 vccd1 vccd1 _03235_ sky130_fd_sc_hd__nor2_1
X_05347_ net457 vssd1 vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__inv_2
X_08135_ top.cb_syn.char_path_n\[102\] net380 net339 top.cb_syn.char_path_n\[100\]
+ net184 vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout118_X net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08066_ _02506_ _04546_ _04553_ vssd1 vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout699_A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07017_ _03665_ _03669_ _03667_ _03664_ vssd1 vssd1 vccd1 vccd1 _03675_ sky130_fd_sc_hd__a211o_1
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout866_A net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08968_ top.WB.CPU_DAT_O\[24\] net1346 net322 vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__mux2_1
X_08899_ top.cb_syn.max_index\[7\] _05067_ _05068_ vssd1 vssd1 vccd1 vccd1 _05069_
+ sky130_fd_sc_hd__o21a_1
X_07919_ top.findLeastValue.sum\[4\] top.hTree.tree_reg\[4\] net278 vssd1 vssd1 vccd1
+ vccd1 _04441_ sky130_fd_sc_hd__mux2_1
X_10930_ clknet_leaf_32_clk _01485_ _00285_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.zeroes\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05507__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10861_ clknet_leaf_46_clk _01447_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[53\]
+ sky130_fd_sc_hd__dfxtp_1
X_10792_ clknet_leaf_53_clk _00032_ _00211_ vssd1 vssd1 vccd1 vccd1 top.histogram.eof_n
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__06845__S _03424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05602__X _02690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XTAP_TAPCELL_ROW_14_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11413_ clknet_leaf_101_clk _01961_ _00768_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[19\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__05691__B2 top.WB.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11344_ clknet_leaf_63_clk _01892_ _00699_ vssd1 vssd1 vccd1 vccd1 top.cw2\[4\] sky130_fd_sc_hd__dfrtp_1
X_11275_ clknet_leaf_79_clk net1445 _00630_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_106_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__09185__A2 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08080__B net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10226_ net816 net656 vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__and2_1
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10115__B net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold4 top.controller.fin_HG vssd1 vssd1 vccd1 vccd1 net957 sky130_fd_sc_hd__dlygate4sd3_1
X_10157_ net816 net656 vssd1 vssd1 vccd1 vccd1 _00771_ sky130_fd_sc_hd__and2_1
X_10088_ net867 net707 vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__and2_1
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05512__X _02615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06250_ net502 net368 _02572_ _03114_ _03112_ vssd1 vssd1 vccd1 vccd1 _03117_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_96_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05682__A1 top.histogram.sram_out\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06181_ _02943_ _03049_ _03050_ net495 net466 vssd1 vssd1 vccd1 vccd1 _03051_ sky130_fd_sc_hd__o221a_1
Xhold415 top.cb_syn.char_path\[60\] vssd1 vssd1 vccd1 vccd1 net1368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold426 top.cb_syn.char_path\[104\] vssd1 vssd1 vccd1 vccd1 net1379 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold404 top.path\[116\] vssd1 vssd1 vccd1 vccd1 net1357 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold459 top.cb_syn.count\[7\] vssd1 vssd1 vccd1 vccd1 net1412 sky130_fd_sc_hd__dlygate4sd3_1
X_09940_ net761 net601 vssd1 vssd1 vccd1 vccd1 _00554_ sky130_fd_sc_hd__and2_1
Xhold448 top.hTree.tree_reg\[36\] vssd1 vssd1 vccd1 vccd1 net1401 sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 top.path\[5\] vssd1 vssd1 vccd1 vccd1 net1390 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_115_Right_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09871_ net790 net630 vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__and2_1
XANTENNA__10025__B net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08822_ top.path\[1\] net328 _05004_ net434 net437 vssd1 vssd1 vccd1 vccd1 _05005_
+ sky130_fd_sc_hd__o221a_1
X_05965_ _02529_ _02779_ _02901_ net1602 vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__o22a_1
X_08753_ _04932_ _04933_ _04934_ net437 net520 vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__a221o_1
XANTENNA__09306__S top.translation.index\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07704_ top.findLeastValue.least2\[1\] top.hTree.tree_reg\[47\] net281 vssd1 vssd1
+ vccd1 vccd1 _04269_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout182_A net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08684_ _04875_ _04134_ vssd1 vssd1 vccd1 vccd1 _04885_ sky130_fd_sc_hd__and2b_2
X_05896_ _02870_ vssd1 vssd1 vccd1 vccd1 _02871_ sky130_fd_sc_hd__inv_2
XFILLER_81_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07635_ net489 _04210_ vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout447_A net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07566_ top.cb_syn.max_index\[5\] _04149_ top.cb_syn.max_index\[6\] vssd1 vssd1 vccd1
+ vccd1 _04156_ sky130_fd_sc_hd__o21ai_1
XFILLER_80_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09305_ top.histogram.total\[13\] net327 _05238_ net433 net521 vssd1 vssd1 vccd1
+ vccd1 _05240_ sky130_fd_sc_hd__o221a_1
X_06517_ net1524 _03275_ vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__xor2_1
X_09236_ net518 top.header_synthesis.char_added vssd1 vssd1 vccd1 vccd1 _05203_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout235_X net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07497_ top.cb_syn.char_path_n\[60\] top.cb_syn.char_path_n\[59\] top.cb_syn.char_path_n\[58\]
+ top.cb_syn.char_path_n\[57\] net401 net352 vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout614_A net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06448_ _03269_ _03270_ top.controller.state_reg\[4\] vssd1 vssd1 vccd1 vccd1 _03271_
+ sky130_fd_sc_hd__o21a_1
X_09167_ net449 net295 top.histogram.state\[5\] vssd1 vssd1 vccd1 vccd1 _05165_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout402_X net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06379_ top.hist_data_o\[13\] _03182_ vssd1 vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__xor2_1
XFILLER_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09098_ net468 top.sram_interface.word_cnt\[7\] _02777_ _05117_ vssd1 vssd1 vccd1
+ vccd1 _05118_ sky130_fd_sc_hd__a31o_1
X_08118_ top.cb_syn.char_path_n\[110\] net195 _04586_ vssd1 vssd1 vccd1 vccd1 _01756_
+ sky130_fd_sc_hd__o21a_1
X_08049_ top.cb_syn.end_cnt\[6\] top.cb_syn.end_cnt\[5\] _04541_ vssd1 vssd1 vccd1
+ vccd1 _04543_ sky130_fd_sc_hd__or3_1
X_11060_ clknet_leaf_27_clk _01608_ _00415_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[90\]
+ sky130_fd_sc_hd__dfrtp_1
X_10011_ net818 net658 vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__and2_1
XFILLER_103_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08127__B1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10913_ clknet_leaf_38_clk _01471_ _00268_ vssd1 vssd1 vccd1 vccd1 top.header_synthesis.bit1
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_80_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10844_ clknet_leaf_107_clk _01430_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_4_11_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10775_ clknet_leaf_15_clk _01374_ _00194_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05664__A1 top.histogram.sram_out\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11327_ clknet_leaf_52_clk _01875_ _00682_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.curr_index\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08366__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11258_ clknet_leaf_105_clk _01806_ _00613_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11189_ clknet_leaf_27_clk _01737_ _00544_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[91\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__05719__A2 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10209_ net826 net666 vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__and2_1
XFILLER_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_19_Left_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05750_ top.compVal\[44\] net172 net158 top.WB.CPU_DAT_O\[12\] vssd1 vssd1 vccd1
+ vccd1 _02329_ sky130_fd_sc_hd__a22o_1
XFILLER_82_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_05681_ top.hTree.node_reg\[32\] net311 _02755_ net480 vssd1 vssd1 vccd1 vccd1 _02756_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_46_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07420_ _04001_ _04013_ _04018_ vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__a21o_1
XFILLER_50_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07351_ net270 _03967_ _03968_ net275 top.findLeastValue.sum\[5\] vssd1 vssd1 vccd1
+ vccd1 _01901_ sky130_fd_sc_hd__a32o_1
X_06302_ net550 top.sram_interface.word_cnt\[13\] net541 net459 vssd1 vssd1 vccd1
+ vccd1 _03166_ sky130_fd_sc_hd__o31a_1
X_07282_ _03684_ _03898_ vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__xor2_1
X_06233_ _02974_ net562 vssd1 vssd1 vccd1 vccd1 _03101_ sky130_fd_sc_hd__and2b_1
X_09021_ top.WB.CPU_DAT_O\[4\] net1362 net320 vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_28_Left_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06164_ _02565_ _02973_ _03030_ _03034_ vssd1 vssd1 vccd1 vccd1 _03035_ sky130_fd_sc_hd__o31a_1
Xhold201 top.cb_syn.char_path\[63\] vssd1 vssd1 vccd1 vccd1 net1154 sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 top.cb_syn.char_path\[100\] vssd1 vssd1 vccd1 vccd1 net1187 sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 top.cb_syn.char_path\[7\] vssd1 vssd1 vccd1 vccd1 net1165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 top.path\[20\] vssd1 vssd1 vccd1 vccd1 net1176 sky130_fd_sc_hd__dlygate4sd3_1
X_06095_ top.cb_syn.char_index\[6\] _02578_ _02963_ _02967_ vssd1 vssd1 vccd1 vccd1
+ _02968_ sky130_fd_sc_hd__a31o_1
Xhold256 top.sram_interface.word_cnt\[11\] vssd1 vssd1 vccd1 vccd1 net1209 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold245 top.path\[70\] vssd1 vssd1 vccd1 vccd1 net1198 sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 top.path\[83\] vssd1 vssd1 vccd1 vccd1 net1220 sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 top.histogram.sram_out\[10\] vssd1 vssd1 vccd1 vccd1 net1231 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout714 net716 vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06080__B2 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout703 net706 vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__clkbuf_2
X_09923_ net776 net616 vssd1 vssd1 vccd1 vccd1 _00537_ sky130_fd_sc_hd__and2_1
Xhold289 top.cb_syn.char_path\[36\] vssd1 vssd1 vccd1 vccd1 net1242 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout397_A net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09854_ net739 net579 vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__and2_1
Xfanout736 net737 vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_0_Left_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout747 net748 vssd1 vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__clkbuf_2
Xfanout725 net727 vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__clkbuf_2
Xfanout758 net759 vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__clkbuf_2
XFILLER_85_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout769 net772 vssd1 vssd1 vccd1 vccd1 net769 sky130_fd_sc_hd__clkbuf_2
X_08805_ top.path\[20\] net408 net326 top.path\[21\] net521 vssd1 vssd1 vccd1 vccd1
+ _04988_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_37_Left_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06997_ top.findLeastValue.val1\[18\] top.findLeastValue.val1\[17\] top.findLeastValue.val1\[16\]
+ top.findLeastValue.val1\[15\] vssd1 vssd1 vccd1 vccd1 _03655_ sky130_fd_sc_hd__and4_1
X_09785_ net758 net598 vssd1 vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__and2_1
X_08736_ top.cb_syn.zeroes\[5\] top.cb_syn.zeroes\[4\] top.cb_syn.zeroes\[3\] top.cb_syn.zeroes\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04920_ sky130_fd_sc_hd__or4_1
XANTENNA__05591__B1 _02679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05948_ top.WB.CPU_DAT_O\[7\] net1250 net307 vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__mux2_1
X_08667_ _04132_ _04867_ _04869_ vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout352_X net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05879_ top.sram_interface.zero_cnt\[0\] _02853_ net1655 vssd1 vssd1 vccd1 vccd1
+ _02856_ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_72_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout731_A net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08447__Y _04805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07618_ net394 net285 vssd1 vssd1 vccd1 vccd1 _04199_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout829_A net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08598_ _04819_ net518 _04817_ vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__mux2_1
X_07549_ net540 _02869_ _04132_ _04139_ vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_62_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_46_Left_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_87_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10560_ net854 net694 vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__and2_1
X_09219_ top.controller.fin_reg\[5\] _05190_ net1709 top.controller.fin_reg\[7\] vssd1
+ vssd1 vccd1 vccd1 _05191_ sky130_fd_sc_hd__or4b_1
X_10491_ net826 net666 vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__and2_1
XFILLER_107_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_10_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11112_ clknet_leaf_6_clk _01660_ _00467_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_25_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_55_Left_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08348__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11043_ clknet_leaf_110_clk _01591_ _00398_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[73\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_3_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_3_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__05582__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09312__A2 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_64_Left_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11876_ clknet_leaf_100_clk _02392_ _01231_ vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__dfrtp_1
X_10827_ clknet_leaf_78_clk _01413_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_10758_ clknet_leaf_44_clk _01357_ _00177_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[52\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06834__A0 top.findLeastValue.least1\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10689_ clknet_leaf_114_clk _01288_ _00108_ vssd1 vssd1 vccd1 vccd1 top.path\[65\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_114_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07485__S1 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_73_Left_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06920_ top.compVal\[23\] top.findLeastValue.val1\[23\] net161 vssd1 vssd1 vccd1
+ vccd1 _03602_ sky130_fd_sc_hd__mux2_1
X_06851_ net470 net288 vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__nor2_1
X_06782_ top.findLeastValue.wipe_the_char_1 net167 _03553_ vssd1 vssd1 vccd1 vccd1
+ _03554_ sky130_fd_sc_hd__a21o_1
X_09570_ net795 net635 vssd1 vssd1 vccd1 vccd1 _00184_ sky130_fd_sc_hd__and2_1
X_05802_ net556 _02821_ net461 vssd1 vssd1 vccd1 vccd1 _02822_ sky130_fd_sc_hd__o21ai_1
X_05733_ top.findLeastValue.alternator_timer\[3\] top.findLeastValue.alternator_timer\[2\]
+ net414 vssd1 vssd1 vccd1 vccd1 _02768_ sky130_fd_sc_hd__o21ai_1
X_08521_ net1373 top.cb_syn.char_path_n\[55\] net230 vssd1 vssd1 vccd1 vccd1 _01573_
+ sky130_fd_sc_hd__mux2_1
XFILLER_70_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08452_ net1189 top.cb_syn.char_path_n\[124\] net231 vssd1 vssd1 vccd1 vccd1 _01642_
+ sky130_fd_sc_hd__mux2_1
X_07403_ top.dut.bit_buf\[12\] top.dut.bit_buf\[5\] net722 vssd1 vssd1 vccd1 vccd1
+ _04003_ sky130_fd_sc_hd__mux2_1
X_05664_ top.histogram.sram_out\[3\] net367 net422 top.hTree.node_reg\[3\] _02741_
+ vssd1 vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__a221o_1
XANTENNA__05413__A top.translation.index\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout145_A _02595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08383_ net509 _04740_ _04741_ vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__a21oi_1
X_05595_ _02682_ _02683_ net472 vssd1 vssd1 vccd1 vccd1 _02684_ sky130_fd_sc_hd__o21a_1
X_07334_ _03727_ _03956_ _03730_ vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_21_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07265_ _03699_ _03906_ vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__or2_1
XANTENNA__06825__B1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06216_ net478 _03078_ _03079_ net460 _03084_ vssd1 vssd1 vccd1 vccd1 _03085_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout312_A net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09004_ top.WB.CPU_DAT_O\[21\] net1378 net318 vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__mux2_1
X_07196_ _03850_ _03853_ vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__or2_1
XFILLER_105_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06147_ net497 _02550_ _02572_ _03017_ _03016_ vssd1 vssd1 vccd1 vccd1 _03018_ sky130_fd_sc_hd__a221o_1
X_06078_ net548 net368 net413 net469 vssd1 vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__o211a_1
XANTENNA__07250__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout779_A net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout533 net534 vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__clkbuf_2
Xfanout511 top.cb_syn.end_cnt\[1\] vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__clkbuf_4
Xfanout500 top.findLeastValue.histo_index\[4\] vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__buf_2
X_09906_ net787 net627 vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout681_A net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout522 top.translation.index\[2\] vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__clkbuf_4
Xfanout555 top.sram_interface.word_cnt\[3\] vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__clkbuf_4
Xfanout544 net547 vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__clkbuf_4
Xfanout566 net567 vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__clkbuf_2
X_09837_ net778 net618 vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__and2_1
XFILLER_58_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout577 net585 vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__clkbuf_2
Xfanout588 net597 vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__clkbuf_2
Xfanout599 net602 vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__clkbuf_2
X_09768_ net775 net615 vssd1 vssd1 vccd1 vccd1 _00382_ sky130_fd_sc_hd__and2_1
XANTENNA__05564__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08750__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08719_ _04902_ _04905_ _04908_ _04898_ net1638 vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__a32o_1
XFILLER_27_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06108__A2 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09699_ net863 net703 vssd1 vssd1 vccd1 vccd1 _00313_ sky130_fd_sc_hd__and2_1
X_11730_ clknet_leaf_121_clk _02263_ _01085_ vssd1 vssd1 vccd1 vccd1 top.path\[61\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_1_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout734_X net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11661_ clknet_leaf_15_clk _02194_ _01016_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_42_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05867__B2 top.WB.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11592_ clknet_leaf_45_clk _02140_ _00947_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10612_ net739 net579 vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__and2_1
XANTENNA__06816__B1 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10543_ net832 net672 vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__and2_1
XANTENNA__05610__X _02697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10474_ net873 net713 vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_75_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11026_ clknet_leaf_26_clk _01574_ _00381_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08741__B1 top.header_synthesis.bit1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05555__B1 _02649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05858__B2 top.WB.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11859_ clknet_leaf_100_clk _02375_ _01214_ vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09049__A1 top.WB.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05380_ top.findLeastValue.val2\[25\] vssd1 vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__inv_2
XANTENNA__07859__S net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06807__B1 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07050_ _03682_ _03706_ _03707_ _03677_ vssd1 vssd1 vccd1 vccd1 _03708_ sky130_fd_sc_hd__o211a_1
X_06001_ _02903_ _02925_ vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__nor2_1
XFILLER_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_81_Left_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 DAT_O[8] sky130_fd_sc_hd__buf_2
XFILLER_99_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06035__A1 top.WB.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08980__A0 top.WB.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07607__B _04188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07952_ top.findLeastValue.least1\[3\] top.findLeastValue.least2\[3\] _04462_ vssd1
+ vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__mux2_1
X_06903_ top.findLeastValue.val2\[32\] net153 net125 _03593_ vssd1 vssd1 vccd1 vccd1
+ _01974_ sky130_fd_sc_hd__o22a_1
X_07883_ net442 net1571 net251 top.findLeastValue.sum\[12\] _04412_ vssd1 vssd1 vccd1
+ vccd1 _01817_ sky130_fd_sc_hd__a221o_1
XFILLER_83_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05546__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06834_ top.findLeastValue.least1\[7\] _02481_ _03424_ vssd1 vssd1 vccd1 vccd1 _03556_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__06938__S net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09622_ net759 net599 vssd1 vssd1 vccd1 vccd1 _00236_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_90_Left_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09553_ net732 net572 vssd1 vssd1 vccd1 vccd1 _00167_ sky130_fd_sc_hd__and2_1
X_06765_ top.findLeastValue.histo_index\[6\] net413 net118 net135 net1577 vssd1 vssd1
+ vccd1 vccd1 _02071_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout262_A net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08504_ net1190 top.cb_syn.char_path_n\[72\] net226 vssd1 vssd1 vccd1 vccd1 _01590_
+ sky130_fd_sc_hd__mux2_1
X_05716_ net28 net416 net309 top.WB.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 _02342_
+ sky130_fd_sc_hd__o22a_1
X_06696_ _03479_ _03480_ _03478_ vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__a21oi_1
X_09484_ net727 net567 vssd1 vssd1 vccd1 vccd1 _00098_ sky130_fd_sc_hd__and2_1
XANTENNA__07299__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08435_ net509 _04777_ _04793_ vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__a21o_1
X_05647_ net1395 net138 _02727_ net174 vssd1 vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__a22o_1
XANTENNA__05849__B2 top.WB.CPU_DAT_O\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08366_ top.cb_syn.char_path_n\[121\] net392 net331 top.cb_syn.char_path_n\[122\]
+ net507 vssd1 vssd1 vccd1 vccd1 _04725_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout527_A net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05578_ net457 top.hTree.node_reg\[49\] net361 net420 top.hTree.node_reg\[17\] vssd1
+ vssd1 vccd1 vccd1 _02670_ sky130_fd_sc_hd__a32o_1
X_07317_ _03725_ _03944_ _03716_ vssd1 vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout315_X net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08297_ top.cb_syn.char_path_n\[21\] net383 net342 top.cb_syn.char_path_n\[19\] net187
+ vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__a221o_1
XFILLER_109_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07248_ _03830_ _03893_ vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__nand2_1
X_07179_ _03817_ _03820_ _03831_ _03672_ vssd1 vssd1 vccd1 vccd1 _03837_ sky130_fd_sc_hd__a211o_1
X_10190_ net863 net703 vssd1 vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__and2_1
XANTENNA__06026__A1 top.WB.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08420__C1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08971__A0 top.WB.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout341 net349 vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__buf_2
Xfanout330 net332 vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout352 net353 vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout374 net377 vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__buf_2
Xfanout363 net364 vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__buf_2
Xfanout385 net386 vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__buf_2
XFILLER_86_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05537__B1 _02634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout396 net397 vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__buf_2
X_11713_ clknet_leaf_121_clk _02246_ _01068_ vssd1 vssd1 vccd1 vccd1 top.path\[44\]
+ sky130_fd_sc_hd__dfrtp_1
X_11644_ clknet_leaf_113_clk _02177_ _00999_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput27 DAT_I[3] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
Xinput16 DAT_I[22] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
X_11575_ clknet_leaf_109_clk _02123_ _00930_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput38 gpio_in[4] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_1
X_10526_ net860 net700 vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__and2_1
X_10457_ net729 net569 vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__and2_1
XFILLER_108_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09195__A _03325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06017__A1 top.WB.CPU_DAT_O\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10388_ net756 net596 vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__and2_1
XANTENNA__08962__A0 top.WB.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09923__A net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05528__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_11009_ clknet_leaf_12_clk _01557_ _00364_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_52_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06550_ _02426_ top.findLeastValue.val1\[23\] top.findLeastValue.val1\[22\] _02427_
+ vssd1 vssd1 vccd1 vccd1 _03339_ sky130_fd_sc_hd__o22a_1
X_05501_ top.histogram.sram_out\[30\] net365 _02604_ _02605_ vssd1 vssd1 vccd1 vccd1
+ _02606_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_51_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06481_ net1511 _03289_ vssd1 vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__nor2_1
XANTENNA__07730__X _04290_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05432_ top.header_synthesis.write_num_lefts vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__inv_2
X_08220_ top.cb_syn.char_path_n\[59\] net207 _04637_ vssd1 vssd1 vccd1 vccd1 _01705_
+ sky130_fd_sc_hd__o21a_1
XFILLER_60_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08151_ top.cb_syn.char_path_n\[94\] net387 net346 top.cb_syn.char_path_n\[92\] net191
+ vssd1 vssd1 vccd1 vccd1 _04603_ sky130_fd_sc_hd__a221o_1
XANTENNA__08245__A2 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05363_ top.findLeastValue.val1\[27\] vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08082_ net1505 net190 _04568_ vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__a21o_1
X_07102_ _03759_ vssd1 vssd1 vccd1 vccd1 _03760_ sky130_fd_sc_hd__inv_2
X_07033_ top.findLeastValue.val1\[30\] top.findLeastValue.val2\[30\] vssd1 vssd1 vccd1
+ vccd1 _03691_ sky130_fd_sc_hd__nand2_1
XANTENNA__06008__A1 top.WB.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07618__A net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08953__A0 top.WB.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10044__A net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08984_ top.WB.CPU_DAT_O\[8\] net1397 net323 vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07935_ top.findLeastValue.sum\[1\] _04453_ net395 vssd1 vssd1 vccd1 vccd1 _04454_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout477_A net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09605_ net804 net644 vssd1 vssd1 vccd1 vccd1 _00219_ sky130_fd_sc_hd__and2_1
XANTENNA__05519__B1 _02619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07866_ net483 _04397_ vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__or2_1
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07797_ net430 _04342_ _04343_ net263 vssd1 vssd1 vccd1 vccd1 _04344_ sky130_fd_sc_hd__o211a_1
X_06817_ top.findLeastValue.val1\[13\] net129 net113 top.compVal\[13\] vssd1 vssd1
+ vccd1 vccd1 _02021_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_39_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_09536_ net749 net589 vssd1 vssd1 vccd1 vccd1 _00150_ sky130_fd_sc_hd__and2_1
X_06748_ _03530_ _03535_ _03532_ vssd1 vssd1 vccd1 vccd1 _03536_ sky130_fd_sc_hd__or3b_1
XANTENNA__09130__B1 _02899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09467_ net752 net592 vssd1 vssd1 vccd1 vccd1 _00081_ sky130_fd_sc_hd__and2_1
X_08418_ top.cb_syn.char_path_n\[35\] top.cb_syn.char_path_n\[36\] net513 vssd1 vssd1
+ vccd1 vccd1 _04777_ sky130_fd_sc_hd__mux2_1
X_06679_ _02443_ top.findLeastValue.val2\[6\] top.findLeastValue.val2\[5\] _02444_
+ vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout811_A net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09398_ top.hTree.nulls\[53\] _04242_ net406 vssd1 vssd1 vccd1 vccd1 _05276_ sky130_fd_sc_hd__mux2_1
X_08349_ net509 _04706_ _04707_ vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__a21o_1
X_11360_ clknet_leaf_97_clk _01908_ _00715_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[12\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_118_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__08912__A _04187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10311_ net818 net658 vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__and2_1
XANTENNA__06798__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11291_ clknet_leaf_84_clk _01839_ _00646_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05766__D_N top.TRN_sram_complete vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08944__A0 top.WB.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10242_ net834 net674 vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__and2_1
X_10173_ net842 net682 vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__and2_1
XANTENNA_input38_A gpio_in[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout160 _02594_ vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__clkbuf_4
Xfanout182 net194 vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__buf_2
Xfanout171 _02845_ vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__clkbuf_2
Xfanout193 net194 vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__buf_2
XFILLER_86_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10401__B net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05930__A0 top.WB.CPU_DAT_O\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11627_ clknet_leaf_53_clk top.dut.out_valid_next _00982_ vssd1 vssd1 vccd1 vccd1
+ top.dut.out_valid sky130_fd_sc_hd__dfrtp_1
XANTENNA__10129__A net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06238__A1 top.cb_syn.char_index\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11558_ clknet_leaf_123_clk _02106_ _00913_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xhold608 top.cw1\[3\] vssd1 vssd1 vccd1 vccd1 net1561 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06789__A2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10509_ net813 net653 vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__and2_1
Xhold619 top.cw2\[3\] vssd1 vssd1 vccd1 vccd1 net1572 sky130_fd_sc_hd__dlygate4sd3_1
X_11489_ clknet_leaf_90_clk _02037_ _00844_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[29\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_94_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08935__A0 top.WB.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07738__A1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05981_ net1506 _02909_ vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__xor2_1
X_07720_ top.hTree.tree_reg\[44\] top.findLeastValue.sum\[44\] net249 vssd1 vssd1
+ vccd1 vccd1 _04282_ sky130_fd_sc_hd__mux2_1
XANTENNA__06961__A2 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07651_ top.findLeastValue.least1\[2\] net249 _04224_ vssd1 vssd1 vccd1 vccd1 _04226_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_92_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07582_ top.cb_syn.max_index\[4\] _04136_ _04166_ _04169_ vssd1 vssd1 vccd1 vccd1
+ _04170_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_36_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06602_ _02406_ top.findLeastValue.val1\[45\] top.findLeastValue.val1\[46\] vssd1
+ vssd1 vccd1 vccd1 _03391_ sky130_fd_sc_hd__a21oi_1
X_06533_ _02812_ _02816_ vssd1 vssd1 vccd1 vccd1 _03323_ sky130_fd_sc_hd__nand2_1
X_09321_ top.translation.totalEn _05032_ _04925_ top.translation.writeEn vssd1 vssd1
+ vccd1 vccd1 _05256_ sky130_fd_sc_hd__and4bb_1
X_09252_ top.header_synthesis.header\[7\] top.cb_syn.char_index\[7\] net519 vssd1
+ vssd1 vccd1 vccd1 _05211_ sky130_fd_sc_hd__mux2_1
X_06464_ top.histogram.total\[21\] top.histogram.total\[20\] _03286_ vssd1 vssd1 vccd1
+ vccd1 _03287_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_16_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09183_ _02932_ _04478_ _05095_ _02526_ vssd1 vssd1 vccd1 vccd1 _05173_ sky130_fd_sc_hd__a211oi_1
XANTENNA__08218__A2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08203_ top.cb_syn.char_path_n\[68\] net380 net340 top.cb_syn.char_path_n\[66\] net184
+ vssd1 vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__a221o_1
X_05415_ net521 vssd1 vssd1 vccd1 vccd1 _02523_ sky130_fd_sc_hd__inv_2
X_06395_ top.hist_data_o\[6\] _03174_ _03176_ top.hist_data_o\[7\] vssd1 vssd1 vccd1
+ vccd1 _03234_ sky130_fd_sc_hd__a31o_1
XFILLER_119_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05346_ top.hTree.write_HT_fin vssd1 vssd1 vccd1 vccd1 _02454_ sky130_fd_sc_hd__inv_2
X_08134_ top.cb_syn.char_path_n\[102\] net202 _04594_ vssd1 vssd1 vccd1 vccd1 _01748_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__07521__S0 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08065_ net512 _04553_ _04551_ vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__a21o_1
XFILLER_108_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08926__A0 top.WB.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07016_ top.findLeastValue.val1\[39\] top.findLeastValue.val2\[39\] _03673_ vssd1
+ vssd1 vccd1 vccd1 _03674_ sky130_fd_sc_hd__a21oi_1
XFILLER_88_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout594_A net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08878__S net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout382_X net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout859_A net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08967_ top.WB.CPU_DAT_O\[25\] net1332 net322 vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__mux2_1
X_08898_ top.cb_syn.max_index\[7\] _05067_ _04187_ vssd1 vssd1 vccd1 vccd1 _05068_
+ sky130_fd_sc_hd__a21oi_1
X_07918_ net440 net1584 net251 top.findLeastValue.sum\[5\] _04440_ vssd1 vssd1 vccd1
+ vccd1 _01810_ sky130_fd_sc_hd__a221o_1
XFILLER_84_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09351__B1 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07849_ top.findLeastValue.sum\[18\] top.hTree.tree_reg\[18\] net278 vssd1 vssd1
+ vccd1 vccd1 _04385_ sky130_fd_sc_hd__mux2_1
XFILLER_16_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout647_X net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10860_ clknet_leaf_46_clk _01446_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[52\]
+ sky130_fd_sc_hd__dfxtp_1
X_09519_ net740 net580 vssd1 vssd1 vccd1 vccd1 _00133_ sky130_fd_sc_hd__and2_1
X_10791_ clknet_leaf_51_clk _00031_ _00210_ vssd1 vssd1 vccd1 vccd1 top.histogram.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11412_ clknet_leaf_100_clk _01960_ _00767_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[18\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__08642__A net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07968__A1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11343_ clknet_leaf_64_clk _01891_ _00698_ vssd1 vssd1 vccd1 vccd1 top.cw2\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_4_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11274_ clknet_leaf_106_clk _01822_ _00629_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10225_ net816 net656 vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__and2_1
X_10156_ net813 net653 vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__and2_1
X_10087_ net872 net712 vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__and2_1
Xhold5 top.controller.fin_FLV vssd1 vssd1 vccd1 vccd1 net958 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload3_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05903__B1 top.CB_write_complete vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10989_ clknet_leaf_22_clk _01537_ _00344_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06056__B net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05682__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06180_ top.hist_addr\[6\] _03022_ vssd1 vssd1 vccd1 vccd1 _03050_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_96_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07503__S0 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold405 top.cb_syn.char_path\[25\] vssd1 vssd1 vccd1 vccd1 net1358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold427 top.path\[46\] vssd1 vssd1 vccd1 vccd1 net1380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold416 top.path\[72\] vssd1 vssd1 vccd1 vccd1 net1369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 _01841_ vssd1 vssd1 vccd1 vccd1 net1402 sky130_fd_sc_hd__dlygate4sd3_1
Xhold438 top.path\[81\] vssd1 vssd1 vccd1 vccd1 net1391 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_98_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09870_ net778 net618 vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__and2_1
XANTENNA__08908__B1 _04188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08821_ top.path\[2\] top.path\[3\] net528 vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__mux2_1
X_05964_ top.sram_interface.word_cnt\[1\] net468 _02548_ _02777_ vssd1 vssd1 vccd1
+ vccd1 _02901_ sky130_fd_sc_hd__and4_1
XANTENNA__08136__A1 top.cb_syn.char_path_n\[101\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08752_ net522 _04927_ _04930_ _02522_ vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__a211o_1
X_08683_ _04134_ _04883_ _04875_ vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__a21o_1
X_07703_ net263 _04267_ _04268_ net1023 net447 vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__a32o_1
XANTENNA__05416__A net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout175_A net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05895_ top.cb_syn.wait_cycle _02526_ vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__nor2_1
X_07634_ net489 _04211_ vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_49_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06946__S net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07565_ net532 top.cb_syn.h_element\[51\] net539 top.cb_syn.h_element\[60\] _04135_
+ vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout342_A net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07496_ top.cb_syn.char_path_n\[56\] top.cb_syn.char_path_n\[55\] top.cb_syn.char_path_n\[54\]
+ top.cb_syn.char_path_n\[53\] net401 net352 vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__mux4_1
XANTENNA__08844__C1 top.translation.index\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09304_ top.histogram.total\[12\] net409 vssd1 vssd1 vccd1 vccd1 _05239_ sky130_fd_sc_hd__or2_1
X_06516_ _03277_ _03312_ vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__nor2_1
XANTENNA__05422__Y _02530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09235_ net518 net1599 _03251_ vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_start
+ sky130_fd_sc_hd__o21a_1
X_06447_ top.dut.out_valid top.histogram.eof_n top.histogram.out_of_init vssd1 vssd1
+ vccd1 vccd1 _03270_ sky130_fd_sc_hd__and3b_4
XFILLER_119_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_fanout228_X net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout607_A net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_119_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_09166_ net366 _05101_ _05103_ top.histogram.eof_n vssd1 vssd1 vccd1 vccd1 _00032_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__06870__B2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05673__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06378_ net1142 _03223_ net300 vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__mux2_1
X_09097_ net562 top.sram_interface.word_cnt\[9\] _02561_ net478 vssd1 vssd1 vccd1
+ vccd1 _05117_ sky130_fd_sc_hd__o211a_1
X_08117_ top.cb_syn.char_path_n\[111\] net373 net333 top.cb_syn.char_path_n\[109\]
+ net178 vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__a221o_1
X_05329_ top.compVal\[12\] vssd1 vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_116_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08048_ top.cb_syn.end_cnt\[5\] net246 _04541_ top.cb_syn.end_cnt\[6\] vssd1 vssd1
+ vccd1 vccd1 _04542_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout597_X net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10010_ net818 net658 vssd1 vssd1 vccd1 vccd1 _00624_ sky130_fd_sc_hd__and2_1
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09999_ net820 net660 vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__and2_1
XANTENNA__07806__A net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09324__B1 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10912_ clknet_leaf_32_clk top.header_synthesis.next_zero_count\[7\] _00267_ vssd1
+ vssd1 vccd1 vccd1 top.cb_syn.zero_count\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_84_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11892_ clknet_leaf_53_clk net919 _01247_ vssd1 vssd1 vccd1 vccd1 top.dut.bits_in_buf\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10843_ clknet_leaf_84_clk _01429_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07638__A0 top.findLeastValue.least1\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10774_ clknet_leaf_107_clk _01373_ _00193_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05664__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11326_ clknet_leaf_52_clk _01874_ _00681_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.curr_index\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11257_ clknet_leaf_90_clk _01805_ _00612_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11188_ clknet_leaf_27_clk _01736_ _00543_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[90\]
+ sky130_fd_sc_hd__dfrtp_2
X_10208_ net826 net666 vssd1 vssd1 vccd1 vccd1 _00822_ sky130_fd_sc_hd__and2_1
X_10139_ net830 net670 vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__and2_1
XANTENNA__09931__A net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05680_ _02753_ _02754_ vssd1 vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_46_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05523__X _02624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_07350_ _03763_ _03765_ vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__nand2_1
XANTENNA__08981__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06301_ top.sram_interface.word_cnt\[9\] net316 net480 vssd1 vssd1 vccd1 vccd1 _03165_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_100_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07597__S _04144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06301__B1 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09020_ top.WB.CPU_DAT_O\[5\] net1471 net319 vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__mux2_1
X_07281_ net268 _03917_ _03918_ net273 net1581 vssd1 vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__a32o_1
X_06232_ net495 _03098_ _03099_ _02943_ net467 vssd1 vssd1 vccd1 vccd1 _03100_ sky130_fd_sc_hd__o221a_1
XANTENNA__05655__A2 top.sram_interface.word_cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06163_ top.cb_syn.curr_index\[7\] _02558_ _03028_ net460 vssd1 vssd1 vccd1 vccd1
+ _03034_ sky130_fd_sc_hd__a22oi_1
Xhold202 top.cb_syn.char_path\[93\] vssd1 vssd1 vccd1 vccd1 net1155 sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 top.histogram.sram_out\[24\] vssd1 vssd1 vccd1 vccd1 net1177 sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 top.cb_syn.char_path\[82\] vssd1 vssd1 vccd1 vccd1 net1188 sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 top.path\[66\] vssd1 vssd1 vccd1 vccd1 net1166 sky130_fd_sc_hd__dlygate4sd3_1
X_06094_ net414 _02965_ _02966_ net470 vssd1 vssd1 vccd1 vccd1 _02967_ sky130_fd_sc_hd__o211a_1
Xhold257 top.cb_syn.char_path\[78\] vssd1 vssd1 vccd1 vccd1 net1210 sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 top.path\[4\] vssd1 vssd1 vccd1 vccd1 net1221 sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 top.path\[119\] vssd1 vssd1 vccd1 vccd1 net1199 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout715 net716 vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__buf_1
XANTENNA__06080__A2 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout704 net705 vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__clkbuf_2
Xhold279 top.cb_syn.char_path\[24\] vssd1 vssd1 vccd1 vccd1 net1232 sky130_fd_sc_hd__dlygate4sd3_1
X_09922_ net774 net614 vssd1 vssd1 vccd1 vccd1 _00536_ sky130_fd_sc_hd__and2_1
XFILLER_100_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09853_ net738 net578 vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__and2_1
Xfanout737 net745 vssd1 vssd1 vccd1 vccd1 net737 sky130_fd_sc_hd__clkbuf_2
Xfanout748 net757 vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__clkbuf_2
Xfanout726 net727 vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10052__A net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08804_ net432 _04986_ vssd1 vssd1 vccd1 vccd1 _04987_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout292_A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09784_ net758 net598 vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__and2_1
Xfanout759 net762 vssd1 vssd1 vccd1 vccd1 net759 sky130_fd_sc_hd__clkbuf_2
X_08735_ top.header_synthesis.count\[3\] _02540_ _03259_ _03260_ vssd1 vssd1 vccd1
+ vccd1 _04919_ sky130_fd_sc_hd__or4_1
X_06996_ top.findLeastValue.val1\[22\] top.findLeastValue.val1\[21\] top.findLeastValue.val1\[20\]
+ top.findLeastValue.val1\[19\] vssd1 vssd1 vccd1 vccd1 _03654_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout557_A net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05947_ top.WB.CPU_DAT_O\[8\] net1382 net306 vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__mux2_1
X_08666_ _04868_ _04555_ vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__and2b_1
X_05878_ _02855_ net1683 vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__and2b_1
XFILLER_26_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07868__B1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08597_ net439 _02861_ _04818_ vssd1 vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__o21ai_1
X_07617_ _02459_ _02473_ _02801_ _04196_ vssd1 vssd1 vccd1 vccd1 _04198_ sky130_fd_sc_hd__or4_2
XANTENNA__09052__S net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07548_ top.cb_syn.setup top.cb_syn.curr_state\[0\] vssd1 vssd1 vccd1 vccd1 _04139_
+ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_24_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_101_Left_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07479_ _04049_ _04051_ vssd1 vssd1 vccd1 vccd1 _04070_ sky130_fd_sc_hd__nor2_2
XANTENNA__08904__B _04187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08293__B1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08832__A2 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09218_ _05188_ _05190_ vssd1 vssd1 vccd1 vccd1 _00016_ sky130_fd_sc_hd__nor2_1
XANTENNA__06843__A1 top.findLeastValue.histo_index\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10490_ net826 net666 vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__and2_1
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_09149_ net541 _05154_ _05156_ net550 vssd1 vssd1 vccd1 vccd1 _05157_ sky130_fd_sc_hd__a22o_1
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_11111_ clknet_leaf_6_clk _01659_ _00466_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__05608__X _02695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11042_ clknet_leaf_11_clk _01590_ _00397_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[72\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_110_Left_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input20_A DAT_I[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11875_ clknet_leaf_70_clk _02391_ _01230_ vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__dfrtp_1
XFILLER_45_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07323__A2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10826_ clknet_leaf_78_clk _01412_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_44_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_43_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10757_ clknet_leaf_44_clk _01356_ _00176_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08823__A2 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05637__A2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10688_ clknet_leaf_114_clk _01287_ _00107_ vssd1 vssd1 vccd1 vccd1 top.path\[64\]
+ sky130_fd_sc_hd__dfrtp_1
X_11309_ clknet_leaf_76_clk _01857_ _00664_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[52\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05518__X _02620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06850_ top.findLeastValue.least2\[0\] net136 _03547_ net126 _03564_ vssd1 vssd1
+ vccd1 vccd1 _01998_ sky130_fd_sc_hd__a32o_1
XFILLER_95_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05801_ net550 net548 top.sram_interface.word_cnt\[13\] net541 vssd1 vssd1 vccd1
+ vccd1 _02821_ sky130_fd_sc_hd__or4_1
XANTENNA__08976__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06781_ net167 _03546_ _03545_ net414 vssd1 vssd1 vccd1 vccd1 _03553_ sky130_fd_sc_hd__and4bb_4
XFILLER_48_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08520_ net1224 top.cb_syn.char_path_n\[56\] net230 vssd1 vssd1 vccd1 vccd1 _01574_
+ sky130_fd_sc_hd__mux2_1
X_05732_ top.findLeastValue.histo_index\[8\] top.findLeastValue.histo_index\[7\] vssd1
+ vssd1 vccd1 vccd1 _02767_ sky130_fd_sc_hd__or2_4
XANTENNA__09380__B _04271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08451_ net1330 top.cb_syn.char_path_n\[125\] net231 vssd1 vssd1 vccd1 vccd1 _01643_
+ sky130_fd_sc_hd__mux2_1
X_05663_ top.hTree.node_reg\[35\] net311 _02740_ net480 vssd1 vssd1 vccd1 vccd1 _02741_
+ sky130_fd_sc_hd__a22o_1
XFILLER_51_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07402_ _04001_ vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__inv_2
X_08382_ top.cb_syn.char_path_n\[101\] net391 net330 top.cb_syn.char_path_n\[102\]
+ net438 vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__a221o_1
X_05594_ top.cb_syn.char_path\[14\] net557 net312 top.cb_syn.char_path\[110\] vssd1
+ vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__a22o_1
XANTENNA__08814__A2 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07333_ _03727_ _03730_ _03956_ vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_21_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07264_ _03700_ _03900_ vssd1 vssd1 vccd1 vccd1 _03906_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout138_A net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06215_ _02971_ _03083_ _02564_ vssd1 vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__and3b_1
X_09003_ top.WB.CPU_DAT_O\[22\] net1080 net318 vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__mux2_1
XANTENNA__06244__B _02767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07195_ _03851_ _03852_ vssd1 vssd1 vccd1 vccd1 _03853_ sky130_fd_sc_hd__nand2_1
X_06146_ top.cw2\[7\] _03005_ vssd1 vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__xor2_1
X_06077_ _02942_ _02948_ _02950_ net449 vssd1 vssd1 vccd1 vccd1 _02951_ sky130_fd_sc_hd__a31oi_1
XFILLER_104_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__07250__A1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout501 top.findLeastValue.histo_index\[4\] vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__buf_1
Xfanout512 top.cb_syn.end_cnt\[1\] vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__clkbuf_2
X_09905_ net788 net628 vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__and2_1
XANTENNA__09047__S net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout523 top.translation.index\[1\] vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__buf_4
Xfanout534 net535 vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__clkbuf_2
XFILLER_98_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout545 net547 vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__clkbuf_2
Xfanout556 top.sram_interface.word_cnt\[1\] vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__buf_2
XFILLER_58_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout674_A net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09836_ net778 net618 vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__and2_1
Xfanout578 net579 vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__clkbuf_2
XFILLER_46_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout589 net590 vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__clkbuf_2
Xfanout567 net574 vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07790__S net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout462_X net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09767_ net775 net615 vssd1 vssd1 vccd1 vccd1 _00381_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout841_A net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06979_ top.findLeastValue.val2\[46\] top.findLeastValue.val2\[45\] top.findLeastValue.val2\[44\]
+ top.findLeastValue.val2\[43\] vssd1 vssd1 vccd1 vccd1 _03637_ sky130_fd_sc_hd__and4_1
X_08718_ top.cb_syn.i\[4\] _04900_ vssd1 vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__or2_1
X_09698_ net867 net707 vssd1 vssd1 vccd1 vccd1 _00312_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_29_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08649_ top.cb_syn.cb_length\[2\] _02927_ vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_1_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11660_ clknet_leaf_14_clk _02193_ _01015_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_11591_ clknet_leaf_44_clk _02139_ _00946_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10611_ net739 net579 vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_115_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_115_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08805__A2 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10542_ net832 net672 vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__and2_1
XFILLER_22_381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__05619__A2 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10473_ net728 net568 vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_75_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07777__C1 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06044__A2 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06170__A net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11025_ clknet_leaf_20_clk _01573_ _00380_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07553__X _04144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11858_ clknet_leaf_115_clk _02374_ _01213_ vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__dfrtp_1
X_11789_ clknet_leaf_75_clk _00024_ _01144_ vssd1 vssd1 vccd1 vccd1 top.hTree.state\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_106_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_106_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10809_ clknet_leaf_105_clk _01395_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06000_ top.sram_interface.init_counter\[0\] _02902_ vssd1 vssd1 vccd1 vccd1 _02925_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__05491__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_71_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 DAT_O[9] sky130_fd_sc_hd__buf_2
XFILLER_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07951_ net1629 _04465_ _04461_ vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__mux2_1
X_06902_ top.compVal\[32\] top.findLeastValue.val1\[32\] net165 vssd1 vssd1 vccd1
+ vccd1 _03593_ sky130_fd_sc_hd__mux2_1
XFILLER_110_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07882_ net425 _04410_ _04411_ net258 vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_86_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09621_ net797 net637 vssd1 vssd1 vccd1 vccd1 _00235_ sky130_fd_sc_hd__and2_1
X_06833_ top.findLeastValue.least2\[8\] net153 net125 _03555_ vssd1 vssd1 vccd1 vccd1
+ _02006_ sky130_fd_sc_hd__o22a_1
XFILLER_95_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06764_ net287 _03442_ vssd1 vssd1 vccd1 vccd1 _03552_ sky130_fd_sc_hd__nand2_1
X_09552_ net730 net570 vssd1 vssd1 vccd1 vccd1 _00166_ sky130_fd_sc_hd__and2_1
XFILLER_102_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_05715_ net29 net417 net359 top.WB.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1 _02343_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07299__A1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08503_ net1144 top.cb_syn.char_path_n\[73\] net225 vssd1 vssd1 vccd1 vccd1 _01591_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout255_A net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06695_ _03458_ _03474_ _03477_ _03482_ vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__a211o_1
X_09483_ net723 net563 vssd1 vssd1 vccd1 vccd1 _00097_ sky130_fd_sc_hd__and2_1
XANTENNA__07299__B2 top.findLeastValue.sum\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08434_ top.cb_syn.char_path_n\[33\] net393 net332 top.cb_syn.char_path_n\[34\] net508
+ vssd1 vssd1 vccd1 vccd1 _04793_ sky130_fd_sc_hd__a221o_1
X_05646_ top.hTree.node_reg\[38\] net310 _02725_ _02726_ vssd1 vssd1 vccd1 vccd1 _02727_
+ sky130_fd_sc_hd__a211o_1
XANTENNA__06954__S net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05849__A2 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08365_ top.cb_syn.char_path_n\[123\] top.cb_syn.char_path_n\[124\] net515 vssd1
+ vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_24_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05577_ _02667_ _02668_ net472 vssd1 vssd1 vccd1 vccd1 _02669_ sky130_fd_sc_hd__o21a_1
X_07316_ _03776_ _03780_ _03721_ vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_34_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08296_ top.cb_syn.char_path_n\[21\] net204 _04675_ vssd1 vssd1 vccd1 vccd1 _01667_
+ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout210_X net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07247_ top.findLeastValue.val1\[32\] top.findLeastValue.val2\[32\] _03887_ vssd1
+ vssd1 vccd1 vccd1 _03893_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_4_2_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_2_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_39_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout791_A net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07178_ _03821_ _03825_ _03835_ vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__o21ba_1
XANTENNA__07785__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06129_ top.cw2\[3\] _03000_ vssd1 vssd1 vccd1 vccd1 _03001_ sky130_fd_sc_hd__or2_1
XANTENNA__08420__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout331 net332 vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout320 _05088_ vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__buf_2
Xfanout353 _04073_ vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__clkbuf_2
Xfanout342 net349 vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__buf_2
Xfanout375 net377 vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_70_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout364 net367 vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__clkbuf_4
Xfanout386 net390 vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_70_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout397 net398 vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__buf_2
XFILLER_59_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09819_ net735 net575 vssd1 vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__and2_1
XFILLER_15_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_53_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ clknet_leaf_118_clk _02245_ _01067_ vssd1 vssd1 vccd1 vccd1 top.path\[43\]
+ sky130_fd_sc_hd__dfrtp_1
X_11643_ clknet_leaf_113_clk _02176_ _00998_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput17 DAT_I[23] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
Xinput28 DAT_I[4] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
X_11574_ clknet_leaf_109_clk _02122_ _00929_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput39 gpio_in[5] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__buf_1
X_10525_ net858 net698 vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__and2_1
XFILLER_108_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09203__A2 _04188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10456_ net729 net569 vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__and2_1
X_10387_ net756 net596 vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__and2_1
XFILLER_96_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09923__B net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08175__C1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11008_ clknet_leaf_12_clk _01556_ _00363_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_92_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05500_ net458 top.hTree.node_reg\[62\] net362 net422 top.hTree.node_reg\[30\] vssd1
+ vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__a32o_1
X_06480_ net1478 _03290_ vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__xor2_1
X_05431_ top.sram_interface.word_cnt\[2\] vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__inv_2
XANTENNA__05531__X _02631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08150_ top.cb_syn.char_path_n\[94\] net209 _04602_ vssd1 vssd1 vccd1 vccd1 _01740_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__05700__B2 top.WB.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07101_ _03747_ _03757_ _03758_ vssd1 vssd1 vccd1 vccd1 _03759_ sky130_fd_sc_hd__and3_1
X_05362_ top.findLeastValue.val1\[28\] vssd1 vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08081_ top.cb_syn.char_path_n\[127\] net206 net345 vssd1 vssd1 vccd1 vccd1 _04568_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09386__A net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07032_ top.findLeastValue.val1\[30\] top.findLeastValue.val2\[30\] vssd1 vssd1 vccd1
+ vccd1 _03690_ sky130_fd_sc_hd__and2_1
XANTENNA__07618__B net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06014__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10044__B net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08983_ top.WB.CPU_DAT_O\[9\] net1447 net323 vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__mux2_1
XANTENNA__09392__Y _05272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07934_ top.findLeastValue.sum\[1\] top.hTree.tree_reg\[1\] net278 vssd1 vssd1 vccd1
+ vccd1 _04453_ sky130_fd_sc_hd__mux2_1
X_07865_ top.hTree.tree_reg\[15\] top.findLeastValue.sum\[15\] net247 vssd1 vssd1
+ vccd1 vccd1 _04398_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09604_ net852 net692 vssd1 vssd1 vccd1 vccd1 _00218_ sky130_fd_sc_hd__and2_1
XANTENNA__10060__A net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07796_ net489 _04341_ vssd1 vssd1 vccd1 vccd1 _04343_ sky130_fd_sc_hd__or2_1
X_06816_ top.findLeastValue.val1\[14\] net128 net112 top.compVal\[14\] vssd1 vssd1
+ vccd1 vccd1 _02022_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_39_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout160_X net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09535_ net749 net589 vssd1 vssd1 vccd1 vccd1 _00149_ sky130_fd_sc_hd__and2_1
X_06747_ _02416_ top.findLeastValue.val2\[32\] _03529_ vssd1 vssd1 vccd1 vccd1 _03535_
+ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout637_A net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09130__A1 _02763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06678_ _02444_ top.findLeastValue.val2\[5\] top.findLeastValue.val2\[4\] _02445_
+ vssd1 vssd1 vccd1 vccd1 _03466_ sky130_fd_sc_hd__o22a_1
X_09466_ net749 net589 vssd1 vssd1 vccd1 vccd1 _00080_ sky130_fd_sc_hd__and2_1
X_08417_ top.cb_syn.char_path_n\[39\] top.cb_syn.char_path_n\[40\] net513 vssd1 vssd1
+ vccd1 vccd1 _04776_ sky130_fd_sc_hd__mux2_1
X_05629_ net1194 net138 _02712_ net174 vssd1 vssd1 vccd1 vccd1 _02379_ sky130_fd_sc_hd__a22o_1
X_09397_ net977 net241 _05274_ _05275_ vssd1 vssd1 vccd1 vccd1 _01446_ sky130_fd_sc_hd__a22o_1
X_08348_ top.cb_syn.char_path_n\[73\] net391 net330 top.cb_syn.char_path_n\[74\] net508
+ vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__a221o_1
X_08279_ top.cb_syn.char_path_n\[30\] net385 net344 top.cb_syn.char_path_n\[28\] net189
+ vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__a221o_1
XFILLER_20_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11290_ clknet_leaf_85_clk net1423 _00645_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[33\]
+ sky130_fd_sc_hd__dfrtp_1
X_10310_ net824 net664 vssd1 vssd1 vccd1 vccd1 _00924_ sky130_fd_sc_hd__and2_1
X_10241_ net828 net668 vssd1 vssd1 vccd1 vccd1 _00855_ sky130_fd_sc_hd__and2_1
XFILLER_105_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06955__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05758__B2 top.WB.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10172_ net842 net682 vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__and2_1
XANTENNA__08157__C1 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout183 net194 vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__clkbuf_2
Xfanout150 net151 vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__clkbuf_4
Xfanout161 net163 vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__clkbuf_4
Xfanout172 _02782_ vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__buf_2
XANTENNA__05616__X _02702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout194 _04566_ vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08172__A2 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06447__X _03270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11626_ clknet_leaf_36_clk _02174_ _00981_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.pulse_first
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05694__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11557_ clknet_leaf_123_clk _02105_ _00912_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_116_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold609 top.hTree.tree_reg\[16\] vssd1 vssd1 vccd1 vccd1 net1562 sky130_fd_sc_hd__dlygate4sd3_1
X_10508_ net813 net653 vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__and2_1
XFILLER_109_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_11488_ clknet_leaf_97_clk _02036_ _00843_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[28\]
+ sky130_fd_sc_hd__dfstp_2
X_10439_ net876 net716 vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_94_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05749__B2 top.WB.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05980_ net1728 top.sram_interface.init_counter\[9\] _02915_ net1100 vssd1 vssd1
+ vccd1 vccd1 _02219_ sky130_fd_sc_hd__a31o_1
XANTENNA__08699__A0 _04875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07650_ top.findLeastValue.least1\[2\] top.hTree.tree_reg\[57\] net279 vssd1 vssd1
+ vccd1 vccd1 _04225_ sky130_fd_sc_hd__mux2_1
XANTENNA__08984__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07581_ net537 _04165_ _04168_ net531 vssd1 vssd1 vccd1 vccd1 _04169_ sky130_fd_sc_hd__a22o_1
XFILLER_25_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06601_ top.compVal\[36\] _02465_ _02466_ top.compVal\[35\] vssd1 vssd1 vccd1 vccd1
+ _03390_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_36_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06532_ net466 _03316_ _03322_ vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__a21oi_1
X_09320_ _05237_ _05244_ _05249_ _05254_ net520 top.translation.index\[4\] vssd1 vssd1
+ vccd1 vccd1 _05255_ sky130_fd_sc_hd__mux4_2
X_09251_ net1124 _05210_ net296 vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_header\[6\]
+ sky130_fd_sc_hd__mux2_1
X_08202_ top.cb_syn.char_path_n\[68\] net201 _04628_ vssd1 vssd1 vccd1 vccd1 _01714_
+ sky130_fd_sc_hd__o21a_1
X_06463_ top.histogram.total\[19\] _03285_ vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_16_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09182_ _04534_ _05171_ _05172_ net474 net535 vssd1 vssd1 vccd1 vccd1 _00009_ sky130_fd_sc_hd__o32a_1
XANTENNA__06009__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05414_ top.translation.index\[3\] vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__inv_2
X_06394_ net1170 _03233_ net300 vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__mux2_1
XANTENNA__08623__B1 _04826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05345_ net1034 vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__inv_2
X_08133_ top.cb_syn.char_path_n\[103\] net382 net341 top.cb_syn.char_path_n\[101\]
+ net186 vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout120_A net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08064_ net516 _04538_ vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__or2_1
XANTENNA__07521__S1 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout218_A net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07015_ top.findLeastValue.val1\[39\] top.findLeastValue.val2\[39\] top.findLeastValue.val2\[38\]
+ top.findLeastValue.val1\[38\] vssd1 vssd1 vccd1 vccd1 _03673_ sky130_fd_sc_hd__o211a_1
XFILLER_88_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08966_ top.WB.CPU_DAT_O\[26\] net1141 net322 vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__mux2_1
XANTENNA__09055__S net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08897_ top.cb_syn.max_index\[6\] top.cb_syn.max_index\[5\] _05065_ vssd1 vssd1 vccd1
+ vccd1 _05067_ sky130_fd_sc_hd__and3_1
XANTENNA__08154__A2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout754_A net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_95_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_95_clk sky130_fd_sc_hd__clkbuf_8
X_07917_ net425 _04438_ _04439_ net258 vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__o211a_1
X_07848_ net445 net1399 net253 top.findLeastValue.sum\[19\] _04384_ vssd1 vssd1 vccd1
+ vccd1 _01824_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout542_X net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09103__A1 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07779_ top.findLeastValue.sum\[32\] top.hTree.tree_reg\[32\] net286 vssd1 vssd1
+ vccd1 vccd1 _04329_ sky130_fd_sc_hd__mux2_1
X_09518_ net732 net572 vssd1 vssd1 vccd1 vccd1 _00132_ sky130_fd_sc_hd__and2_1
X_10790_ clknet_leaf_51_clk _00030_ _00209_ vssd1 vssd1 vccd1 vccd1 top.histogram.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout807_X net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09449_ net844 net684 vssd1 vssd1 vccd1 vccd1 _00063_ sky130_fd_sc_hd__and2_1
X_11411_ clknet_leaf_99_clk _01959_ _00766_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[17\]
+ sky130_fd_sc_hd__dfstp_1
X_11342_ clknet_leaf_64_clk _01890_ _00697_ vssd1 vssd1 vccd1 vccd1 top.cw2\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__07512__S1 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11273_ clknet_leaf_106_clk net1563 _00628_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10224_ net814 net654 vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__and2_1
X_10155_ net811 net651 vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__and2_1
XANTENNA__05600__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold6 top.sram_interface.init_counter\[18\] vssd1 vssd1 vccd1 vccd1 net959 sky130_fd_sc_hd__dlygate4sd3_1
X_10086_ net874 net714 vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_86_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_86_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_47_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07353__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10988_ clknet_leaf_22_clk _01536_ _00343_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08853__B1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09929__A net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05667__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11609_ clknet_leaf_60_clk _02157_ _00964_ vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__dfrtp_1
XANTENNA__06056__C net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07503__S1 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_10_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_8
Xhold406 top.cb_syn.char_path\[98\] vssd1 vssd1 vccd1 vccd1 net1359 sky130_fd_sc_hd__dlygate4sd3_1
Xhold417 top.path\[23\] vssd1 vssd1 vccd1 vccd1 net1370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold428 top.cb_syn.char_path\[123\] vssd1 vssd1 vccd1 vccd1 net1381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold439 top.path\[53\] vssd1 vssd1 vccd1 vccd1 net1392 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08369__C1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08820_ net434 _05001_ _05002_ vssd1 vssd1 vccd1 vccd1 _05003_ sky130_fd_sc_hd__o21a_1
XANTENNA__06919__B1 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09383__B _04266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05963_ net294 _02900_ vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_77_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_clk sky130_fd_sc_hd__clkbuf_8
X_08751_ top.path\[64\] top.path\[65\] top.path\[66\] top.path\[67\] net527 net523
+ vssd1 vssd1 vccd1 vccd1 _04934_ sky130_fd_sc_hd__mux4_1
X_08682_ top.cb_syn.zeroes\[6\] _04881_ vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__nand2_1
X_05894_ top.cb_syn.wait_cycle _02553_ vssd1 vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__or2_1
XANTENNA__06147__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07702_ net490 _04264_ vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__or2_1
X_07633_ top.findLeastValue.least1\[5\] net250 _04209_ vssd1 vssd1 vccd1 vccd1 _04211_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_49_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07895__A1 top.findLeastValue.sum\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout168_A net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_07564_ top.cb_syn.h_element\[60\] top.cb_syn.h_element\[51\] _04145_ vssd1 vssd1
+ vccd1 vccd1 _04154_ sky130_fd_sc_hd__mux2_1
XANTENNA__07631__B net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07495_ top.cb_syn.char_path_n\[52\] top.cb_syn.char_path_n\[51\] top.cb_syn.char_path_n\[50\]
+ top.cb_syn.char_path_n\[49\] net400 net351 vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__mux4_1
X_09303_ top.histogram.total\[14\] top.histogram.total\[15\] net526 vssd1 vssd1 vccd1
+ vccd1 _05238_ sky130_fd_sc_hd__mux2_1
X_06515_ net1729 _03275_ net1503 vssd1 vssd1 vccd1 vccd1 _03312_ sky130_fd_sc_hd__a21oi_1
X_09234_ _02540_ _05192_ _05202_ _04913_ vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_enable
+ sky130_fd_sc_hd__a31o_1
X_06446_ top.histogram.eof_n top.histogram.state\[1\] vssd1 vssd1 vccd1 vccd1 _03269_
+ sky130_fd_sc_hd__and2b_2
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06962__S net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09165_ net450 top.histogram.state\[2\] net295 _05164_ net1600 vssd1 vssd1 vccd1
+ vccd1 _00031_ sky130_fd_sc_hd__a32o_1
XFILLER_21_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_119_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_107_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_08116_ top.cb_syn.char_path_n\[111\] net197 _04585_ vssd1 vssd1 vccd1 vccd1 _01757_
+ sky130_fd_sc_hd__o21a_1
X_06377_ _03183_ _03222_ vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__nor2_1
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09096_ net469 _02775_ _02778_ _05113_ _05115_ vssd1 vssd1 vccd1 vccd1 _05116_ sky130_fd_sc_hd__a311o_1
X_05328_ top.compVal\[13\] vssd1 vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__inv_2
X_08047_ top.cb_syn.end_cnt\[4\] net505 net507 _04540_ vssd1 vssd1 vccd1 vccd1 _04541_
+ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_116_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09021__A0 top.WB.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09998_ net836 net676 vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__and2_1
X_08949_ top.WB.CPU_DAT_O\[24\] top.cb_syn.h_element\[56\] net369 vssd1 vssd1 vccd1
+ vccd1 _01361_ sky130_fd_sc_hd__mux2_1
XFILLER_48_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_68_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_57_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09324__A1 top.header_synthesis.bit1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout757_X net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10911_ clknet_leaf_32_clk top.header_synthesis.next_zero_count\[6\] _00266_ vssd1
+ vssd1 vccd1 vccd1 top.cb_syn.zero_count\[6\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__06138__B2 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11891_ clknet_leaf_54_clk top.dut.bits_in_buf_next\[2\] _01246_ vssd1 vssd1 vccd1
+ vccd1 top.dut.bits_in_buf\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07541__B net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10842_ clknet_leaf_84_clk _01428_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_hold714_A top.histogram.sram_out\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10956__Q top.controller.fin_reg\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10773_ clknet_leaf_15_clk _01372_ _00192_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05649__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08063__A1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07497__S0 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11325_ clknet_leaf_51_clk _01873_ _00680_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.curr_index\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11256_ clknet_leaf_75_clk _01804_ _00611_ vssd1 vssd1 vccd1 vccd1 top.hTree.nullSumIndex\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09012__A0 top.WB.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08366__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11187_ clknet_leaf_27_clk _01735_ _00542_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[89\]
+ sky130_fd_sc_hd__dfrtp_1
X_10207_ net831 net671 vssd1 vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__and2_1
X_10138_ net830 net670 vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__and2_1
XANTENNA__08771__C1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_59_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_clk sky130_fd_sc_hd__clkbuf_8
X_10069_ net850 net690 vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__and2_1
XANTENNA__09931__B net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09423__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06300_ _02417_ top.hist_addr\[0\] _02942_ top.sram_interface.init_counter\[0\] _02418_
+ vssd1 vssd1 vccd1 vccd1 _03164_ sky130_fd_sc_hd__a221o_1
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07280_ _03683_ _03916_ vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__or2_1
X_06231_ top.sram_interface.init_counter\[4\] _02944_ vssd1 vssd1 vccd1 vccd1 _03099_
+ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_100_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06635__X _03424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_116_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06162_ _02963_ _03032_ _02578_ vssd1 vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__or3b_1
XANTENNA__07488__S0 _04072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_06093_ top.findLeastValue.histo_index\[7\] net549 net368 vssd1 vssd1 vccd1 vccd1
+ _02966_ sky130_fd_sc_hd__a21o_1
Xhold203 top.cb_syn.char_path\[22\] vssd1 vssd1 vccd1 vccd1 net1156 sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 top.path\[17\] vssd1 vssd1 vccd1 vccd1 net1178 sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 top.path\[27\] vssd1 vssd1 vccd1 vccd1 net1167 sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 net92 vssd1 vssd1 vccd1 vccd1 net1200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 top.cb_syn.char_path\[124\] vssd1 vssd1 vccd1 vccd1 net1189 sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 top.hTree.tree_reg\[60\] vssd1 vssd1 vccd1 vccd1 net1222 sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ net774 net614 vssd1 vssd1 vccd1 vccd1 _00535_ sky130_fd_sc_hd__and2_1
Xhold258 top.hTree.nulls\[50\] vssd1 vssd1 vccd1 vccd1 net1211 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09003__A0 top.WB.CPU_DAT_O\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout705 net706 vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__clkbuf_2
Xfanout716 net717 vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__10333__A net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout738 net739 vssd1 vssd1 vccd1 vccd1 net738 sky130_fd_sc_hd__clkbuf_2
X_09852_ net736 net576 vssd1 vssd1 vccd1 vccd1 _00466_ sky130_fd_sc_hd__and2_1
Xfanout727 net734 vssd1 vssd1 vccd1 vccd1 net727 sky130_fd_sc_hd__clkbuf_2
Xfanout749 net750 vssd1 vssd1 vccd1 vccd1 net749 sky130_fd_sc_hd__clkbuf_2
XFILLER_100_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_08803_ top.path\[22\] top.path\[23\] net524 vssd1 vssd1 vccd1 vccd1 _04986_ sky130_fd_sc_hd__mux2_1
XANTENNA__08762__C1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09783_ net762 net602 vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__and2_1
XANTENNA__06022__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08734_ _03261_ _04917_ _03251_ vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__a21boi_1
XANTENNA_fanout285_A net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10052__B net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06995_ top.findLeastValue.val1\[30\] top.findLeastValue.val1\[29\] top.findLeastValue.val1\[28\]
+ top.findLeastValue.val1\[27\] vssd1 vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__and4_1
XANTENNA__05591__A2 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05946_ top.WB.CPU_DAT_O\[9\] net1350 net306 vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__mux2_1
X_08665_ top.cb_syn.h_element\[63\] _04507_ vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__nor2_1
X_05877_ top.sram_interface.zero_cnt\[2\] top.sram_interface.zero_cnt\[1\] top.sram_interface.zero_cnt\[0\]
+ _02853_ vssd1 vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout452_A net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07868__B2 top.findLeastValue.sum\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07868__A1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08596_ net531 net534 top.cb_syn.curr_state\[5\] _02867_ vssd1 vssd1 vccd1 vccd1
+ _04818_ sky130_fd_sc_hd__or4_1
X_07616_ _02801_ _04196_ _02813_ vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__or3b_2
XFILLER_14_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07547_ net535 top.cb_syn.wait_cycle vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout717_A net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07478_ _04061_ _04068_ vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_62_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06429_ top.header_synthesis.count\[2\] _03256_ vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout505_X net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09217_ top.controller.fin_reg\[1\] top.controller.fin_reg\[2\] top.controller.fin_reg\[3\]
+ top.controller.fin_reg\[4\] vssd1 vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__or4_1
XFILLER_108_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09148_ net452 _02530_ _05155_ vssd1 vssd1 vccd1 vccd1 _05156_ sky130_fd_sc_hd__o21ai_1
X_09079_ net1679 _05098_ _05099_ top.hTree.state\[9\] vssd1 vssd1 vccd1 vccd1 _00026_
+ sky130_fd_sc_hd__a22o_1
X_11110_ clknet_leaf_6_clk _01658_ _00465_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[12\]
+ sky130_fd_sc_hd__dfrtp_2
Xhold770 top.histogram.total\[23\] vssd1 vssd1 vccd1 vccd1 net1723 sky130_fd_sc_hd__dlygate4sd3_1
X_11041_ clknet_leaf_12_clk _01589_ _00396_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[71\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08348__A2 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08753__C1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05582__A2 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input13_A DAT_I[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06531__A1 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11874_ clknet_leaf_23_clk _02390_ _01229_ vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__dfrtp_1
X_10825_ clknet_leaf_107_clk _01411_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_43_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10756_ clknet_leaf_44_clk _01355_ _00175_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10687_ clknet_leaf_120_clk _01286_ _00106_ vssd1 vssd1 vccd1 vccd1 top.path\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11308_ clknet_leaf_72_clk _01856_ _00663_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[51\]
+ sky130_fd_sc_hd__dfrtp_1
X_11239_ clknet_leaf_30_clk _01787_ _00594_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_05800_ _02803_ _02819_ vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__or2_1
X_06780_ top.findLeastValue.least1\[0\] net136 net118 net504 vssd1 vssd1 vccd1 vccd1
+ _02056_ sky130_fd_sc_hd__a22o_1
XANTENNA__05573__A2 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05731_ top.findLeastValue.histo_index\[8\] top.findLeastValue.histo_index\[7\] vssd1
+ vssd1 vccd1 vccd1 _02766_ sky130_fd_sc_hd__nor2_1
X_08450_ net1246 top.cb_syn.char_path_n\[126\] net231 vssd1 vssd1 vccd1 vccd1 _01644_
+ sky130_fd_sc_hd__mux2_1
X_05662_ _02738_ _02739_ vssd1 vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__or2_1
X_07401_ _03996_ net297 vssd1 vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__nor2_2
X_08381_ top.cb_syn.char_path_n\[103\] top.cb_syn.char_path_n\[104\] net513 vssd1
+ vssd1 vccd1 vccd1 _04740_ sky130_fd_sc_hd__mux2_1
X_05593_ top.cb_syn.char_path\[78\] net551 net542 top.cb_syn.char_path\[46\] vssd1
+ vssd1 vccd1 vccd1 _02682_ sky130_fd_sc_hd__a22o_1
X_07332_ _03729_ _03955_ vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__or2_1
XANTENNA__08275__A1 top.cb_syn.char_path_n\[32\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07263_ net268 _03902_ _03905_ net273 net1662 vssd1 vssd1 vccd1 vccd1 _01926_ sky130_fd_sc_hd__a32o_1
XANTENNA__06825__A2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06214_ top.TRN_char_index\[2\] top.TRN_char_index\[1\] top.TRN_char_index\[3\] vssd1
+ vssd1 vccd1 vccd1 _03083_ sky130_fd_sc_hd__a21o_1
XANTENNA__06017__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09002_ top.WB.CPU_DAT_O\[23\] net1437 net318 vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__mux2_1
X_07194_ top.findLeastValue.val1\[42\] top.findLeastValue.val2\[42\] vssd1 vssd1 vccd1
+ vccd1 _03852_ sky130_fd_sc_hd__or2_1
X_06145_ _02573_ _03010_ _03015_ _02574_ vssd1 vssd1 vccd1 vccd1 _03016_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_113_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06076_ top.sram_interface.init_counter\[10\] top.sram_interface.init_counter\[9\]
+ _02947_ vssd1 vssd1 vccd1 vccd1 _02950_ sky130_fd_sc_hd__nand3_1
Xfanout502 top.findLeastValue.histo_index\[2\] vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__buf_2
X_09904_ net788 net628 vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__and2_1
Xfanout513 net514 vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__clkbuf_4
Xfanout524 net526 vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__clkbuf_4
XFILLER_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout535 top.cb_syn.char_path_n\[0\] vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__buf_2
X_09835_ net777 net617 vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__and2_1
Xfanout546 net547 vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__clkbuf_4
Xfanout557 net558 vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input5_A DAT_I[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout579 net585 vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__clkbuf_2
Xfanout568 net571 vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__clkbuf_2
X_09766_ net775 net615 vssd1 vssd1 vccd1 vccd1 _00380_ sky130_fd_sc_hd__and2_1
XANTENNA__05564__A2 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06978_ top.findLeastValue.val2\[42\] top.findLeastValue.val2\[41\] top.findLeastValue.val2\[40\]
+ top.findLeastValue.val2\[39\] vssd1 vssd1 vccd1 vccd1 _03636_ sky130_fd_sc_hd__and4_1
X_08717_ net1701 _04907_ _04904_ vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__o21a_1
X_09697_ net801 net641 vssd1 vssd1 vccd1 vccd1 _00311_ sky130_fd_sc_hd__and2_1
XFILLER_66_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05929_ top.WB.CPU_DAT_O\[26\] net1169 net305 vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout834_A net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout455_X net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08648_ net1538 _04855_ vssd1 vssd1 vccd1 vccd1 _01495_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_1_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07710__A0 top.findLeastValue.least2\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08579_ _04808_ net1523 _04807_ vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__mux2_1
XANTENNA__08915__B _04187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11590_ clknet_leaf_45_clk _02138_ _00945_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10610_ net738 net578 vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__and2_1
XANTENNA__06816__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10541_ net833 net673 vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__and2_1
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10472_ net731 net571 vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__and2_1
XANTENNA__11130__Q top.cb_syn.char_path_n\[32\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07547__A net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11024_ clknet_leaf_20_clk _01572_ _00379_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05555__A2 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11857_ clknet_leaf_86_clk _02373_ _01212_ vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__dfrtp_1
X_11788_ clknet_leaf_74_clk _00023_ _01143_ vssd1 vssd1 vccd1 vccd1 top.hTree.state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10808_ clknet_leaf_83_clk _01394_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08257__A1 top.cb_syn.char_path_n\[41\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10739_ clknet_leaf_118_clk _01338_ _00158_ vssd1 vssd1 vccd1 vccd1 top.path\[115\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06807__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09937__A net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 SEL_O[0] sky130_fd_sc_hd__buf_2
XANTENNA__09301__S0 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05529__X _02629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07950_ top.findLeastValue.least1\[4\] top.findLeastValue.least2\[4\] _04462_ vssd1
+ vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__mux2_1
X_06901_ top.findLeastValue.val2\[33\] net152 net125 _03592_ vssd1 vssd1 vccd1 vccd1
+ _01975_ sky130_fd_sc_hd__o22a_1
XANTENNA__08987__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07881_ net482 _04409_ vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__or2_1
X_09620_ net797 net637 vssd1 vssd1 vccd1 vccd1 _00234_ sky130_fd_sc_hd__and2_1
XFILLER_95_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05546__A2 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06832_ _02459_ net167 _03553_ vssd1 vssd1 vccd1 vccd1 _03555_ sky130_fd_sc_hd__a21oi_1
X_06763_ net287 _03442_ vssd1 vssd1 vccd1 vccd1 _03551_ sky130_fd_sc_hd__and2_1
X_09551_ net730 net570 vssd1 vssd1 vccd1 vccd1 _00165_ sky130_fd_sc_hd__and2_1
XFILLER_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05714_ net30 net416 net309 top.WB.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1 _02344_
+ sky130_fd_sc_hd__o22a_1
X_08502_ net1110 top.cb_syn.char_path_n\[74\] net225 vssd1 vssd1 vccd1 vccd1 _01592_
+ sky130_fd_sc_hd__mux2_1
X_06694_ _02438_ top.findLeastValue.val2\[11\] _03478_ _03479_ _03481_ vssd1 vssd1
+ vccd1 vccd1 _03482_ sky130_fd_sc_hd__a2111o_1
X_09482_ net725 net565 vssd1 vssd1 vccd1 vccd1 _00096_ sky130_fd_sc_hd__and2_1
X_08433_ net438 _04781_ _04780_ net505 vssd1 vssd1 vccd1 vccd1 _04792_ sky130_fd_sc_hd__o211a_1
XFILLER_24_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05645_ top.histogram.sram_out\[6\] net363 net419 top.hTree.node_reg\[6\] vssd1 vssd1
+ vccd1 vccd1 _02726_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout150_A net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08364_ top.cb_syn.char_path_n\[125\] top.cb_syn.char_path_n\[126\] top.cb_syn.char_path_n\[127\]
+ top.cb_syn.curr_path\[127\] net515 net511 vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__mux4_1
XANTENNA__06536__A net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout248_A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05576_ top.cb_syn.char_path\[17\] net557 net312 top.cb_syn.char_path\[113\] vssd1
+ vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__a22o_1
X_07315_ net268 _03921_ _03943_ net273 net1566 vssd1 vssd1 vccd1 vccd1 _01912_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_34_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08295_ top.cb_syn.char_path_n\[22\] net383 net342 top.cb_syn.char_path_n\[20\] net187
+ vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout415_A net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07246_ net1711 net277 net272 _03892_ vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__a22o_1
X_07177_ _03824_ _03827_ _03834_ _03826_ vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__a31o_1
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06128_ top.cw2\[2\] top.cw2\[1\] top.cw2\[0\] vssd1 vssd1 vccd1 vccd1 _03000_ sky130_fd_sc_hd__and3_1
XANTENNA__08420__A1 top.cb_syn.char_path_n\[41\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06059_ net1030 net142 net137 vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__a21o_1
XANTENNA__08420__B2 top.cb_syn.char_path_n\[42\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout332 _04697_ vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__clkbuf_2
Xfanout310 net311 vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout321 net322 vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__clkbuf_4
Xfanout354 _03986_ vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__buf_2
Xfanout365 net366 vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__clkbuf_4
Xfanout343 net349 vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_70_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout387 net389 vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__buf_2
XANTENNA__05537__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout376 net377 vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__clkbuf_2
Xfanout398 _04195_ vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__clkbuf_4
XFILLER_46_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09818_ net735 net575 vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__and2_1
X_09749_ net760 net600 vssd1 vssd1 vccd1 vccd1 _00363_ sky130_fd_sc_hd__and2_1
XANTENNA__07533__C net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_53_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ clknet_leaf_116_clk _02244_ _01066_ vssd1 vssd1 vccd1 vccd1 top.path\[42\]
+ sky130_fd_sc_hd__dfrtp_1
X_11642_ clknet_leaf_102_clk _02175_ _00997_ vssd1 vssd1 vccd1 vccd1 top.hist_data_o\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_11573_ clknet_leaf_108_clk _02121_ _00928_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput18 DAT_I[24] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
X_10524_ net863 net703 vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__and2_1
Xinput29 DAT_I[5] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06733__X _03521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06880__S net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10455_ net730 net570 vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__and2_1
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10386_ net813 net653 vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__and2_1
XANTENNA__08175__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05528__A2 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11007_ clknet_leaf_13_clk _01555_ _00362_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_38_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05430_ net546 vssd1 vssd1 vccd1 vccd1 _02538_ sky130_fd_sc_hd__inv_2
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_05361_ top.findLeastValue.val1\[32\] vssd1 vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_99_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07100_ top.findLeastValue.val1\[3\] top.findLeastValue.val2\[3\] vssd1 vssd1 vccd1
+ vccd1 _03758_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_31_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08080_ net439 net389 vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__nand2_1
XANTENNA__09386__B _04261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07031_ _03686_ _03688_ vssd1 vssd1 vccd1 vccd1 _03689_ sky130_fd_sc_hd__nor2_1
XANTENNA__06091__A top.cb_syn.char_index\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08982_ top.WB.CPU_DAT_O\[10\] net1355 net323 vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__mux2_1
X_07933_ net443 net1438 net254 top.findLeastValue.sum\[2\] _04452_ vssd1 vssd1 vccd1
+ vccd1 _01807_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout198_A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07864_ top.findLeastValue.sum\[15\] top.hTree.tree_reg\[15\] net283 vssd1 vssd1
+ vccd1 vccd1 _04397_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_09603_ net804 net644 vssd1 vssd1 vccd1 vccd1 _00217_ sky130_fd_sc_hd__and2_1
XANTENNA__05519__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06815_ top.findLeastValue.val1\[15\] net129 net113 top.compVal\[15\] vssd1 vssd1
+ vccd1 vccd1 _02023_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout365_A net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10060__B net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07795_ top.findLeastValue.sum\[29\] _04341_ net397 vssd1 vssd1 vccd1 vccd1 _04342_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09534_ net750 net590 vssd1 vssd1 vccd1 vccd1 _00148_ sky130_fd_sc_hd__and2_1
X_06746_ _02410_ top.findLeastValue.val2\[39\] top.findLeastValue.val2\[35\] _02413_
+ vssd1 vssd1 vccd1 vccd1 _03534_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout153_X net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06677_ _03462_ _03463_ _03464_ vssd1 vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__a21o_1
X_09465_ net749 net589 vssd1 vssd1 vccd1 vccd1 _00079_ sky130_fd_sc_hd__and2_1
XFILLER_36_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_08416_ top.cb_syn.end_cnt\[5\] _04760_ _04774_ vssd1 vssd1 vccd1 vccd1 _04775_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_50_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05628_ top.histogram.sram_out\[9\] net363 net419 top.hTree.node_reg\[9\] _02711_
+ vssd1 vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__a221o_1
X_09396_ top.hTree.nulls\[52\] net405 net244 vssd1 vssd1 vccd1 vccd1 _05275_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout418_X net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05559_ _02652_ _02653_ net472 vssd1 vssd1 vccd1 vccd1 _02654_ sky130_fd_sc_hd__o21a_1
X_08347_ top.cb_syn.char_path_n\[75\] top.cb_syn.char_path_n\[76\] net513 vssd1 vssd1
+ vccd1 vccd1 _04706_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout320_X net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08278_ top.cb_syn.char_path_n\[30\] net207 _04666_ vssd1 vssd1 vccd1 vccd1 _01676_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_59_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07229_ _03661_ _03879_ _03660_ vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__a21bo_1
X_10240_ net834 net674 vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__and2_1
X_10171_ net832 net672 vssd1 vssd1 vccd1 vccd1 _00785_ sky130_fd_sc_hd__and2_1
Xfanout140 _02595_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_110_Right_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10251__A net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout151 net153 vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__clkbuf_2
Xfanout173 _02782_ vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout162 net163 vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__clkbuf_4
Xfanout184 net186 vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__buf_2
Xfanout195 net196 vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__buf_2
XANTENNA_hold744_A top.findLeastValue.sum\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07904__A0 top.findLeastValue.sum\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_70_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11625_ clknet_leaf_53_clk _02173_ _00980_ vssd1 vssd1 vccd1 vccd1 top.histogram.out_of_init
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_85_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05694__B2 top.WB.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08632__A1 _04826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11556_ clknet_leaf_122_clk _02104_ _00911_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10507_ net817 net657 vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__and2_1
XFILLER_109_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_11487_ clknet_leaf_97_clk _02035_ _00842_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[27\]
+ sky130_fd_sc_hd__dfstp_1
X_10438_ net873 net713 vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__and2_1
X_10369_ net855 net695 vssd1 vssd1 vccd1 vccd1 _00983_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_94_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_23_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07371__A1 top.findLeastValue.histo_index\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_1_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_1_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09360__A2 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_38_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07580_ _04149_ _04167_ vssd1 vssd1 vccd1 vccd1 _04168_ sky130_fd_sc_hd__nand2_1
X_06600_ top.compVal\[33\] _02468_ _02469_ top.compVal\[32\] vssd1 vssd1 vccd1 vccd1
+ _03389_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_36_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06531_ net466 _03321_ net957 vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__a21oi_1
X_09250_ top.header_synthesis.header\[6\] top.cb_syn.char_index\[6\] net519 vssd1
+ vssd1 vccd1 vccd1 _05210_ sky130_fd_sc_hd__mux2_1
XFILLER_61_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08201_ top.cb_syn.char_path_n\[69\] net380 net339 top.cb_syn.char_path_n\[67\] net184
+ vssd1 vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_16_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06462_ top.histogram.total\[18\] top.histogram.total\[17\] _03284_ vssd1 vssd1 vccd1
+ vccd1 _03285_ sky130_fd_sc_hd__and3_1
XANTENNA__08871__A1 top.translation.index\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09181_ _02553_ _02862_ _04893_ vssd1 vssd1 vccd1 vccd1 _05172_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_103_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05413_ top.translation.index\[4\] vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__inv_2
X_06393_ _03179_ _03232_ vssd1 vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__nor2_1
X_05344_ top.sram_interface.CB_write_counter\[0\] vssd1 vssd1 vccd1 vccd1 _02452_
+ sky130_fd_sc_hd__inv_2
X_08132_ top.cb_syn.char_path_n\[103\] net199 _04593_ vssd1 vssd1 vccd1 vccd1 _01749_
+ sky130_fd_sc_hd__o21a_1
X_08063_ net535 net246 _04552_ _04551_ net1658 vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__o32a_1
XFILLER_108_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_07014_ _03664_ _03666_ _03667_ _03671_ vssd1 vssd1 vccd1 vccd1 _03672_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout113_A net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06025__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08965_ top.WB.CPU_DAT_O\[27\] net1321 net322 vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__mux2_1
XFILLER_69_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07916_ net482 _04437_ vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__or2_1
X_08896_ top.cb_syn.max_index\[5\] _05065_ vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__nand2_1
XFILLER_68_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07847_ net428 _04382_ _04383_ net262 vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__o211a_1
XFILLER_17_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout368_X net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07778_ net443 net1422 net254 top.findLeastValue.sum\[33\] _04328_ vssd1 vssd1 vccd1
+ vccd1 _01838_ sky130_fd_sc_hd__a221o_1
X_06729_ top.compVal\[24\] _02489_ _03509_ vssd1 vssd1 vccd1 vccd1 _03517_ sky130_fd_sc_hd__o21ai_1
X_09517_ net732 net572 vssd1 vssd1 vccd1 vccd1 _00131_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout535_X net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09448_ net847 net687 vssd1 vssd1 vccd1 vccd1 _00062_ sky130_fd_sc_hd__and2_1
XFILLER_40_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09379_ net1007 _05263_ net244 vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__mux2_1
XFILLER_12_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_11410_ clknet_leaf_100_clk _01958_ _00765_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[16\]
+ sky130_fd_sc_hd__dfstp_2
X_11341_ clknet_leaf_68_clk _01889_ _00696_ vssd1 vssd1 vccd1 vccd1 top.cw2\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09100__A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10246__A net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07822__C1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11272_ clknet_leaf_79_clk _01820_ _00627_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10223_ net809 net649 vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__and2_1
XANTENNA_input43_A gpio_in[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10154_ net810 net650 vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__and2_1
X_10085_ net871 net711 vssd1 vssd1 vccd1 vccd1 _00699_ sky130_fd_sc_hd__and2_1
Xhold7 top.sram_interface.CB_read_counter vssd1 vssd1 vccd1 vccd1 net960 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07353__B2 top.findLeastValue.sum\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10987_ clknet_leaf_7_clk _01535_ _00342_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09929__B net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11608_ clknet_leaf_60_clk _02156_ _00963_ vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_96_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold407 top.cb_syn.char_path\[120\] vssd1 vssd1 vccd1 vccd1 net1360 sky130_fd_sc_hd__dlygate4sd3_1
X_11539_ clknet_leaf_2_clk _02087_ _00894_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold418 top.path\[21\] vssd1 vssd1 vccd1 vccd1 net1371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold429 top.path\[40\] vssd1 vssd1 vccd1 vccd1 net1382 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_98_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09030__A1 top.WB.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05537__X _02636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09318__C1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05962_ _02895_ _02899_ top.TRN_sram_complete vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__o21a_1
X_08750_ top.path\[68\] net411 net329 top.path\[69\] net522 vssd1 vssd1 vccd1 vccd1
+ _04933_ sky130_fd_sc_hd__o221a_1
X_08681_ _04881_ vssd1 vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__inv_2
X_05893_ top.cb_syn.wait_cycle _02553_ vssd1 vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__nor2_1
X_07701_ net491 _04266_ vssd1 vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__nand2_1
X_07632_ top.findLeastValue.least1\[5\] top.hTree.tree_reg\[60\] net280 vssd1 vssd1
+ vccd1 vccd1 _04210_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_105_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07563_ net1624 _04144_ _04152_ _04153_ vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__o22a_1
XANTENNA__07631__C net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_09302_ _05234_ _05235_ _05236_ _02523_ vssd1 vssd1 vccd1 vccd1 _05237_ sky130_fd_sc_hd__a22o_1
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07494_ _04079_ _04084_ _04069_ vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__mux2_1
XANTENNA__08844__B2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06514_ net1504 _03277_ vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__xor2_1
X_09233_ net519 _05201_ _04922_ _03251_ vssd1 vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__o211ai_1
XANTENNA_fanout230_A net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06445_ top.histogram.total\[14\] top.histogram.total\[13\] top.histogram.total\[12\]
+ vssd1 vssd1 vccd1 vccd1 _03268_ sky130_fd_sc_hd__and3_1
X_09164_ _03270_ net295 _05164_ net1690 vssd1 vssd1 vccd1 vccd1 _00030_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout328_A net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08743__B net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08115_ top.cb_syn.char_path_n\[112\] net373 net335 top.cb_syn.char_path_n\[110\]
+ net180 vssd1 vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__a221o_1
X_06376_ top.hist_data_o\[14\] _03184_ vssd1 vssd1 vccd1 vccd1 _03222_ sky130_fd_sc_hd__nor2_1
XFILLER_119_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09095_ net463 _02894_ _02899_ _02876_ net479 vssd1 vssd1 vccd1 vccd1 _05115_ sky130_fd_sc_hd__a32o_1
X_05327_ top.compVal\[14\] vssd1 vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout116_X net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08046_ net511 net516 vssd1 vssd1 vccd1 vccd1 _04540_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout697_A net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05447__X _02555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_103_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09997_ net846 net686 vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__and2_1
X_08948_ top.WB.CPU_DAT_O\[25\] top.cb_syn.h_element\[57\] _05086_ vssd1 vssd1 vccd1
+ vccd1 _01362_ sky130_fd_sc_hd__mux2_1
XANTENNA__05594__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08879_ net556 _02565_ vssd1 vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__nor2_1
XANTENNA__09324__A2 top.header_synthesis.enable vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10910_ clknet_leaf_32_clk top.header_synthesis.next_zero_count\[5\] _00265_ vssd1
+ vssd1 vccd1 vccd1 top.cb_syn.zero_count\[5\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__06138__A2 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11890_ clknet_leaf_54_clk top.dut.bits_in_buf_next\[1\] _01245_ vssd1 vssd1 vccd1
+ vccd1 top.dut.bits_in_buf\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10841_ clknet_leaf_78_clk _01427_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_80_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10772_ clknet_leaf_15_clk _01371_ _00191_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08835__A1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06846__B1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07497__S1 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11324_ clknet_leaf_51_clk _01872_ _00679_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.curr_index\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11255_ clknet_leaf_75_clk _01803_ _00610_ vssd1 vssd1 vccd1 vccd1 top.hTree.nullSumIndex\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10206_ net830 net670 vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__and2_1
XANTENNA__07285__A _03782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11186_ clknet_leaf_19_clk _01734_ _00541_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[88\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__05585__B1 _02674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10137_ net831 net671 vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__and2_1
X_10068_ net850 net690 vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08826__A1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06837__A0 top.findLeastValue.least1\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06230_ top.hist_addr\[4\] _03021_ vssd1 vssd1 vccd1 vccd1 _03098_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_100_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06301__A2 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06161_ top.cb_syn.char_index\[5\] _02962_ vssd1 vssd1 vccd1 vccd1 _03032_ sky130_fd_sc_hd__nor2_1
XANTENNA__07488__S1 _04071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06092_ _02480_ _02481_ vssd1 vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__nor2_1
Xhold204 top.histogram.sram_out\[31\] vssd1 vssd1 vccd1 vccd1 net1157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 top.cb_syn.char_path\[19\] vssd1 vssd1 vccd1 vccd1 net1179 sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 net79 vssd1 vssd1 vccd1 vccd1 net1168 sky130_fd_sc_hd__dlygate4sd3_1
X_09920_ net743 net583 vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__and2_1
Xhold259 top.path\[3\] vssd1 vssd1 vccd1 vccd1 net1212 sky130_fd_sc_hd__dlygate4sd3_1
Xhold248 top.path\[0\] vssd1 vssd1 vccd1 vccd1 net1201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 top.cb_syn.char_path\[72\] vssd1 vssd1 vccd1 vccd1 net1190 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_98_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xfanout706 net717 vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__clkbuf_2
Xfanout717 net718 vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__clkbuf_4
XFILLER_98_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__10333__B net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout739 net745 vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__clkbuf_2
Xfanout728 net731 vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__clkbuf_2
X_09851_ net737 net577 vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__and2_1
XFILLER_105_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__05576__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09782_ net758 net598 vssd1 vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__and2_1
X_08802_ top.path\[17\] net326 _04984_ vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__o21a_1
X_06994_ top.findLeastValue.val1\[26\] net496 top.findLeastValue.val1\[24\] top.findLeastValue.val1\[23\]
+ vssd1 vssd1 vccd1 vccd1 _03652_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08733_ top.header_synthesis.enable top.header_synthesis.write_char_path top.header_synthesis.char_added
+ vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__and3_1
X_05945_ top.WB.CPU_DAT_O\[10\] net1218 net306 vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__mux2_1
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout278_A _04198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08664_ _04129_ _04866_ vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__nor2_1
X_05876_ top.sram_interface.zero_cnt\[2\] _02449_ top.sram_interface.zero_cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__o21ai_1
XFILLER_81_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08595_ _04557_ _04558_ _04560_ _04816_ vssd1 vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__or4b_1
X_07615_ _02795_ _02799_ vssd1 vssd1 vccd1 vccd1 _04196_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout445_A net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07546_ top.cb_syn.curr_state\[0\] _04136_ vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__or2_1
XANTENNA__08817__A1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07477_ _04048_ _04060_ vssd1 vssd1 vccd1 vccd1 _04068_ sky130_fd_sc_hd__nand2_1
X_09216_ _05188_ _05189_ vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout233_X net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout612_A net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06428_ top.header_synthesis.count\[1\] top.header_synthesis.count\[0\] _03245_ vssd1
+ vssd1 vccd1 vccd1 _03256_ sky130_fd_sc_hd__and3_1
XANTENNA__05500__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09147_ top.sram_interface.TRN_counter\[2\] top.sram_interface.TRN_counter\[1\] top.sram_interface.TRN_counter\[0\]
+ net465 vssd1 vssd1 vccd1 vccd1 _05155_ sky130_fd_sc_hd__or4b_1
XANTENNA_fanout400_X net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06359_ net1214 _03211_ net302 vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__mux2_1
XFILLER_107_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09078_ _02820_ net257 vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__or2_1
XANTENNA__09585__A net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07253__B1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_15_Left_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08029_ top.cb_syn.count\[1\] top.cb_syn.count\[0\] vssd1 vssd1 vccd1 vccd1 _04526_
+ sky130_fd_sc_hd__or2_1
Xhold771 top.findLeastValue.sum\[30\] vssd1 vssd1 vccd1 vccd1 net1724 sky130_fd_sc_hd__dlygate4sd3_1
Xhold760 top.compVal\[9\] vssd1 vssd1 vccd1 vccd1 net1713 sky130_fd_sc_hd__dlygate4sd3_1
X_11040_ clknet_leaf_12_clk _01588_ _00395_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[70\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_76_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_24_Left_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10967__Q top.cb_syn.char_index\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11873_ clknet_leaf_23_clk _02389_ _01228_ vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__dfrtp_1
XFILLER_60_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10824_ clknet_leaf_107_clk _01410_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_43_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06819__B1 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10755_ clknet_leaf_47_clk _01354_ _00174_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_10686_ clknet_leaf_120_clk _01285_ _00105_ vssd1 vssd1 vccd1 vccd1 top.path\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09233__A1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_33_Left_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06047__A1 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07244__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11307_ clknet_leaf_84_clk _01855_ _00662_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08992__A0 top.WB.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11238_ clknet_leaf_30_clk _01786_ _00593_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05558__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11169_ clknet_leaf_11_clk _01717_ _00524_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[71\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_42_Left_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05730_ top.findLeastValue.alternator_timer\[2\] _02764_ _02763_ top.findLeastValue.alternator_timer\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__a211oi_1
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05661_ top.cb_syn.char_path\[3\] net558 net316 top.cb_syn.char_path\[99\] vssd1
+ vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__a22o_1
X_07400_ top.dut.bits_in_buf_next\[2\] net297 vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__or2_2
X_08380_ net510 _04737_ _04738_ vssd1 vssd1 vccd1 vccd1 _04739_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07889__S net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05730__B1 _02763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05592_ net1168 net138 _02681_ net174 vssd1 vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__a22o_1
X_07331_ _03734_ _03954_ _03732_ vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_0_clk_X clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09389__B _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_51_Left_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07262_ _03694_ _03901_ vssd1 vssd1 vccd1 vccd1 _03905_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_21_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06213_ top.TRN_char_index\[3\] _02974_ vssd1 vssd1 vccd1 vccd1 _03082_ sky130_fd_sc_hd__nor2_1
X_09001_ top.WB.CPU_DAT_O\[24\] net1414 net317 vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__mux2_1
X_07193_ top.findLeastValue.val1\[42\] top.findLeastValue.val2\[42\] vssd1 vssd1 vccd1
+ vccd1 _03851_ sky130_fd_sc_hd__nand2_1
X_06144_ net497 net549 _03014_ vssd1 vssd1 vccd1 vccd1 _03015_ sky130_fd_sc_hd__and3_1
XANTENNA__08513__S net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08983__A0 top.WB.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06075_ net1049 net144 net137 _02949_ vssd1 vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__a211o_1
XANTENNA__07637__B net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout503 top.findLeastValue.histo_index\[1\] vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__buf_2
X_09903_ net789 net629 vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__and2_1
Xfanout514 top.cb_syn.end_cnt\[0\] vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_4_9_0_clk_X clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout536 top.cb_syn.curr_state\[4\] vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__buf_2
X_09834_ net777 net617 vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__and2_1
Xfanout547 top.sram_interface.word_cnt\[10\] vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__buf_2
XANTENNA__05549__B1 _02644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_60_Left_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout525 net526 vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__buf_2
XFILLER_86_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07653__A net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout558 net560 vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__clkbuf_4
Xfanout569 net571 vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08749__A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout562_A top.sram_interface.word_cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09765_ net773 net613 vssd1 vssd1 vccd1 vccd1 _00379_ sky130_fd_sc_hd__and2_1
X_06977_ _03631_ _03632_ _03633_ _03634_ vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__and4_1
X_08716_ _04898_ _04902_ vssd1 vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__nor2_1
X_09696_ net794 net634 vssd1 vssd1 vccd1 vccd1 _00310_ sky130_fd_sc_hd__and2_1
X_05928_ top.WB.CPU_DAT_O\[27\] net1376 net305 vssd1 vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__mux2_1
XFILLER_26_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08647_ _04845_ _04847_ net193 vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__a21o_1
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout350_X net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05859_ top.compVal\[8\] net170 net156 top.WB.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1
+ _02283_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_1_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout448_X net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07799__S net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08578_ top.cb_syn.h_element\[62\] top.cb_syn.h_element\[53\] net532 vssd1 vssd1
+ vccd1 vccd1 _04808_ sky130_fd_sc_hd__mux2_1
XANTENNA__05901__A _02875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10519__A net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07529_ _04108_ _04119_ _04067_ vssd1 vssd1 vccd1 vccd1 _04120_ sky130_fd_sc_hd__mux2_1
X_10540_ net763 net603 vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__and2_1
X_10471_ net728 net568 vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__and2_1
XANTENNA__06029__A1 top.WB.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07777__A1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08974__A0 top.WB.CPU_DAT_O\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xhold590 top.hTree.tree_reg\[37\] vssd1 vssd1 vccd1 vccd1 net1543 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11023_ clknet_leaf_20_clk _01571_ _00378_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06878__S net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11856_ clknet_leaf_70_clk _02372_ _01211_ vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__dfrtp_1
XANTENNA__05712__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10807_ clknet_leaf_51_clk _01393_ _00226_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.max_index\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_11787_ clknet_leaf_75_clk _00022_ _01142_ vssd1 vssd1 vccd1 vccd1 top.hTree.state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10738_ clknet_leaf_118_clk _01337_ _00157_ vssd1 vssd1 vccd1 vccd1 top.path\[114\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09937__B net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10669_ clknet_leaf_119_clk _01268_ _00088_ vssd1 vssd1 vccd1 vccd1 top.path\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 SEL_O[1] sky130_fd_sc_hd__buf_2
XANTENNA__05491__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08965__A0 top.WB.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09301__S1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06900_ top.compVal\[33\] top.findLeastValue.val1\[33\] net167 vssd1 vssd1 vccd1
+ vccd1 _03592_ sky130_fd_sc_hd__mux2_1
X_07880_ top.hTree.tree_reg\[12\] top.findLeastValue.sum\[12\] net247 vssd1 vssd1
+ vccd1 vccd1 _04410_ sky130_fd_sc_hd__mux2_1
X_06831_ net1660 net134 net119 net413 vssd1 vssd1 vccd1 vccd1 _02007_ sky130_fd_sc_hd__a22o_1
XFILLER_83_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06089__A top.cb_syn.char_index\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06762_ net287 net152 vssd1 vssd1 vccd1 vccd1 _03550_ sky130_fd_sc_hd__nand2_1
XANTENNA__05951__A0 top.WB.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09550_ net730 net570 vssd1 vssd1 vccd1 vccd1 _00164_ sky130_fd_sc_hd__and2_1
XANTENNA__07940__A1 top.findLeastValue.sum\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07760__X _04314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05713_ net31 net416 net309 top.WB.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1 _02345_
+ sky130_fd_sc_hd__o22a_1
X_09481_ net725 net565 vssd1 vssd1 vccd1 vccd1 _00095_ sky130_fd_sc_hd__and2_1
X_08501_ net1316 top.cb_syn.char_path_n\[75\] net221 vssd1 vssd1 vccd1 vccd1 _01593_
+ sky130_fd_sc_hd__mux2_1
X_08432_ _02505_ _04786_ _04788_ _04790_ net506 vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__o221a_1
X_06693_ _02436_ top.findLeastValue.val2\[13\] top.findLeastValue.val2\[12\] _02437_
+ vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__a22o_1
XFILLER_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05644_ _02723_ _02724_ net473 vssd1 vssd1 vccd1 vccd1 _02725_ sky130_fd_sc_hd__o21a_1
XANTENNA__05703__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout143_A net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08363_ top.cb_syn.end_cnt\[5\] _04718_ _04721_ vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__or3b_1
X_05575_ top.cb_syn.char_path\[81\] net551 net543 top.cb_syn.char_path\[49\] vssd1
+ vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__a22o_1
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08294_ top.cb_syn.char_path_n\[22\] net204 _04674_ vssd1 vssd1 vccd1 vccd1 _01668_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_34_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07314_ _03782_ _03799_ vssd1 vssd1 vccd1 vccd1 _03943_ sky130_fd_sc_hd__nand2_1
X_07245_ _03824_ _03888_ vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__xor2_1
XANTENNA__11231__Q top.cb_syn.end_cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout310_A net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout408_A _02788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08956__A0 top.WB.CPU_DAT_O\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07176_ top.findLeastValue.val1\[33\] top.findLeastValue.val2\[33\] _03833_ vssd1
+ vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__o21a_1
XFILLER_117_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06127_ top.cw2\[1\] top.cw2\[0\] vssd1 vssd1 vccd1 vccd1 _02999_ sky130_fd_sc_hd__nand2_1
XANTENNA__07000__X _03658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08420__A2 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06058_ net1031 net144 net137 vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout398_X net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout311 _02690_ vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__clkbuf_2
Xfanout300 net303 vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout322 net323 vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__buf_2
Xfanout366 net367 vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__clkbuf_2
Xfanout344 net345 vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__buf_2
Xfanout333 net334 vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__buf_2
Xfanout355 net356 vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06195__B1 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xfanout388 net389 vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__buf_2
Xfanout377 net390 vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_70_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout399 net400 vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__buf_4
X_09817_ net741 net581 vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__and2_1
X_09748_ net765 net605 vssd1 vssd1 vccd1 vccd1 _00362_ sky130_fd_sc_hd__and2_1
XANTENNA__05942__A0 top.WB.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09679_ net783 net623 vssd1 vssd1 vccd1 vccd1 _00293_ sky130_fd_sc_hd__and2_1
X_11710_ clknet_leaf_117_clk _02243_ _01065_ vssd1 vssd1 vccd1 vccd1 top.path\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08418__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11641_ clknet_leaf_56_clk top.dut.bit_buf_next\[13\] _00996_ vssd1 vssd1 vccd1 vccd1
+ top.dut.bit_buf\[13\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10249__A net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11572_ clknet_leaf_113_clk _02120_ _00927_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10523_ net861 net701 vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__and2_1
Xinput19 DAT_I[25] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08947__A0 top.WB.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10454_ net748 net588 vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__and2_1
X_10385_ net812 net652 vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__and2_1
XFILLER_97_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11006_ clknet_leaf_14_clk _01554_ _00361_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05933__A0 top.WB.CPU_DAT_O\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_11839_ clknet_leaf_117_clk _02355_ _01194_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05360_ top.findLeastValue.val1\[33\] vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_99_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07030_ top.findLeastValue.val1\[31\] top.findLeastValue.val2\[31\] vssd1 vssd1 vccd1
+ vccd1 _03688_ sky130_fd_sc_hd__nor2_1
XANTENNA__08938__A0 top.WB.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06413__A1 top.histogram.sram_out\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07755__X _04310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08981_ top.WB.CPU_DAT_O\[11\] net1244 net323 vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__mux2_1
X_07932_ net429 _04450_ _04451_ net260 vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__o211a_1
XANTENNA__06177__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07863_ net441 net1562 net252 top.findLeastValue.sum\[16\] _04396_ vssd1 vssd1 vccd1
+ vccd1 _01821_ sky130_fd_sc_hd__a221o_1
X_09602_ net856 net696 vssd1 vssd1 vccd1 vccd1 _00216_ sky130_fd_sc_hd__and2_1
X_06814_ top.findLeastValue.val1\[16\] net128 net112 net1628 vssd1 vssd1 vccd1 vccd1
+ _02024_ sky130_fd_sc_hd__o22a_1
XANTENNA__05924__A0 top.WB.CPU_DAT_O\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07913__A1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07794_ top.findLeastValue.sum\[29\] top.hTree.tree_reg\[29\] net280 vssd1 vssd1
+ vccd1 vccd1 _04341_ sky130_fd_sc_hd__mux2_1
X_09533_ net750 net590 vssd1 vssd1 vccd1 vccd1 _00147_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_39_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout358_A _02926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06745_ _02410_ top.findLeastValue.val2\[39\] top.findLeastValue.val2\[38\] _02411_
+ vssd1 vssd1 vccd1 vccd1 _03533_ sky130_fd_sc_hd__o22a_1
XFILLER_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout260_A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06676_ _02445_ top.findLeastValue.val2\[4\] top.findLeastValue.val2\[3\] _02446_
+ vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__a22o_1
X_09464_ net754 net594 vssd1 vssd1 vccd1 vccd1 _00078_ sky130_fd_sc_hd__and2_1
X_08415_ net507 _04763_ _04766_ _04773_ top.cb_syn.end_cnt\[4\] vssd1 vssd1 vccd1
+ vccd1 _04774_ sky130_fd_sc_hd__o311a_1
X_09395_ net405 _04246_ vssd1 vssd1 vccd1 vccd1 _05274_ sky130_fd_sc_hd__nand2_1
X_05627_ top.hTree.node_reg\[41\] net310 _02710_ net473 vssd1 vssd1 vccd1 vccd1 _02711_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09858__A net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08346_ top.cb_syn.char_path_n\[77\] top.cb_syn.char_path_n\[78\] top.cb_syn.char_path_n\[79\]
+ top.cb_syn.char_path_n\[80\] net514 net510 vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__mux4_1
XFILLER_51_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout525_A net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05558_ top.cb_syn.char_path\[20\] net558 net313 top.cb_syn.char_path\[116\] vssd1
+ vssd1 vccd1 vccd1 _02653_ sky130_fd_sc_hd__a22o_1
XFILLER_20_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_05489_ net453 _02592_ net160 vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__a21o_1
X_08277_ top.cb_syn.char_path_n\[31\] net386 net345 top.cb_syn.char_path_n\[29\] net190
+ vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout313_X net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07228_ _03660_ _03661_ _03879_ vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__nand3b_1
XANTENNA__08929__A0 top.WB.CPU_DAT_O\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07159_ _03704_ _03782_ _03808_ vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__or3_2
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout682_X net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10170_ net842 net682 vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__and2_1
XANTENNA__06955__A2 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xfanout130 net131 vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__clkbuf_4
Xfanout141 net143 vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__buf_2
Xfanout152 net153 vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09354__B1 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout174 net176 vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__buf_4
Xfanout163 _03423_ vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10251__B net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout185 net186 vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout196 net211 vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__clkbuf_4
XFILLER_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09121__A3 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11624_ clknet_leaf_54_clk _02172_ _00979_ vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08672__A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Left_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05694__A2 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11555_ clknet_leaf_122_clk _02103_ _00910_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10506_ net812 net652 vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__and2_1
X_11486_ clknet_leaf_103_clk _02034_ _00841_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[26\]
+ sky130_fd_sc_hd__dfstp_1
X_10437_ net875 net715 vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__and2_1
XFILLER_7_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10368_ net853 net693 vssd1 vssd1 vccd1 vccd1 _00982_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_94_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10299_ net724 net564 vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__and2_1
XANTENNA__07371__A2 _03553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06530_ top.histogram.eof_n top.dut.out_valid _03319_ vssd1 vssd1 vccd1 vccd1 _03321_
+ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06461_ top.histogram.total\[16\] top.histogram.total\[15\] _03268_ _03281_ vssd1
+ vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__and4_1
XANTENNA__10885__Q top.translation.index\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08200_ top.cb_syn.char_path_n\[69\] net201 _04627_ vssd1 vssd1 vccd1 vccd1 _01715_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_16_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05412_ top.translation.index\[5\] vssd1 vssd1 vccd1 vccd1 _02520_ sky130_fd_sc_hd__inv_2
X_09180_ _02528_ _04554_ vssd1 vssd1 vccd1 vccd1 _05171_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_103_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06392_ top.hist_data_o\[8\] _03178_ vssd1 vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__nor2_1
X_05343_ top.sram_interface.CB_write_counter\[1\] vssd1 vssd1 vccd1 vccd1 _02451_
+ sky130_fd_sc_hd__inv_2
X_08131_ top.cb_syn.char_path_n\[104\] net378 net341 top.cb_syn.char_path_n\[102\]
+ net182 vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__a221o_1
X_08062_ top.cb_syn.end_cnt\[2\] net392 vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07013_ _03669_ _03670_ vssd1 vssd1 vccd1 vccd1 _03671_ sky130_fd_sc_hd__nand2_1
XFILLER_102_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08964_ top.WB.CPU_DAT_O\[28\] net1336 net321 vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__mux2_1
XANTENNA__05446__A top.CB_write_complete vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07915_ top.hTree.tree_reg\[5\] top.findLeastValue.sum\[5\] net247 vssd1 vssd1 vccd1
+ vccd1 _04438_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout475_A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08895_ top.cb_syn.max_index\[4\] top.cb_syn.max_index\[3\] top.cb_syn.max_index\[2\]
+ top.cb_syn.max_index\[1\] vssd1 vssd1 vccd1 vccd1 _05065_ sky130_fd_sc_hd__and4_1
X_07846_ net485 _04381_ vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout642_A net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07777_ net430 _04326_ _04327_ net266 vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__o211a_1
X_09516_ net725 net565 vssd1 vssd1 vccd1 vccd1 _00130_ sky130_fd_sc_hd__and2_1
X_06728_ _03505_ _03508_ _03515_ vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__or3b_1
X_09447_ net847 net687 vssd1 vssd1 vccd1 vccd1 _00061_ sky130_fd_sc_hd__and2_1
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout430_X net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout528_X net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06659_ _02407_ top.findLeastValue.val2\[44\] vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__nand2_1
X_09378_ top.hTree.nulls\[46\] _04275_ net406 vssd1 vssd1 vccd1 vccd1 _05263_ sky130_fd_sc_hd__mux2_1
XFILLER_24_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05676__A2 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10527__A net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08329_ top.cb_syn.char_path_n\[5\] net379 net338 top.cb_syn.char_path_n\[3\] net183
+ vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__a221o_1
X_11340_ clknet_leaf_67_clk _01888_ _00695_ vssd1 vssd1 vccd1 vccd1 top.cw2\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10246__B net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11271_ clknet_leaf_106_clk _01819_ _00626_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10222_ net808 net648 vssd1 vssd1 vccd1 vccd1 _00836_ sky130_fd_sc_hd__and2_1
XFILLER_106_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10153_ net810 net650 vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__and2_1
XANTENNA__05600__A2 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10084_ net871 net711 vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__and2_1
Xhold8 _02311_ vssd1 vssd1 vccd1 vccd1 net961 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_87_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input36_A gpio_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07889__A0 top.findLeastValue.sum\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06886__S net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07353__A2 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10986_ clknet_leaf_7_clk _01534_ _00341_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_70_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05667__A2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11607_ clknet_leaf_61_clk _02155_ _00962_ vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__dfrtp_1
XFILLER_30_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__07813__B1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold408 top.path\[6\] vssd1 vssd1 vccd1 vccd1 net1361 sky130_fd_sc_hd__dlygate4sd3_1
X_11538_ clknet_leaf_0_clk _02086_ _00893_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_109_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08369__A1 _02506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11469_ clknet_leaf_96_clk _02017_ _00824_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[9\]
+ sky130_fd_sc_hd__dfstp_1
Xhold419 top.path\[89\] vssd1 vssd1 vccd1 vccd1 net1372 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10172__A net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09318__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07700_ _02478_ net397 _04265_ vssd1 vssd1 vccd1 vccd1 _04266_ sky130_fd_sc_hd__o21a_1
X_05961_ top.translation.totalEn _02791_ _02897_ _02898_ vssd1 vssd1 vccd1 vccd1 _02899_
+ sky130_fd_sc_hd__a211o_2
X_08680_ _02511_ _04880_ vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__nor2_1
X_05892_ top.cb_syn.h_element\[63\] _02866_ vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__and2_1
XANTENNA__05553__X _02649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07631_ top.hTree.tree_reg\[60\] net397 net286 vssd1 vssd1 vccd1 vccd1 _04209_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_105_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07562_ top.cb_syn.max_index\[7\] _04135_ _04144_ vssd1 vssd1 vccd1 vccd1 _04153_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_80_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06513_ _03279_ _03311_ vssd1 vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__nor2_1
X_09301_ top.histogram.total\[0\] top.histogram.total\[1\] top.histogram.total\[2\]
+ top.histogram.total\[3\] net526 net523 vssd1 vssd1 vccd1 vccd1 _05236_ sky130_fd_sc_hd__mux4_1
XFILLER_34_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07493_ _04080_ _04081_ _04082_ _04083_ _04072_ _04071_ vssd1 vssd1 vccd1 vccd1 _04084_
+ sky130_fd_sc_hd__mux4_1
X_06444_ top.header_synthesis.count\[0\] _03245_ _03267_ vssd1 vssd1 vccd1 vccd1 _02107_
+ sky130_fd_sc_hd__o21a_1
X_09232_ top.header_synthesis.write_zeroes _05200_ top.header_synthesis.enable vssd1
+ vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__a21bo_1
XANTENNA__08516__S net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09163_ net453 net295 net449 vssd1 vssd1 vccd1 vccd1 _05164_ sky130_fd_sc_hd__a21o_1
X_06375_ net1258 _03221_ net301 vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout223_A net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08114_ top.cb_syn.char_path_n\[112\] net197 _04584_ vssd1 vssd1 vccd1 vccd1 _01758_
+ sky130_fd_sc_hd__o21a_1
X_05326_ top.compVal\[15\] vssd1 vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__inv_2
X_09094_ net463 _02894_ vssd1 vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__nand2_1
X_08045_ net512 net515 vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_116_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05728__X _02763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09996_ net848 net688 vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__and2_1
XFILLER_76_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout857_A net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08947_ top.WB.CPU_DAT_O\[26\] top.cb_syn.h_element\[58\] _05086_ vssd1 vssd1 vccd1
+ vccd1 _01363_ sky130_fd_sc_hd__mux2_1
XFILLER_57_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06791__B1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_84_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08878_ _05041_ _05042_ net527 vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__mux2_1
XFILLER_84_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07829_ top.findLeastValue.sum\[22\] top.hTree.tree_reg\[22\] net285 vssd1 vssd1
+ vccd1 vccd1 _04369_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_88_Left_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10840_ clknet_leaf_80_clk _01426_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_80_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10771_ clknet_leaf_14_clk _01370_ _00190_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_99_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05649__A2 top.sram_interface.word_cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_22_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_97_Left_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11323_ clknet_leaf_66_clk _01871_ _00678_ vssd1 vssd1 vccd1 vccd1 top.controller.fin_FINISHED
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_0_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_0_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_37_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11254_ clknet_leaf_75_clk _01802_ _00609_ vssd1 vssd1 vccd1 vccd1 top.hTree.nullSumIndex\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10205_ net830 net670 vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__and2_1
X_11185_ clknet_leaf_19_clk _01733_ _00540_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[87\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06782__B1 _03553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10136_ net831 net671 vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__and2_1
X_10067_ net850 net690 vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__and2_1
XFILLER_47_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkload1_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10969_ clknet_leaf_40_clk _01517_ _00324_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_index\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06837__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06160_ top.cb_syn.char_index\[5\] _02960_ _02579_ vssd1 vssd1 vccd1 vccd1 _03031_
+ sky130_fd_sc_hd__o21ai_1
X_06091_ top.cb_syn.char_index\[6\] _02963_ vssd1 vssd1 vccd1 vccd1 _02964_ sky130_fd_sc_hd__nand2_1
Xhold205 top.cb_syn.char_path\[80\] vssd1 vssd1 vccd1 vccd1 net1158 sky130_fd_sc_hd__dlygate4sd3_1
Xhold216 top.path\[58\] vssd1 vssd1 vccd1 vccd1 net1169 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06651__Y _03440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold249 top.path\[54\] vssd1 vssd1 vccd1 vccd1 net1202 sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 net74 vssd1 vssd1 vccd1 vccd1 net1191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 top.cb_syn.char_path\[13\] vssd1 vssd1 vccd1 vccd1 net1180 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout718 net719 vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__buf_2
Xfanout707 net717 vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__clkbuf_2
Xfanout729 net731 vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__clkbuf_2
X_09850_ net741 net581 vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__and2_1
XFILLER_85_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06773__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09781_ net762 net602 vssd1 vssd1 vccd1 vccd1 _00395_ sky130_fd_sc_hd__and2_1
X_08801_ top.path\[16\] net408 _04983_ net432 net436 vssd1 vssd1 vccd1 vccd1 _04984_
+ sky130_fd_sc_hd__o221a_1
X_06993_ _03647_ _03648_ _03649_ _03650_ vssd1 vssd1 vccd1 vccd1 _03651_ sky130_fd_sc_hd__and4_1
X_08732_ _04913_ _04915_ vssd1 vssd1 vccd1 vccd1 _04916_ sky130_fd_sc_hd__nand2_1
X_05944_ top.WB.CPU_DAT_O\[11\] net1305 net306 vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__mux2_1
X_08663_ _04126_ _04508_ vssd1 vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__and2b_1
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05875_ net550 net468 vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout173_A _02782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08594_ net531 net534 top.cb_syn.curr_state\[5\] net540 vssd1 vssd1 vccd1 vccd1 _04816_
+ sky130_fd_sc_hd__or4_1
X_07614_ top.hTree.write_HT_fin top.hTree.closing vssd1 vssd1 vccd1 vccd1 _04195_
+ sky130_fd_sc_hd__or2_1
X_07545_ net534 net539 _04134_ vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__or3_2
XANTENNA_fanout340_A net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07476_ _04062_ _04066_ vssd1 vssd1 vccd1 vccd1 _04067_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_4_5_0_clk_X clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout438_A _02505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06427_ net1565 _03254_ _03255_ vssd1 vssd1 vccd1 vccd1 _02112_ sky130_fd_sc_hd__a21o_1
X_09215_ top.controller.fin_reg\[1\] top.controller.fin_reg\[2\] top.controller.fin_reg\[4\]
+ top.controller.fin_reg\[3\] vssd1 vssd1 vccd1 vccd1 _05189_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_62_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05500__A1 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09146_ top.sram_interface.CB_write_counter\[1\] top.sram_interface.CB_write_counter\[0\]
+ net479 _05139_ vssd1 vssd1 vccd1 vccd1 _05154_ sky130_fd_sc_hd__a31o_1
X_06358_ _03189_ _03210_ vssd1 vssd1 vccd1 vccd1 _03211_ sky130_fd_sc_hd__nor2_1
X_05309_ net495 vssd1 vssd1 vccd1 vccd1 _02417_ sky130_fd_sc_hd__inv_2
X_06289_ net549 _02573_ _03150_ _03152_ vssd1 vssd1 vccd1 vccd1 _03154_ sky130_fd_sc_hd__a31o_1
X_09077_ _02820_ net257 vssd1 vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__nor2_1
XANTENNA__09585__B net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08028_ _04512_ _04520_ _04525_ _04509_ net1663 vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__a32o_1
XFILLER_116_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold772 top.findLeastValue.sum\[20\] vssd1 vssd1 vccd1 vccd1 net1725 sky130_fd_sc_hd__dlygate4sd3_1
Xhold761 top.findLeastValue.sum\[11\] vssd1 vssd1 vccd1 vccd1 net1714 sky130_fd_sc_hd__dlygate4sd3_1
Xhold750 top.findLeastValue.sum\[43\] vssd1 vssd1 vccd1 vccd1 net1703 sky130_fd_sc_hd__dlygate4sd3_1
X_09979_ net781 net621 vssd1 vssd1 vccd1 vccd1 _00593_ sky130_fd_sc_hd__and2_1
XANTENNA__08753__B2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11872_ clknet_leaf_23_clk _02388_ _01227_ vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__dfrtp_1
XFILLER_44_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_105_Right_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10823_ clknet_leaf_107_clk _01409_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_43_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08808__A2 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_118_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_118_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08364__S0 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10754_ clknet_leaf_44_clk _01353_ _00173_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10685_ clknet_leaf_120_clk _01284_ _00104_ vssd1 vssd1 vccd1 vccd1 top.path\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07244__A1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11306_ clknet_leaf_71_clk _01854_ _00661_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[49\]
+ sky130_fd_sc_hd__dfrtp_1
X_11237_ clknet_leaf_30_clk _01785_ _00592_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11168_ clknet_leaf_13_clk _01716_ _00523_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[70\]
+ sky130_fd_sc_hd__dfrtp_2
X_10119_ net821 net661 vssd1 vssd1 vccd1 vccd1 _00733_ sky130_fd_sc_hd__and2_1
X_11099_ clknet_leaf_42_clk _01647_ _00454_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_05660_ top.cb_syn.char_path\[67\] net552 net543 top.cb_syn.char_path\[35\] vssd1
+ vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__a22o_1
X_05591_ top.histogram.sram_out\[15\] net364 _02679_ _02680_ vssd1 vssd1 vccd1 vccd1
+ _02681_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_109_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_109_clk
+ sky130_fd_sc_hd__clkbuf_8
X_07330_ top.findLeastValue.val1\[8\] top.findLeastValue.val2\[8\] _03775_ vssd1 vssd1
+ vccd1 vccd1 _03954_ sky130_fd_sc_hd__a21bo_1
X_07261_ net268 _03903_ _03904_ net273 net1611 vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__a32o_1
X_09000_ top.WB.CPU_DAT_O\[25\] net1372 net317 vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__mux2_1
X_06212_ top.cb_syn.char_index\[3\] top.cb_syn.char_index\[2\] top.cb_syn.char_index\[1\]
+ _03080_ vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__a31o_1
XANTENNA__05494__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07192_ _03847_ _03849_ vssd1 vssd1 vccd1 vccd1 _03850_ sky130_fd_sc_hd__nand2_1
X_06143_ net499 net501 _03012_ _02767_ vssd1 vssd1 vccd1 vccd1 _03014_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_113_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06074_ net466 net159 _02942_ _02948_ vssd1 vssd1 vccd1 vccd1 _02949_ sky130_fd_sc_hd__and4_1
XANTENNA__07637__C net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09902_ net789 net629 vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__and2_1
Xfanout504 top.findLeastValue.histo_index\[0\] vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__buf_2
Xfanout515 top.cb_syn.end_cnt\[0\] vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__clkbuf_4
Xfanout537 top.cb_syn.curr_state\[4\] vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__dlymetal6s2s_1
X_09833_ net777 net617 vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__and2_1
Xfanout548 net549 vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__buf_2
XANTENNA__07493__X _04084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout526 top.translation.index\[0\] vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout388_A net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout559 net560 vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__clkbuf_4
XFILLER_100_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05454__A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09764_ net773 net613 vssd1 vssd1 vccd1 vccd1 _00378_ sky130_fd_sc_hd__and2_1
X_06976_ top.findLeastValue.val2\[18\] top.findLeastValue.val2\[17\] top.findLeastValue.val2\[16\]
+ top.findLeastValue.val2\[15\] vssd1 vssd1 vccd1 vccd1 _03634_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout176_X net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08715_ _02517_ _04904_ _04906_ vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__o21a_1
X_09695_ net804 net644 vssd1 vssd1 vccd1 vccd1 _00309_ sky130_fd_sc_hd__and2_1
X_05927_ top.WB.CPU_DAT_O\[28\] net1435 net304 vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__mux2_1
XANTENNA__09160__A1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08646_ net1692 _04854_ vssd1 vssd1 vccd1 vccd1 _01496_ sky130_fd_sc_hd__xnor2_1
X_05858_ top.compVal\[9\] net170 net156 top.WB.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1
+ _02284_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_1_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08577_ _04481_ _04535_ vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__nand2_4
X_05789_ top.hTree.state\[7\] top.hTree.state\[8\] vssd1 vssd1 vccd1 vccd1 _02809_
+ sky130_fd_sc_hd__or2_4
XANTENNA__08346__S0 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10519__B net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07528_ _04113_ _04118_ _04069_ vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__mux2_1
X_07459_ top.cb_syn.i\[3\] top.cb_syn.cb_length\[3\] vssd1 vssd1 vccd1 vccd1 _04050_
+ sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout510_X net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10470_ net728 net568 vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__and2_1
X_09129_ net469 net1209 _05135_ net1461 vssd1 vssd1 vccd1 vccd1 _00050_ sky130_fd_sc_hd__a22o_1
XANTENNA__07777__A2 _04326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08005__A top.cb_syn.h_element\[63\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold580 top.hTree.tree_reg\[39\] vssd1 vssd1 vccd1 vccd1 net1533 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11022_ clknet_leaf_20_clk _01570_ _00377_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[52\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold591 _01842_ vssd1 vssd1 vccd1 vccd1 net1544 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_106_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__11139__Q top.cb_syn.char_path_n\[41\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06894__S net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05712__B2 top.WB.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11855_ clknet_leaf_100_clk _02371_ _01210_ vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__dfrtp_1
X_10806_ clknet_leaf_51_clk _01392_ _00225_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.max_index\[6\]
+ sky130_fd_sc_hd__dfrtp_2
X_11786_ clknet_leaf_75_clk _00021_ _01141_ vssd1 vssd1 vccd1 vccd1 top.hTree.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10737_ clknet_leaf_118_clk _01336_ _00156_ vssd1 vssd1 vccd1 vccd1 top.path\[113\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10668_ clknet_leaf_118_clk _01267_ _00087_ vssd1 vssd1 vccd1 vccd1 top.path\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 SEL_O[2] sky130_fd_sc_hd__buf_2
X_10599_ net752 net592 vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__and2_1
XFILLER_99_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06830_ top.findLeastValue.val1\[0\] net130 net114 net1664 vssd1 vssd1 vccd1 vccd1
+ _02008_ sky130_fd_sc_hd__o22a_1
XANTENNA__10180__A net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06761_ net287 net152 vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__and2_1
XANTENNA__09142__A1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06692_ _02436_ top.findLeastValue.val2\[13\] vssd1 vssd1 vccd1 vccd1 _03480_ sky130_fd_sc_hd__nand2_1
X_05712_ net32 net417 net359 top.WB.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 _02346_
+ sky130_fd_sc_hd__a22o_1
X_09480_ net723 net563 vssd1 vssd1 vccd1 vccd1 _00094_ sky130_fd_sc_hd__and2_1
X_08500_ net1442 top.cb_syn.char_path_n\[76\] net221 vssd1 vssd1 vccd1 vccd1 _01594_
+ sky130_fd_sc_hd__mux2_1
X_08431_ top.cb_syn.char_path_n\[57\] net392 net331 top.cb_syn.char_path_n\[58\] net507
+ vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__a221o_1
XFILLER_63_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05561__X _02656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05643_ top.cb_syn.char_path\[6\] net558 net313 top.cb_syn.char_path\[102\] vssd1
+ vssd1 vccd1 vccd1 _02724_ sky130_fd_sc_hd__a22o_1
XANTENNA__05703__B2 top.WB.CPU_DAT_O\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06900__A0 top.compVal\[33\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05574_ net1260 net139 _02666_ net175 vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__a22o_1
X_08362_ top.cb_syn.end_cnt\[4\] _04719_ _04720_ vssd1 vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__or3_1
X_08293_ top.cb_syn.char_path_n\[23\] net383 net342 top.cb_syn.char_path_n\[21\] net187
+ vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__a221o_1
XANTENNA__11512__Q top.findLeastValue.least1\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07313_ net269 _03941_ _03942_ net274 top.findLeastValue.sum\[17\] vssd1 vssd1 vccd1
+ vccd1 _01913_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_34_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05467__B1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07244_ net272 _03890_ _03891_ net277 net1639 vssd1 vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__a32o_1
XFILLER_118_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07175_ top.findLeastValue.val1\[33\] top.findLeastValue.val2\[33\] top.findLeastValue.val2\[32\]
+ top.findLeastValue.val1\[32\] vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__a22o_1
X_06126_ top.findLeastValue.histo_index\[8\] _02481_ _02549_ _02574_ vssd1 vssd1 vccd1
+ vccd1 _02998_ sky130_fd_sc_hd__a31o_1
XANTENNA__06967__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06057_ net1037 net142 net137 vssd1 vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__a21o_1
XANTENNA__06196__A1_N net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08169__C1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout312 net313 vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__clkbuf_4
Xfanout301 net303 vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__clkbuf_2
Xfanout323 net324 vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__clkbuf_4
XFILLER_101_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout345 net349 vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__buf_2
Xfanout334 net336 vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__buf_2
Xfanout356 _02926_ vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08184__A2 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout293_X net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout367 _02567_ vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__buf_2
Xfanout389 net390 vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout378 net390 vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__buf_2
X_09816_ net744 net584 vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__and2_1
X_09747_ net765 net605 vssd1 vssd1 vccd1 vccd1 _00361_ sky130_fd_sc_hd__and2_1
X_06959_ top.findLeastValue.val2\[4\] net149 net122 _03621_ vssd1 vssd1 vccd1 vccd1
+ _01946_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout558_X net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09678_ net782 net622 vssd1 vssd1 vccd1 vccd1 _00292_ sky130_fd_sc_hd__and2_1
XANTENNA__08341__C1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08629_ _04828_ _04835_ _04842_ _04826_ top.cb_syn.num_lefts\[2\] vssd1 vssd1 vccd1
+ vccd1 _01501_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_53_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ clknet_leaf_57_clk top.dut.bit_buf_next\[12\] _00995_ vssd1 vssd1 vccd1 vccd1
+ top.dut.bit_buf\[12\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10249__B net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11571_ clknet_leaf_109_clk _02119_ _00926_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10522_ net865 net705 vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__and2_1
XFILLER_10_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10453_ net748 net588 vssd1 vssd1 vccd1 vccd1 _01067_ sky130_fd_sc_hd__and2_1
XFILLER_108_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10384_ net812 net652 vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__and2_1
XANTENNA__05646__X _02727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05630__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08175__A2 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11005_ clknet_leaf_16_clk _01553_ _00360_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09372__B2 _04298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_13_0_clk_X clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11838_ clknet_leaf_121_clk _02354_ _01193_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[16\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_14_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_40_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_clk sky130_fd_sc_hd__clkbuf_8
X_11769_ clknet_leaf_103_clk _02302_ _01124_ vssd1 vssd1 vccd1 vccd1 top.compVal\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06653__A _03424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06949__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08980_ top.WB.CPU_DAT_O\[12\] net1280 net322 vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__mux2_1
X_07931_ net488 _04449_ vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__or2_1
XFILLER_110_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08166__A2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07862_ net426 _04394_ _04395_ net261 vssd1 vssd1 vccd1 vccd1 _04396_ sky130_fd_sc_hd__o211a_1
XFILLER_113_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09601_ net856 net696 vssd1 vssd1 vccd1 vccd1 _00215_ sky130_fd_sc_hd__and2_1
X_06813_ top.findLeastValue.val1\[17\] net128 net112 net1691 vssd1 vssd1 vccd1 vccd1
+ _02025_ sky130_fd_sc_hd__o22a_1
X_07793_ net441 net1536 net253 net1724 _04340_ vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__a221o_1
X_09532_ net756 net596 vssd1 vssd1 vccd1 vccd1 _00146_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_39_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06744_ _02414_ top.findLeastValue.val2\[34\] vssd1 vssd1 vccd1 vccd1 _03532_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout253_A net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09463_ net754 net594 vssd1 vssd1 vccd1 vccd1 _00077_ sky130_fd_sc_hd__and2_1
X_06675_ _02446_ top.findLeastValue.val2\[3\] top.findLeastValue.val2\[2\] _02447_
+ vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__o22a_1
X_08414_ _02505_ _04769_ _04772_ vssd1 vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__or3_1
X_09394_ net988 net240 _05272_ _05273_ vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__a22o_1
X_05626_ _02708_ _02709_ vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__or2_1
X_08345_ net512 _04702_ _04703_ vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__a21oi_1
X_05557_ top.cb_syn.char_path\[84\] net553 net544 top.cb_syn.char_path\[52\] vssd1
+ vssd1 vccd1 vccd1 _02652_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_50_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_31_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout139_X net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout518_A net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout420_A net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09858__B net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07524__S1 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05488_ net1038 net139 net175 vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__a21o_1
X_08276_ top.cb_syn.char_path_n\[31\] net207 _04665_ vssd1 vssd1 vccd1 vccd1 _01677_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_59_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07227_ _03665_ _03669_ _03877_ _03667_ _03663_ vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__a311o_1
X_07158_ _03806_ _03814_ _03815_ _03801_ vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__o211a_1
X_06109_ top.sram_interface.init_counter\[7\] _02946_ top.sram_interface.init_counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02981_ sky130_fd_sc_hd__a21oi_1
X_07089_ top.findLeastValue.val1\[3\] top.findLeastValue.val2\[3\] vssd1 vssd1 vccd1
+ vccd1 _03747_ sky130_fd_sc_hd__nand2_1
XANTENNA__05612__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout120 net121 vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_98_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_98_clk sky130_fd_sc_hd__clkbuf_8
Xfanout131 net132 vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout675_X net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout142 net143 vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout153 _03548_ vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__buf_2
Xfanout164 net166 vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__clkbuf_4
Xfanout175 net176 vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__buf_4
XANTENNA__06168__B2 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout186 net194 vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__clkbuf_2
Xfanout197 net211 vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09106__A1 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout842_X net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05679__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11623_ clknet_leaf_68_clk _02171_ _00978_ vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08617__B1 _04826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08672__B net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_22_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07515__S1 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06891__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11554_ clknet_leaf_123_clk _02102_ _00909_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_109_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10505_ net809 net649 vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__and2_1
X_11485_ clknet_leaf_102_clk _02033_ _00840_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[25\]
+ sky130_fd_sc_hd__dfstp_1
X_10436_ net873 net713 vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__and2_1
XANTENNA__05851__B1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10367_ net798 net638 vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_94_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10298_ net723 net563 vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__and2_1
XANTENNA__08148__A2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_89_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_89_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_108_Left_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05906__A1 top.CB_read_complete vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08339__S top.cb_syn.end_cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06460_ top.histogram.total\[15\] _03268_ _03281_ vssd1 vssd1 vccd1 vccd1 _03283_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_16_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05411_ top.translation.resEn vssd1 vssd1 vccd1 vccd1 _02519_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_117_Left_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_103_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_13_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_8
X_08130_ top.cb_syn.char_path_n\[104\] net199 _04592_ vssd1 vssd1 vccd1 vccd1 _01750_
+ sky130_fd_sc_hd__o21a_1
X_06391_ net1148 _03231_ net300 vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__mux2_1
X_05342_ top.sram_interface.zero_cnt\[0\] vssd1 vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__inv_2
X_08061_ net439 _04540_ net246 vssd1 vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__a21oi_1
X_07012_ top.findLeastValue.val1\[36\] top.findLeastValue.val2\[36\] vssd1 vssd1 vccd1
+ vccd1 _03670_ sky130_fd_sc_hd__or2_1
XANTENNA__05842__B1 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08963_ top.WB.CPU_DAT_O\[29\] net1343 net321 vssd1 vssd1 vccd1 vccd1 _01348_ sky130_fd_sc_hd__mux2_1
XANTENNA__05446__B top.CB_read_complete vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07914_ top.findLeastValue.sum\[5\] top.hTree.tree_reg\[5\] net283 vssd1 vssd1 vccd1
+ vccd1 _04437_ sky130_fd_sc_hd__mux2_1
X_08894_ _02454_ top.hTree.closing net489 _05063_ vssd1 vssd1 vccd1 vccd1 _05064_
+ sky130_fd_sc_hd__a31o_1
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07845_ top.findLeastValue.sum\[19\] _04381_ net394 vssd1 vssd1 vccd1 vccd1 _04382_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07898__B2 top.findLeastValue.sum\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07362__A3 _03547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07661__B net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07776_ net490 _04325_ vssd1 vssd1 vccd1 vccd1 _04327_ sky130_fd_sc_hd__or2_1
XFILLER_17_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09515_ net725 net565 vssd1 vssd1 vccd1 vccd1 _00129_ sky130_fd_sc_hd__and2_1
X_06727_ _02422_ top.findLeastValue.val2\[28\] _02487_ net494 _03507_ vssd1 vssd1
+ vccd1 vccd1 _03515_ sky130_fd_sc_hd__o221a_1
X_09446_ net867 net707 vssd1 vssd1 vccd1 vccd1 _00060_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout256_X net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06658_ _02406_ top.findLeastValue.val2\[45\] top.findLeastValue.val2\[44\] _02407_
+ vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__o22ai_1
XANTENNA_fanout802_A net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout423_X net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09377_ net1019 net238 net215 _04278_ vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__a22o_1
X_06589_ _03353_ _03369_ _03377_ vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__a21o_1
X_05609_ top.hTree.node_reg\[44\] net310 _02695_ net473 vssd1 vssd1 vccd1 vccd1 _02696_
+ sky130_fd_sc_hd__a22o_1
X_08328_ top.cb_syn.char_path_n\[5\] net200 _04691_ vssd1 vssd1 vccd1 vccd1 _01651_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__11700__Q top.TRN_sram_complete vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10527__B net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08259_ top.cb_syn.char_path_n\[40\] net378 net337 top.cb_syn.char_path_n\[38\] net183
+ vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__a221o_1
XANTENNA__09024__A0 top.WB.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_106_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11270_ clknet_leaf_106_clk _01818_ _00625_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_106_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10221_ net811 net651 vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__and2_1
X_10152_ net814 net654 vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__and2_1
X_10083_ net864 net704 vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__and2_1
XFILLER_87_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold9 top.hTree.state\[10\] vssd1 vssd1 vccd1 vccd1 net962 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input29_A DAT_I[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10985_ clknet_leaf_6_clk _01533_ _00340_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11606_ clknet_leaf_63_clk _02154_ _00961_ vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08066__A1 _02506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06077__B1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11537_ clknet_leaf_0_clk _02085_ _00892_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07813__A1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold409 top.path\[68\] vssd1 vssd1 vccd1 vccd1 net1362 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09015__A0 top.WB.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11468_ clknet_leaf_95_clk _02016_ _00823_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[8\]
+ sky130_fd_sc_hd__dfstp_2
X_10419_ net870 net710 vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__and2_1
X_11399_ clknet_leaf_94_clk _01947_ _00754_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[5\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_97_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__10172__B net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05834__X _02845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05960_ top.translation.write_fin top.TRN_sram_complete top.translation.totalEn vssd1
+ vssd1 vccd1 vccd1 _02898_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07329__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_2_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_119_Right_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05891_ _02864_ _02865_ vssd1 vssd1 vccd1 vccd1 _02866_ sky130_fd_sc_hd__or2_1
XFILLER_93_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07630_ net456 net1055 net257 _04208_ vssd1 vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_105_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07561_ net536 _04146_ _04151_ net530 _04147_ vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__a221o_1
XFILLER_80_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06512_ net1722 _03277_ net1479 vssd1 vssd1 vccd1 vccd1 _03311_ sky130_fd_sc_hd__a21oi_1
X_09300_ top.histogram.total\[4\] net409 net326 top.histogram.total\[5\] net521 vssd1
+ vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__o221a_1
X_07492_ top.cb_syn.char_path_n\[16\] top.cb_syn.char_path_n\[15\] top.cb_syn.char_path_n\[14\]
+ top.cb_syn.char_path_n\[13\] net400 net351 vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__mux4_1
X_06443_ top.header_synthesis.count\[0\] _03245_ _03263_ vssd1 vssd1 vccd1 vccd1 _03267_
+ sky130_fd_sc_hd__a21boi_1
X_09231_ _04489_ _05199_ vssd1 vssd1 vccd1 vccd1 _05200_ sky130_fd_sc_hd__or2_2
X_09162_ net449 net1597 _03321_ _05102_ vssd1 vssd1 vccd1 vccd1 _00029_ sky130_fd_sc_hd__a22o_1
XANTENNA__08057__A1 top.cb_syn.end_cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06374_ top.hist_data_o\[15\] _03183_ vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__xor2_1
XFILLER_119_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08113_ top.cb_syn.char_path_n\[113\] net375 net335 top.cb_syn.char_path_n\[111\]
+ net180 vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__a221o_1
X_05325_ top.compVal\[16\] vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__inv_2
XFILLER_119_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09093_ net452 net479 _05112_ vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout216_A net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09006__A0 top.WB.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08044_ _02873_ _04537_ vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_116_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_1_0_clk_X clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09995_ net846 net686 vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout585_A net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08946_ top.WB.CPU_DAT_O\[27\] top.cb_syn.h_element\[59\] net369 vssd1 vssd1 vccd1
+ vccd1 _01364_ sky130_fd_sc_hd__mux2_1
XFILLER_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05594__A2 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08877_ _05043_ _05047_ _05052_ vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__or3_1
XFILLER_29_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09174__A_N top.cb_syn.char_path_n\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07828_ net445 net1551 net253 top.findLeastValue.sum\[23\] _04368_ vssd1 vssd1 vccd1
+ vccd1 _01828_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_67_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07759_ top.findLeastValue.sum\[36\] top.hTree.tree_reg\[36\] net280 vssd1 vssd1
+ vccd1 vccd1 _04313_ sky130_fd_sc_hd__mux2_1
XANTENNA__09599__A net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10770_ clknet_leaf_78_clk _01369_ _00189_ vssd1 vssd1 vccd1 vccd1 top.hTree.nulls\[46\]
+ sky130_fd_sc_hd__dfrtp_1
X_09429_ net998 vssd1 vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__clkbuf_1
XFILLER_100_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06059__B1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11322_ clknet_leaf_75_clk _01870_ _00677_ vssd1 vssd1 vccd1 vccd1 top.WorR sky130_fd_sc_hd__dfrtp_2
XFILLER_109_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11253_ clknet_leaf_75_clk _01801_ _00608_ vssd1 vssd1 vccd1 vccd1 top.hTree.nullSumIndex\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10204_ net830 net670 vssd1 vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__and2_1
X_11184_ clknet_leaf_19_clk _01732_ _00539_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[86\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05585__A2 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10135_ net832 net672 vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__and2_1
X_10066_ net851 net691 vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__and2_1
XFILLER_94_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_90_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10968_ clknet_leaf_40_clk _01516_ _00323_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_index\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_26_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10899_ clknet_leaf_39_clk top.header_synthesis.next_header\[4\] _00254_ vssd1 vssd1
+ vccd1 vccd1 top.header_synthesis.header\[4\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06090_ top.cb_syn.char_index\[5\] _02962_ vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__and2_1
Xhold206 top.cb_syn.char_path\[16\] vssd1 vssd1 vccd1 vccd1 net1159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold217 top.histogram.sram_out\[8\] vssd1 vssd1 vccd1 vccd1 net1170 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xhold239 top.cb_syn.char_path\[84\] vssd1 vssd1 vccd1 vccd1 net1192 sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 top.hTree.nulls\[53\] vssd1 vssd1 vccd1 vccd1 net1181 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_98_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09972__A net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout719 net44 vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__clkbuf_4
Xfanout708 net717 vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__buf_1
X_08800_ top.path\[18\] top.path\[19\] net524 vssd1 vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__mux2_1
XFILLER_98_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06773__A1 top.findLeastValue.least1\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05576__A2 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09780_ net765 net605 vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08762__A2 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06992_ top.findLeastValue.val1\[34\] top.findLeastValue.val1\[33\] top.findLeastValue.val1\[32\]
+ top.findLeastValue.val1\[31\] vssd1 vssd1 vccd1 vccd1 _03650_ sky130_fd_sc_hd__and4_1
X_08731_ _04914_ _04912_ top.header_synthesis.count\[2\] vssd1 vssd1 vccd1 vccd1 _04915_
+ sky130_fd_sc_hd__mux2_1
X_05943_ top.WB.CPU_DAT_O\[12\] net1342 net306 vssd1 vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__mux2_1
X_08662_ top.cb_syn.wait_cycle _04865_ _04863_ vssd1 vssd1 vccd1 vccd1 _01491_ sky130_fd_sc_hd__mux2_1
X_05874_ net449 _02453_ _02852_ net495 vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__o31a_1
X_07613_ net962 net265 _04194_ vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__a21oi_1
XFILLER_66_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08593_ _04815_ top.cb_syn.char_index\[0\] _04807_ vssd1 vssd1 vccd1 vccd1 _01510_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__11515__Q top.findLeastValue.least1\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout166_A _03423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07544_ _04134_ _02526_ _02498_ vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__and3b_2
X_07475_ _04045_ _04046_ _04061_ vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__and3_1
XANTENNA__09212__A top.controller.fin_reg\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06426_ top.header_synthesis.count\[5\] _03248_ _03252_ vssd1 vssd1 vccd1 vccd1 _03255_
+ sky130_fd_sc_hd__and3b_1
X_09214_ _05187_ _05188_ vssd1 vssd1 vccd1 vccd1 _00015_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_62_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout333_A net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09145_ net469 net1102 net1209 _05135_ vssd1 vssd1 vccd1 vccd1 _00040_ sky130_fd_sc_hd__a22o_1
X_06357_ top.hist_data_o\[21\] _03188_ vssd1 vssd1 vccd1 vccd1 _03210_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout219_X net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout121_X net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06288_ top.cw1\[1\] top.cw1\[0\] vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__or2_1
X_09076_ _03323_ net257 vssd1 vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__or2_1
XANTENNA__07253__A2 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05308_ top.compVal\[32\] vssd1 vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__inv_2
X_08027_ top.cb_syn.count\[1\] top.cb_syn.count\[0\] top.cb_syn.count\[2\] vssd1 vssd1
+ vccd1 vccd1 _04525_ sky130_fd_sc_hd__a21o_1
XFILLER_100_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold751 top.hist_data_o\[19\] vssd1 vssd1 vccd1 vccd1 net1704 sky130_fd_sc_hd__dlygate4sd3_1
Xhold773 top.findLeastValue.sum\[32\] vssd1 vssd1 vccd1 vccd1 net1726 sky130_fd_sc_hd__dlygate4sd3_1
Xhold762 top.hist_data_o\[14\] vssd1 vssd1 vccd1 vccd1 net1715 sky130_fd_sc_hd__dlygate4sd3_1
Xhold740 top.compVal\[1\] vssd1 vssd1 vccd1 vccd1 net1693 sky130_fd_sc_hd__dlygate4sd3_1
X_09978_ net780 net620 vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__and2_1
XANTENNA__05567__A2 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08929_ top.WB.CPU_DAT_O\[25\] net1292 net372 vssd1 vssd1 vccd1 vccd1 _01380_ sky130_fd_sc_hd__mux2_1
XANTENNA__07713__B1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11871_ clknet_leaf_7_clk _02387_ _01226_ vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__dfrtp_1
XFILLER_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11425__Q top.findLeastValue.val2\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10822_ clknet_leaf_106_clk _01408_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_43_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08364__S1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10753_ clknet_leaf_48_clk _01352_ _00172_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06819__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10684_ clknet_leaf_120_clk _01283_ _00103_ vssd1 vssd1 vccd1 vccd1 top.path\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09313__S0 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11305_ clknet_leaf_71_clk _01853_ _00660_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[48\]
+ sky130_fd_sc_hd__dfrtp_1
X_11236_ clknet_leaf_30_clk _01784_ _00591_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_106_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05558__A2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11167_ clknet_leaf_13_clk _01715_ _00522_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[69\]
+ sky130_fd_sc_hd__dfrtp_2
X_10118_ net823 net663 vssd1 vssd1 vccd1 vccd1 _00732_ sky130_fd_sc_hd__and2_1
X_11098_ clknet_leaf_35_clk net1063 _00453_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.end_cond
+ sky130_fd_sc_hd__dfrtp_1
X_10049_ net859 net699 vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__and2_1
X_05590_ net457 top.hTree.node_reg\[47\] net361 net420 top.hTree.node_reg\[15\] vssd1
+ vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__a32o_1
XANTENNA__08347__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09209__B1 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07260_ _03691_ _03902_ _03689_ vssd1 vssd1 vccd1 vccd1 _03904_ sky130_fd_sc_hd__a21bo_1
XFILLER_117_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06211_ _02507_ _02956_ _02578_ vssd1 vssd1 vccd1 vccd1 _03080_ sky130_fd_sc_hd__a21bo_1
X_07191_ top.findLeastValue.val1\[43\] top.findLeastValue.val2\[43\] vssd1 vssd1 vccd1
+ vccd1 _03849_ sky130_fd_sc_hd__or2_1
X_06142_ net501 _03012_ _02767_ vssd1 vssd1 vccd1 vccd1 _03013_ sky130_fd_sc_hd__a21o_1
XANTENNA__08432__A1 _02505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_83_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06073_ top.sram_interface.init_counter\[9\] _02947_ top.sram_interface.init_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02948_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_113_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09901_ net789 net629 vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__and2_1
XFILLER_113_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout505 top.cb_syn.end_cnt\[3\] vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_98_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout538 top.cb_syn.curr_state\[2\] vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__clkbuf_4
Xfanout516 top.cb_syn.end_cnt\[0\] vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09832_ net770 net610 vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__and2_1
XANTENNA__05549__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout527 net528 vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__buf_4
Xfanout549 top.sram_interface.word_cnt\[8\] vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__clkbuf_4
X_09763_ net773 net613 vssd1 vssd1 vccd1 vccd1 _00377_ sky130_fd_sc_hd__and2_1
XANTENNA__07943__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08714_ _04903_ _04905_ top.cb_syn.i\[6\] vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_21_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06975_ top.findLeastValue.val2\[22\] top.findLeastValue.val2\[21\] top.findLeastValue.val2\[20\]
+ top.findLeastValue.val2\[19\] vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout283_A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05454__B net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09694_ net802 net642 vssd1 vssd1 vccd1 vccd1 _00308_ sky130_fd_sc_hd__and2_1
XFILLER_82_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05926_ top.WB.CPU_DAT_O\[29\] net1338 net305 vssd1 vssd1 vccd1 vccd1 _02263_ sky130_fd_sc_hd__mux2_1
X_08645_ _04846_ _04848_ net210 vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__o21ai_1
X_05857_ top.compVal\[10\] net170 net156 top.WB.CPU_DAT_O\[10\] vssd1 vssd1 vccd1
+ vccd1 _02285_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_1_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08576_ _02498_ _04562_ _04806_ net1449 vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout548_A net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout169_X net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_36_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05788_ top.hTree.state\[7\] top.hTree.state\[8\] vssd1 vssd1 vccd1 vccd1 _02808_
+ sky130_fd_sc_hd__nor2_1
X_07527_ _04114_ _04115_ _04116_ _04117_ _04072_ _04071_ vssd1 vssd1 vccd1 vccd1 _04118_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08346__S1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07458_ top.cb_syn.i\[3\] top.cb_syn.cb_length\[3\] vssd1 vssd1 vccd1 vccd1 _04049_
+ sky130_fd_sc_hd__and2b_1
X_07389_ top.dut.bit_buf\[8\] top.dut.bit_buf\[1\] net722 vssd1 vssd1 vccd1 vccd1
+ _03991_ sky130_fd_sc_hd__mux2_1
XFILLER_10_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_20_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06409_ top.hist_data_o\[2\] _03173_ vssd1 vssd1 vccd1 vccd1 _03243_ sky130_fd_sc_hd__xnor2_1
X_09128_ net562 _05131_ _05141_ _02893_ vssd1 vssd1 vccd1 vccd1 _00038_ sky130_fd_sc_hd__a211o_1
XFILLER_108_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09059_ _03270_ _03316_ _05089_ net466 vssd1 vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__o31ai_4
XTAP_TAPCELL_ROW_75_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold570 top.cb_syn.char_index\[7\] vssd1 vssd1 vccd1 vccd1 net1523 sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 top.histogram.total\[22\] vssd1 vssd1 vccd1 vccd1 net1534 sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 top.histogram.wr_r_en\[1\] vssd1 vssd1 vccd1 vccd1 net1545 sky130_fd_sc_hd__dlygate4sd3_1
X_11021_ clknet_leaf_21_clk _01569_ _00376_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_9_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_109_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07934__A0 top.findLeastValue.sum\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05960__A2 top.TRN_sram_complete vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input11_A DAT_I[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11854_ clknet_leaf_86_clk _02370_ _01209_ vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_56_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10805_ clknet_leaf_51_clk _01391_ _00224_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.max_index\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__05712__A2 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11785_ clknet_leaf_74_clk _00020_ _01140_ vssd1 vssd1 vccd1 vccd1 top.hTree.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10736_ clknet_leaf_118_clk _01335_ _00155_ vssd1 vssd1 vccd1 vccd1 top.path\[112\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10667_ clknet_leaf_118_clk _01266_ _00086_ vssd1 vssd1 vccd1 vccd1 top.path\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10598_ net840 net680 vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__and2_1
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 SEL_O[3] sky130_fd_sc_hd__buf_2
X_11219_ clknet_leaf_25_clk _01767_ _00574_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[121\]
+ sky130_fd_sc_hd__dfrtp_2
Xoutput90 net90 vssd1 vssd1 vccd1 vccd1 DAT_O[25] sky130_fd_sc_hd__buf_2
XANTENNA__07925__A0 top.findLeastValue.sum\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06003__X _02926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10180__B net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06760_ _03424_ _03441_ _03547_ net287 vssd1 vssd1 vccd1 vccd1 _03548_ sky130_fd_sc_hd__o211ai_1
XFILLER_102_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06691_ _02437_ top.findLeastValue.val2\[12\] vssd1 vssd1 vccd1 vccd1 _03479_ sky130_fd_sc_hd__nor2_1
X_05711_ net33 net416 net309 top.WB.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1 _02347_
+ sky130_fd_sc_hd__o22a_1
X_08430_ net507 _04782_ _04784_ _04785_ _02504_ vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__o221a_1
X_05642_ top.cb_syn.char_path\[70\] net552 net543 top.cb_syn.char_path\[38\] vssd1
+ vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__a22o_1
XANTENNA__05703__A2 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05573_ top.histogram.sram_out\[18\] net364 _02664_ _02665_ vssd1 vssd1 vccd1 vccd1
+ _02666_ sky130_fd_sc_hd__a211o_1
X_08361_ net508 _04709_ _04711_ _04712_ _02504_ vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__o221a_1
X_08292_ top.cb_syn.char_path_n\[23\] net204 _04673_ vssd1 vssd1 vccd1 vccd1 _01669_
+ sky130_fd_sc_hd__o21a_1
X_07312_ _03785_ _03940_ vssd1 vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__nand2_1
X_07243_ _03821_ _03889_ _03827_ vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__a21bo_1
XANTENNA_fanout129_A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07174_ _03817_ _03820_ _03831_ vssd1 vssd1 vccd1 vccd1 _03832_ sky130_fd_sc_hd__a21o_1
X_06125_ top.cw1\[7\] _02996_ _02573_ vssd1 vssd1 vccd1 vccd1 _02997_ sky130_fd_sc_hd__a21o_1
XFILLER_105_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06056_ net471 net368 net159 net412 vssd1 vssd1 vccd1 vccd1 _02941_ sky130_fd_sc_hd__and4_1
Xfanout302 net303 vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout313 net315 vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__buf_2
Xfanout357 _02926_ vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__clkbuf_4
Xfanout346 net348 vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__clkbuf_4
Xfanout335 net336 vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input3_A DAT_I[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout324 _05087_ vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__buf_2
X_09815_ net740 net580 vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__and2_1
Xfanout368 _02550_ vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout286_X net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout379 net390 vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout665_A net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09746_ net787 net627 vssd1 vssd1 vccd1 vccd1 _00360_ sky130_fd_sc_hd__and2_1
X_06958_ top.compVal\[4\] top.findLeastValue.val1\[4\] net166 vssd1 vssd1 vccd1 vccd1
+ _03621_ sky130_fd_sc_hd__mux2_1
X_09677_ net800 net640 vssd1 vssd1 vccd1 vccd1 _00291_ sky130_fd_sc_hd__and2_1
X_05909_ top.sram_interface.CB_write_counter\[1\] _02452_ vssd1 vssd1 vccd1 vccd1
+ _02882_ sky130_fd_sc_hd__nor2_1
XFILLER_27_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08628_ top.cb_syn.num_lefts\[1\] top.cb_syn.num_lefts\[0\] top.cb_syn.num_lefts\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout453_X net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06889_ top.findLeastValue.val2\[39\] net150 net123 _03586_ vssd1 vssd1 vccd1 vccd1
+ _01981_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_53_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_fanout718_X net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08559_ net1146 top.cb_syn.char_path_n\[17\] net222 vssd1 vssd1 vccd1 vccd1 _01535_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11570_ clknet_leaf_106_clk _02118_ _00925_ vssd1 vssd1 vccd1 vccd1 top.histogram.sram_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10521_ net861 net701 vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__and2_1
XANTENNA__07852__C1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10452_ net747 net587 vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__and2_1
X_10383_ net813 net653 vssd1 vssd1 vccd1 vccd1 _00997_ sky130_fd_sc_hd__and2_1
XANTENNA__08450__S net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11004_ clknet_leaf_17_clk _01552_ _00359_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_88_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06758__X _03546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05662__X _02740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11837_ clknet_leaf_115_clk _02353_ _01192_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__05697__B2 top.WB.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11768_ clknet_leaf_102_clk _02301_ _01123_ vssd1 vssd1 vccd1 vccd1 top.compVal\[26\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__05449__A1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10719_ clknet_leaf_3_clk _01318_ _00138_ vssd1 vssd1 vccd1 vccd1 top.path\[95\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11699_ clknet_leaf_66_clk _02232_ _01054_ vssd1 vssd1 vccd1 vccd1 top.FLV_done sky130_fd_sc_hd__dfrtp_1
XANTENNA__08399__A0 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07930_ top.findLeastValue.sum\[2\] _04449_ net398 vssd1 vssd1 vccd1 vccd1 _04450_
+ sky130_fd_sc_hd__mux2_1
X_07861_ net483 _04393_ vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__or2_1
XFILLER_110_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09600_ net851 net691 vssd1 vssd1 vccd1 vccd1 _00214_ sky130_fd_sc_hd__and2_1
X_07792_ net428 _04338_ _04339_ net259 vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__o211a_1
X_06812_ top.findLeastValue.val1\[18\] net128 net112 top.compVal\[18\] vssd1 vssd1
+ vccd1 vccd1 _02026_ sky130_fd_sc_hd__o22a_1
X_09531_ net756 net596 vssd1 vssd1 vccd1 vccd1 _00145_ sky130_fd_sc_hd__and2_1
X_06743_ top.compVal\[37\] _02485_ vssd1 vssd1 vccd1 vccd1 _03531_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_108_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09462_ net751 net591 vssd1 vssd1 vccd1 vccd1 _00076_ sky130_fd_sc_hd__and2_1
X_06674_ _02448_ top.findLeastValue.val2\[0\] _03459_ _03460_ _03461_ vssd1 vssd1
+ vccd1 vccd1 _03462_ sky130_fd_sc_hd__a311o_1
XANTENNA__08874__A1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08413_ net511 _04770_ _04771_ vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__a21oi_1
X_09393_ top.hTree.nulls\[51\] net405 net244 vssd1 vssd1 vccd1 vccd1 _05273_ sky130_fd_sc_hd__o21a_1
X_05625_ top.cb_syn.char_path\[9\] net558 net313 top.cb_syn.char_path\[105\] vssd1
+ vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__a22o_1
X_08344_ top.cb_syn.char_path_n\[89\] net393 net331 top.cb_syn.char_path_n\[90\] net507
+ vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__a221o_1
X_05556_ net1074 net144 _02651_ _02589_ vssd1 vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__a22o_1
XFILLER_51_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05487_ net160 _02592_ vssd1 vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__and2b_1
X_08275_ top.cb_syn.char_path_n\[32\] net386 net345 top.cb_syn.char_path_n\[30\] net190
+ vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout413_A net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07226_ _03665_ _03669_ _03877_ _03667_ vssd1 vssd1 vccd1 vccd1 _03878_ sky130_fd_sc_hd__a31o_1
XFILLER_22_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05860__B2 top.WB.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09051__A1 top.WB.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07157_ _03803_ _03800_ vssd1 vssd1 vccd1 vccd1 _03815_ sky130_fd_sc_hd__nand2b_1
X_06108_ net1383 net143 _02980_ net159 vssd1 vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__a22o_1
XANTENNA__05747__X _02782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07675__A net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout782_A net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07088_ top.findLeastValue.val1\[3\] top.findLeastValue.val2\[3\] vssd1 vssd1 vccd1
+ vccd1 _03746_ sky130_fd_sc_hd__and2_1
X_06039_ _02927_ _02929_ vssd1 vssd1 vccd1 vccd1 _02930_ sky130_fd_sc_hd__or2_1
XFILLER_59_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout121 net124 vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__clkbuf_4
Xfanout143 net144 vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__clkbuf_2
Xfanout154 net155 vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__clkbuf_4
Xfanout132 net133 vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__clkbuf_2
Xfanout165 net166 vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__clkbuf_4
Xfanout176 _02589_ vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__clkbuf_4
XFILLER_87_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout187 net194 vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__buf_2
Xfanout198 net211 vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__clkbuf_2
XANTENNA__05923__A _02892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09729_ net769 net609 vssd1 vssd1 vccd1 vccd1 _00343_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout835_X net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07668__A2 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11622_ clknet_leaf_39_clk _02170_ _00977_ vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08617__A1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11553_ clknet_leaf_123_clk _02101_ _00908_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10504_ net753 net593 vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__and2_1
X_11484_ clknet_leaf_103_clk _02032_ _00839_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[24\]
+ sky130_fd_sc_hd__dfstp_2
X_10435_ net875 net715 vssd1 vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__and2_1
XANTENNA__05851__B2 top.WB.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09042__A1 top.WB.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10366_ net852 net692 vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_94_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05603__A1 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10297_ net724 net564 vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__and2_1
XFILLER_2_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06800__B1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05410_ top.cb_syn.i\[5\] vssd1 vssd1 vccd1 vccd1 _02518_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_06390_ top.hist_data_o\[9\] _03179_ vssd1 vssd1 vccd1 vccd1 _03231_ sky130_fd_sc_hd__xor2_1
X_05341_ top.sram_interface.zero_cnt\[1\] vssd1 vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__inv_2
XANTENNA__06095__A1 top.cb_syn.char_index\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08060_ _04550_ net246 net505 _04549_ vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07292__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07011_ top.findLeastValue.val1\[36\] top.findLeastValue.val2\[36\] vssd1 vssd1 vccd1
+ vccd1 _03669_ sky130_fd_sc_hd__nand2_1
XANTENNA__09033__A1 top.WB.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05842__B2 top.WB.CPU_DAT_O\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__05567__X _02661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08962_ top.WB.CPU_DAT_O\[30\] net1101 net321 vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__mux2_1
X_08893_ net492 _02809_ vssd1 vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__nor2_1
X_07913_ net442 net1578 net252 top.findLeastValue.sum\[6\] _04436_ vssd1 vssd1 vccd1
+ vccd1 _01811_ sky130_fd_sc_hd__a221o_1
XFILLER_69_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07844_ top.findLeastValue.sum\[19\] top.hTree.tree_reg\[19\] net278 vssd1 vssd1
+ vccd1 vccd1 _04381_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout196_A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09215__A top.controller.fin_reg\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07661__C net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07775_ top.findLeastValue.sum\[33\] _04325_ net396 vssd1 vssd1 vccd1 vccd1 _04326_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout363_A net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09514_ net725 net565 vssd1 vssd1 vccd1 vccd1 _00128_ sky130_fd_sc_hd__and2_1
X_06726_ _02419_ top.findLeastValue.val2\[31\] vssd1 vssd1 vccd1 vccd1 _03514_ sky130_fd_sc_hd__nor2_1
X_09445_ net847 net687 vssd1 vssd1 vccd1 vccd1 _00059_ sky130_fd_sc_hd__and2_1
X_06657_ _02406_ top.findLeastValue.val2\[45\] top.findLeastValue.val2\[46\] vssd1
+ vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout628_A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout249_X net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05608_ _02693_ _02694_ vssd1 vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout151_X net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05530__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06588_ _03373_ _03375_ _03376_ _03374_ vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__or4b_1
X_09376_ net1039 net236 net214 _04282_ vssd1 vssd1 vccd1 vccd1 _01438_ sky130_fd_sc_hd__a22o_1
X_05539_ top.cb_syn.char_path\[87\] net553 net544 top.cb_syn.char_path\[55\] vssd1
+ vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__a22o_1
X_08327_ top.cb_syn.char_path_n\[6\] net379 net338 top.cb_syn.char_path_n\[4\] net183
+ vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout416_X net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07807__C1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08258_ top.cb_syn.char_path_n\[40\] net200 _04656_ vssd1 vssd1 vccd1 vccd1 _01686_
+ sky130_fd_sc_hd__o21a_1
X_07209_ _03860_ net271 vssd1 vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__nand2_1
X_10220_ net808 net648 vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__and2_1
X_08189_ top.cb_syn.char_path_n\[75\] net378 net337 top.cb_syn.char_path_n\[73\] net182
+ vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__a221o_1
XANTENNA__05597__B1 _02684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10151_ net810 net650 vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__and2_1
X_10082_ net864 net704 vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__and2_1
XFILLER_114_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__06010__A1 top.WB.CPU_DAT_O\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10984_ clknet_leaf_6_clk _01532_ _00339_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08838__A1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06849__A0 top.findLeastValue.least1\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05521__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11605_ clknet_leaf_63_clk _02153_ _00960_ vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08903__S _05072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11536_ clknet_leaf_1_clk _02084_ _00891_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11467_ clknet_leaf_95_clk _02015_ _00822_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[7\]
+ sky130_fd_sc_hd__dfstp_1
X_10418_ net870 net710 vssd1 vssd1 vccd1 vccd1 _01032_ sky130_fd_sc_hd__and2_1
X_11398_ clknet_leaf_94_clk _01946_ _00753_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[4\]
+ sky130_fd_sc_hd__dfstp_1
X_10349_ net869 net709 vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__and2_1
XANTENNA__05588__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09318__A2 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07329__A1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05890_ top.cb_syn.h_element\[61\] top.cb_syn.h_element\[60\] top.cb_syn.h_element\[59\]
+ top.cb_syn.h_element\[62\] vssd1 vssd1 vccd1 vccd1 _02865_ sky130_fd_sc_hd__or4b_1
XFILLER_66_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07560_ top.cb_syn.max_index\[7\] _04150_ vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_49_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06511_ net1636 _03279_ vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__xor2_1
X_09230_ _04488_ _05198_ _04484_ vssd1 vssd1 vccd1 vccd1 _05199_ sky130_fd_sc_hd__o21a_1
X_07491_ top.cb_syn.char_path_n\[12\] top.cb_syn.char_path_n\[11\] top.cb_syn.char_path_n\[10\]
+ top.cb_syn.char_path_n\[9\] net399 net350 vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__mux4_1
X_06442_ _03256_ _03263_ _03266_ vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__and3b_1
XANTENNA__05512__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09161_ net450 net1472 _05102_ _05107_ _05163_ vssd1 vssd1 vccd1 vccd1 _00028_ sky130_fd_sc_hd__a311o_1
X_06373_ net1094 net299 _03220_ vssd1 vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__a21o_1
XANTENNA__11801__Q top.compVal\[33\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09092_ _02937_ _05111_ vssd1 vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__nor2_2
X_08112_ top.cb_syn.char_path_n\[113\] net197 _04583_ vssd1 vssd1 vccd1 vccd1 _01759_
+ sky130_fd_sc_hd__o21a_1
X_05324_ top.compVal\[17\] vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__inv_2
XFILLER_107_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08043_ net535 top.cb_syn.curr_state\[5\] _04535_ vssd1 vssd1 vccd1 vccd1 _04537_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout209_A net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06333__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09994_ net847 net687 vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__and2_1
XFILLER_1_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout480_A net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08945_ top.WB.CPU_DAT_O\[28\] top.cb_syn.h_element\[60\] net369 vssd1 vssd1 vccd1
+ vccd1 _01365_ sky130_fd_sc_hd__mux2_1
XANTENNA__06791__A2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08876_ net527 _05040_ top.translation.index\[1\] vssd1 vssd1 vccd1 vccd1 _05052_
+ sky130_fd_sc_hd__o21a_1
X_07827_ net428 _04366_ _04367_ net267 vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout366_X net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout745_A net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07758_ net444 net1543 net254 top.findLeastValue.sum\[37\] _04312_ vssd1 vssd1 vccd1
+ vccd1 _01842_ sky130_fd_sc_hd__a221o_1
X_06709_ _02430_ top.findLeastValue.val2\[19\] top.findLeastValue.val2\[18\] _02431_
+ vssd1 vssd1 vccd1 vccd1 _03497_ sky130_fd_sc_hd__o22a_1
XFILLER_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09599__B net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07689_ net490 _04256_ vssd1 vssd1 vccd1 vccd1 _04257_ sky130_fd_sc_hd__nand2_1
X_09428_ net1016 vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__clkbuf_1
X_09359_ net1010 net242 net218 _04350_ vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__a22o_1
X_11321_ clknet_leaf_71_clk net963 _00676_ vssd1 vssd1 vccd1 vccd1 top.HT_fin_reg
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_78_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11252_ clknet_leaf_74_clk _01800_ _00607_ vssd1 vssd1 vccd1 vccd1 top.hTree.nullSumIndex\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11183_ clknet_leaf_17_clk _01731_ _00538_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[85\]
+ sky130_fd_sc_hd__dfrtp_2
X_10203_ net831 net671 vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__and2_1
XANTENNA_input41_A gpio_in[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10134_ net836 net676 vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__and2_1
XFILLER_94_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06782__A2 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10065_ net851 net691 vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__and2_1
XFILLER_63_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10967_ clknet_leaf_40_clk _01515_ _00322_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_index\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__06298__B2 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10898_ clknet_leaf_39_clk top.header_synthesis.next_header\[3\] _00253_ vssd1 vssd1
+ vccd1 vccd1 top.header_synthesis.header\[3\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_26_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07798__A1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08995__A0 top.WB.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11519_ clknet_leaf_65_clk _02067_ _00874_ vssd1 vssd1 vccd1 vccd1 top.cw1\[2\] sky130_fd_sc_hd__dfrtp_1
Xhold207 top.cb_syn.char_path\[79\] vssd1 vssd1 vccd1 vccd1 net1160 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold218 top.cb_syn.char_path\[94\] vssd1 vssd1 vccd1 vccd1 net1171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 top.path\[95\] vssd1 vssd1 vccd1 vccd1 net1182 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09972__B net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout709 net710 vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08869__A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06991_ top.findLeastValue.val1\[38\] top.findLeastValue.val1\[37\] top.findLeastValue.val1\[36\]
+ top.findLeastValue.val1\[35\] vssd1 vssd1 vccd1 vccd1 _03649_ sky130_fd_sc_hd__and4_1
X_08730_ top.cb_syn.num_lefts\[0\] top.cb_syn.num_lefts\[6\] top.cb_syn.num_lefts\[7\]
+ top.cb_syn.num_lefts\[5\] top.header_synthesis.count\[1\] top.header_synthesis.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04914_ sky130_fd_sc_hd__mux4_1
XFILLER_100_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05942_ top.WB.CPU_DAT_O\[13\] net1365 net306 vssd1 vssd1 vccd1 vccd1 _02247_ sky130_fd_sc_hd__mux2_1
X_05873_ _02760_ _02851_ vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__and2_1
X_08661_ _02554_ _02866_ _02870_ _04864_ vssd1 vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__a31o_1
X_07612_ top.hTree.state\[1\] net265 net955 vssd1 vssd1 vccd1 vccd1 _04194_ sky130_fd_sc_hd__a21oi_1
XANTENNA__05733__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08592_ top.cb_syn.h_element\[55\] top.cb_syn.h_element\[46\] net533 vssd1 vssd1
+ vccd1 vccd1 _04815_ sky130_fd_sc_hd__mux2_1
X_07543_ net530 net536 vssd1 vssd1 vccd1 vccd1 _04134_ sky130_fd_sc_hd__or2_2
XANTENNA_fanout159_A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07474_ _04044_ _04063_ vssd1 vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09212__B top.controller.fin_reg\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06289__A1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06425_ _03245_ _03248_ _03246_ vssd1 vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__a21oi_1
X_09213_ top.controller.fin_reg\[5\] top.controller.fin_reg\[6\] top.controller.fin_reg\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05188_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_62_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09144_ net546 _05139_ _05153_ vssd1 vssd1 vccd1 vccd1 _00039_ sky130_fd_sc_hd__a21o_1
XANTENNA__05500__A3 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout326_A net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06852__A net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08543__S net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06356_ net1499 _03209_ net302 vssd1 vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__mux2_1
XANTENNA__08986__A0 top.WB.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09075_ net538 net431 _04869_ _05097_ vssd1 vssd1 vccd1 vccd1 _00005_ sky130_fd_sc_hd__a211o_1
X_06287_ _02572_ _02999_ _03151_ net368 net504 vssd1 vssd1 vccd1 vccd1 _03152_ sky130_fd_sc_hd__a32o_1
X_05307_ top.compVal\[33\] vssd1 vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__inv_2
X_08026_ _04514_ _04520_ _04524_ _04509_ top.cb_syn.count\[3\] vssd1 vssd1 vccd1 vccd1
+ _01786_ sky130_fd_sc_hd__a32o_1
Xhold730 top.sram_interface.zero_cnt\[2\] vssd1 vssd1 vccd1 vccd1 net1683 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout695_A net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold741 top.cw1\[7\] vssd1 vssd1 vccd1 vccd1 net1694 sky130_fd_sc_hd__dlygate4sd3_1
Xhold752 top.sram_interface.counter_HTREE\[2\] vssd1 vssd1 vccd1 vccd1 net1705 sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 top.findLeastValue.sum\[20\] vssd1 vssd1 vccd1 vccd1 net1716 sky130_fd_sc_hd__dlygate4sd3_1
Xhold774 top.findLeastValue.sum\[34\] vssd1 vssd1 vccd1 vccd1 net1727 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09977_ net780 net620 vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__and2_1
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08928_ top.WB.CPU_DAT_O\[26\] net1327 net371 vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__mux2_1
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09163__B1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07713__A1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08859_ _05040_ vssd1 vssd1 vccd1 vccd1 _05041_ sky130_fd_sc_hd__inv_2
X_11870_ clknet_leaf_7_clk _02386_ _01225_ vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09403__A net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10821_ clknet_leaf_106_clk _01407_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_10752_ clknet_leaf_47_clk _01351_ _00171_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.h_element\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10683_ clknet_leaf_119_clk _01282_ _00102_ vssd1 vssd1 vccd1 vccd1 top.path\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08453__S net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08426__C1 _02505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06762__A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09313__S1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08977__A0 top.WB.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11304_ clknet_leaf_70_clk _01852_ _00659_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[47\]
+ sky130_fd_sc_hd__dfrtp_1
X_11235_ clknet_leaf_29_clk _01783_ _00590_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_106_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input44_X net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11166_ clknet_leaf_16_clk _01714_ _00521_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[68\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11097_ clknet_leaf_28_clk _01645_ _00452_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[127\]
+ sky130_fd_sc_hd__dfrtp_1
X_10117_ net821 net661 vssd1 vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__and2_1
X_10048_ net837 net677 vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__and2_1
Xhold90 net60 vssd1 vssd1 vccd1 vccd1 net1043 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08901__B1 _04188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05715__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_11_Left_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09209__A1 top.cb_syn.char_path_n\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06210_ top.cb_syn.max_index\[5\] _03025_ _03027_ top.hTree.nullSumIndex\[4\] vssd1
+ vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__a22o_1
XANTENNA__11351__Q top.findLeastValue.sum\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08968__A0 top.WB.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07190_ top.findLeastValue.val1\[43\] top.findLeastValue.val2\[43\] vssd1 vssd1 vccd1
+ vccd1 _03848_ sky130_fd_sc_hd__nor2_1
X_06141_ net502 net503 net504 top.findLeastValue.histo_index\[3\] vssd1 vssd1 vccd1
+ vccd1 _03012_ sky130_fd_sc_hd__a31o_1
XFILLER_8_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06072_ top.sram_interface.init_counter\[8\] top.sram_interface.init_counter\[7\]
+ _02946_ vssd1 vssd1 vccd1 vccd1 _02947_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_20_Left_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09900_ net790 net630 vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__and2_1
XFILLER_6_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_113_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout506 top.cb_syn.end_cnt\[3\] vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__clkbuf_2
Xfanout539 net540 vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__buf_2
Xfanout517 top.cb_syn.char_path_n\[1\] vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__buf_2
XANTENNA_clkload13_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09831_ net771 net611 vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__and2_1
Xfanout528 top.translation.index\[0\] vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__clkbuf_4
X_09762_ net773 net613 vssd1 vssd1 vccd1 vccd1 _00376_ sky130_fd_sc_hd__and2_1
XANTENNA__05954__A0 top.WB.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07943__B2 top.findLeastValue.sum\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07943__A1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06974_ top.findLeastValue.val2\[30\] top.findLeastValue.val2\[29\] top.findLeastValue.val2\[28\]
+ top.findLeastValue.val2\[27\] vssd1 vssd1 vccd1 vccd1 _03632_ sky130_fd_sc_hd__and4_1
X_08713_ net538 _04897_ vssd1 vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__nor2_2
X_05925_ top.WB.CPU_DAT_O\[30\] net1173 net305 vssd1 vssd1 vccd1 vccd1 _02264_ sky130_fd_sc_hd__mux2_1
X_09693_ net800 net640 vssd1 vssd1 vccd1 vccd1 _00307_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout276_A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08644_ net1609 _04850_ vssd1 vssd1 vccd1 vccd1 _01497_ sky130_fd_sc_hd__xnor2_1
X_05856_ top.compVal\[11\] net170 net156 top.WB.CPU_DAT_O\[11\] vssd1 vssd1 vccd1
+ vccd1 _02286_ sky130_fd_sc_hd__a22o_1
XANTENNA__05706__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08575_ net1149 net517 net234 vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__mux2_1
X_05787_ top.findLeastValue.least1\[8\] top.findLeastValue.least2\[8\] vssd1 vssd1
+ vccd1 vccd1 _02807_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_1_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07526_ top.cb_syn.char_path_n\[112\] top.cb_syn.char_path_n\[111\] top.cb_syn.char_path_n\[110\]
+ top.cb_syn.char_path_n\[109\] net400 net351 vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout443_A net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout708_A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07457_ _04046_ _04047_ vssd1 vssd1 vccd1 vccd1 _04048_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout231_X net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout329_X net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07388_ _03988_ _03989_ _03987_ vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__mux2_1
XANTENNA__08959__A0 top.WB.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06408_ net1667 net299 _03242_ vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__a21o_1
XFILLER_108_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09127_ top.sram_interface.CB_write_counter\[1\] _02452_ net479 net541 _02690_ vssd1
+ vssd1 vccd1 vccd1 _05141_ sky130_fd_sc_hd__a41o_1
X_06339_ net1420 _03200_ net302 vssd1 vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__mux2_1
X_09058_ net454 _02405_ vssd1 vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__nor2_1
X_08009_ _04511_ vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_75_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold560 top.histogram.total\[21\] vssd1 vssd1 vccd1 vccd1 net1513 sky130_fd_sc_hd__dlygate4sd3_1
Xhold571 top.histogram.total\[4\] vssd1 vssd1 vccd1 vccd1 net1524 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold582 top.hTree.state\[5\] vssd1 vssd1 vccd1 vccd1 net1535 sky130_fd_sc_hd__dlygate4sd3_1
X_11020_ clknet_leaf_21_clk _01568_ _00375_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_9_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold593 top.hTree.tree_reg\[9\] vssd1 vssd1 vccd1 vccd1 net1546 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05945__A0 top.WB.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_TAPCELL_ROW_28_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11853_ clknet_leaf_116_clk _02369_ _01208_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[31\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_17_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10804_ clknet_leaf_48_clk _01390_ _00223_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.max_index\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_56_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11784_ clknet_leaf_72_clk _00019_ _01139_ vssd1 vssd1 vccd1 vccd1 top.hTree.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10735_ clknet_leaf_119_clk _01334_ _00154_ vssd1 vssd1 vccd1 vccd1 top.path\[111\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10666_ clknet_leaf_116_clk _01265_ _00085_ vssd1 vssd1 vccd1 vccd1 top.path\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10597_ net841 net681 vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__and2_1
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 STB_O sky130_fd_sc_hd__buf_2
XANTENNA_output72_A net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11218_ clknet_leaf_24_clk _01766_ _00573_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[120\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_95_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput91 net91 vssd1 vssd1 vccd1 vccd1 DAT_O[26] sky130_fd_sc_hd__buf_2
X_11149_ clknet_leaf_21_clk _01697_ _00504_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[51\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 DAT_O[16] sky130_fd_sc_hd__buf_2
XANTENNA__05936__A0 top.WB.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__09127__B1 _02690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09142__A3 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06690_ _02436_ top.findLeastValue.val2\[13\] vssd1 vssd1 vccd1 vccd1 _03478_ sky130_fd_sc_hd__nor2_1
X_05710_ net3 net417 net359 top.WB.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1 _02348_
+ sky130_fd_sc_hd__a22o_1
XFILLER_63_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05641_ net1411 net145 _02722_ net177 vssd1 vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__a22o_1
X_08360_ net438 _04705_ _04708_ net505 vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__o211a_1
XFILLER_17_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05572_ net457 top.hTree.node_reg\[50\] net361 net420 top.hTree.node_reg\[18\] vssd1
+ vssd1 vccd1 vccd1 _02665_ sky130_fd_sc_hd__a32o_1
XFILLER_51_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07311_ _03785_ _03940_ vssd1 vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__or2_1
X_08291_ top.cb_syn.char_path_n\[24\] net383 net342 top.cb_syn.char_path_n\[22\] net187
+ vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__a221o_1
X_07242_ _03822_ _03827_ _03889_ vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__or3b_1
X_07173_ _03828_ _03829_ _03830_ vssd1 vssd1 vccd1 vccd1 _03831_ sky130_fd_sc_hd__or3_1
X_06124_ top.cw1\[6\] _02995_ vssd1 vssd1 vccd1 vccd1 _02996_ sky130_fd_sc_hd__and2_1
XANTENNA__08821__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06967__A2 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06055_ net1363 net141 _02940_ net159 vssd1 vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__a22o_1
Xfanout303 _03171_ vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__buf_2
Xfanout314 net315 vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06341__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout347 net348 vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__clkbuf_2
Xfanout336 net349 vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__clkbuf_2
X_09814_ net742 net582 vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_6_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout358 _02926_ vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__clkbuf_2
Xfanout369 net370 vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05927__A0 top.WB.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout560_A top.sram_interface.word_cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09745_ net788 net628 vssd1 vssd1 vccd1 vccd1 _00359_ sky130_fd_sc_hd__and2_1
X_06957_ top.findLeastValue.val2\[5\] net151 net122 _03620_ vssd1 vssd1 vccd1 vccd1
+ _01947_ sky130_fd_sc_hd__o22a_1
XFILLER_27_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09676_ net799 net639 vssd1 vssd1 vccd1 vccd1 _00290_ sky130_fd_sc_hd__and2_1
X_05908_ top.sram_interface.CB_write_counter\[0\] _02561_ _02880_ vssd1 vssd1 vccd1
+ vccd1 _02881_ sky130_fd_sc_hd__o21ai_1
X_06888_ top.compVal\[39\] top.findLeastValue.val1\[39\] net166 vssd1 vssd1 vccd1
+ vccd1 _03586_ sky130_fd_sc_hd__mux2_1
XFILLER_39_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08627_ _04830_ _04835_ _04841_ _04826_ net1688 vssd1 vssd1 vccd1 vccd1 _01502_ sky130_fd_sc_hd__a32o_1
X_05839_ top.compVal\[28\] net171 net157 top.WB.CPU_DAT_O\[28\] vssd1 vssd1 vccd1
+ vccd1 _02303_ sky130_fd_sc_hd__a22o_1
XFILLER_54_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout446_X net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout825_A net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08558_ net1312 top.cb_syn.char_path_n\[18\] net222 vssd1 vssd1 vccd1 vccd1 _01536_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07527__S0 _04072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07900__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07509_ top.cb_syn.char_path_n\[92\] top.cb_syn.char_path_n\[91\] top.cb_syn.char_path_n\[90\]
+ top.cb_syn.char_path_n\[89\] net402 net353 vssd1 vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__mux4_1
X_08489_ net1254 top.cb_syn.char_path_n\[87\] net230 vssd1 vssd1 vccd1 vccd1 _01605_
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10520_ net861 net701 vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__and2_1
XFILLER_52_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10451_ net748 net588 vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__and2_1
XFILLER_108_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10382_ net854 net694 vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__and2_1
XANTENNA__08801__C1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold390 top.path\[125\] vssd1 vssd1 vccd1 vccd1 net1343 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09357__B1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05630__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11003_ clknet_leaf_17_clk _01551_ _00358_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[33\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout870 net877 vssd1 vssd1 vccd1 vccd1 net870 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_88_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_82_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__07518__S0 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11836_ clknet_leaf_100_clk _02352_ _01191_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_14_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__07810__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_97_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11767_ clknet_leaf_102_clk _02300_ _01122_ vssd1 vssd1 vccd1 vccd1 top.compVal\[25\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__05449__A2 _02555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07843__B1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10718_ clknet_leaf_2_clk _01317_ _00137_ vssd1 vssd1 vccd1 vccd1 top.path\[94\]
+ sky130_fd_sc_hd__dfrtp_1
X_11698_ clknet_leaf_61_clk _02231_ _01053_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_99_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10649_ clknet_leaf_60_clk _01248_ _00068_ vssd1 vssd1 vccd1 vccd1 top.hist_addr\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_20_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08399__A1 top.cb_syn.char_path_n\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06949__A2 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_35_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09348__B1 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07860_ top.hTree.tree_reg\[16\] top.findLeastValue.sum\[16\] net249 vssd1 vssd1
+ vccd1 vccd1 _04394_ sky130_fd_sc_hd__mux2_1
XANTENNA__07374__A2 _03553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07791_ net486 _04337_ vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__or2_1
XANTENNA__09325__X top.translation.writeBin vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06811_ top.findLeastValue.val1\[19\] net128 net112 top.compVal\[19\] vssd1 vssd1
+ vccd1 vccd1 _02027_ sky130_fd_sc_hd__o22a_1
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_06742_ _02415_ top.findLeastValue.val2\[33\] vssd1 vssd1 vccd1 vccd1 _03530_ sky130_fd_sc_hd__and2_1
X_09530_ net749 net589 vssd1 vssd1 vccd1 vccd1 _00144_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_108_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09461_ net751 net591 vssd1 vssd1 vccd1 vccd1 _00075_ sky130_fd_sc_hd__and2_1
X_06673_ top.compVal\[1\] top.findLeastValue.val2\[1\] vssd1 vssd1 vccd1 vccd1 _03461_
+ sky130_fd_sc_hd__and2b_1
XFILLER_36_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08412_ top.cb_syn.char_path_n\[21\] net392 net331 top.cb_syn.char_path_n\[22\] net506
+ vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__a221o_1
X_09392_ net407 _04251_ vssd1 vssd1 vccd1 vccd1 _05272_ sky130_fd_sc_hd__nand2_1
X_05624_ top.cb_syn.char_path\[73\] net552 net542 top.cb_syn.char_path\[41\] vssd1
+ vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout141_A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07509__S0 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08343_ top.cb_syn.char_path_n\[91\] top.cb_syn.char_path_n\[92\] net516 vssd1 vssd1
+ vccd1 vccd1 _04702_ sky130_fd_sc_hd__mux2_1
X_05555_ top.histogram.sram_out\[21\] net364 _02649_ _02650_ vssd1 vssd1 vccd1 vccd1
+ _02651_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_50_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07720__S net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08274_ top.cb_syn.char_path_n\[32\] net208 _04664_ vssd1 vssd1 vccd1 vccd1 _01678_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__07834__A0 top.findLeastValue.sum\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_108_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05486_ _02544_ _02593_ net177 vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__a21o_1
X_07225_ _03832_ _03836_ _03671_ vssd1 vssd1 vccd1 vccd1 _03877_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout406_A net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06860__A net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05860__A2 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07156_ _03795_ _03810_ _03813_ _03798_ vssd1 vssd1 vccd1 vccd1 _03814_ sky130_fd_sc_hd__o2bb2a_1
X_06107_ _02955_ _02969_ _02979_ vssd1 vssd1 vccd1 vccd1 _02980_ sky130_fd_sc_hd__or3_1
X_07087_ top.findLeastValue.val1\[4\] top.findLeastValue.val2\[4\] vssd1 vssd1 vccd1
+ vccd1 _03745_ sky130_fd_sc_hd__or2_1
X_06038_ top.cb_syn.cb_length\[6\] top.cb_syn.cb_length\[5\] _02928_ vssd1 vssd1 vccd1
+ vccd1 _02929_ sky130_fd_sc_hd__or3_1
XFILLER_0_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05612__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout775_A net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout122 net124 vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__clkbuf_4
Xfanout144 net145 vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__buf_2
XFILLER_59_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout133 _03444_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__buf_2
Xfanout155 net157 vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__clkbuf_4
Xfanout177 _02589_ vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__clkbuf_8
Xfanout188 net194 vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__clkbuf_2
Xfanout199 net203 vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__buf_2
Xfanout166 _03423_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__clkbuf_2
X_07989_ _04483_ _04491_ vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__nand2_1
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09728_ net739 net579 vssd1 vssd1 vccd1 vccd1 _00342_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09659_ net785 net625 vssd1 vssd1 vccd1 vccd1 _00273_ sky130_fd_sc_hd__and2_1
XFILLER_55_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05679__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ clknet_leaf_64_clk _02169_ _00976_ vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__dfrtp_1
XFILLER_23_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11552_ clknet_leaf_123_clk _02100_ _00907_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10503_ net809 net649 vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__and2_1
X_11483_ clknet_leaf_98_clk _02031_ _00838_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[23\]
+ sky130_fd_sc_hd__dfstp_1
X_10434_ net873 net713 vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__and2_1
XANTENNA__05851__A2 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10365_ net853 net693 vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_94_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05603__A2 _02689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10296_ net723 net563 vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__and2_1
Xteam_05_950 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] team_05_950/LO sky130_fd_sc_hd__conb_1
XANTENNA__07805__S net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05833__B _02843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06648__C top.compVal\[33\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06867__A1 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11819_ clknet_leaf_56_clk _02335_ _01174_ vssd1 vssd1 vccd1 vccd1 top.TRN_char_index\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_16_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05340_ top.compVal\[0\] vssd1 vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__inv_2
XFILLER_21_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06619__A1 top.compVal\[33\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07292__A1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07292__B2 top.findLeastValue.sum\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07010_ _03666_ _03667_ vssd1 vssd1 vccd1 vccd1 _03668_ sky130_fd_sc_hd__nor2_1
XANTENNA__05842__A2 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05296__A net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08961_ top.WB.CPU_DAT_O\[31\] net1320 net321 vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__mux2_1
XFILLER_102_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08892_ _02795_ net492 top.findLeastValue.least1\[8\] top.hTree.write_HT_fin vssd1
+ vssd1 vccd1 vccd1 _05062_ sky130_fd_sc_hd__and4b_1
X_07912_ net426 _04434_ _04435_ net258 vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__o211a_1
XANTENNA__08544__A1 top.cb_syn.char_path_n\[32\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07843_ net441 net1554 net253 net1725 _04380_ vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__a221o_1
XFILLER_56_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05583__X _02674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07715__S net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_3_Left_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09215__B top.controller.fin_reg\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07774_ top.findLeastValue.sum\[33\] top.hTree.tree_reg\[33\] net280 vssd1 vssd1
+ vccd1 vccd1 _04325_ sky130_fd_sc_hd__mux2_1
XFILLER_83_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09513_ net733 net573 vssd1 vssd1 vccd1 vccd1 _00127_ sky130_fd_sc_hd__and2_1
X_06725_ net494 _02487_ top.findLeastValue.val2\[26\] _02424_ vssd1 vssd1 vccd1 vccd1
+ _03513_ sky130_fd_sc_hd__a22o_1
X_06656_ top.cw1\[7\] net135 vssd1 vssd1 vccd1 vccd1 _02072_ sky130_fd_sc_hd__and2_1
X_09444_ net860 net700 vssd1 vssd1 vccd1 vccd1 _00058_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout356_A _02926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06855__A net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05607_ top.cb_syn.char_path\[12\] net557 net312 top.cb_syn.char_path\[108\] vssd1
+ vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout144_X net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06587_ _02438_ top.findLeastValue.val1\[11\] vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__and2_1
X_09375_ net1293 net236 net214 _04286_ vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__a22o_1
X_05538_ net1406 net140 _02636_ net175 vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__a22o_1
X_08326_ top.cb_syn.char_path_n\[6\] net199 _04690_ vssd1 vssd1 vccd1 vccd1 _01652_
+ sky130_fd_sc_hd__o21a_1
X_05469_ _02562_ net316 vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout311_X net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_49_Left_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08257_ top.cb_syn.char_path_n\[41\] net378 net337 top.cb_syn.char_path_n\[39\] net182
+ vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__a221o_1
XFILLER_20_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_08188_ top.cb_syn.char_path_n\[75\] net199 _04621_ vssd1 vssd1 vccd1 vccd1 _01721_
+ sky130_fd_sc_hd__o21a_1
X_07208_ _03855_ _03857_ _03859_ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__and3_1
X_07139_ _03795_ _03796_ vssd1 vssd1 vccd1 vccd1 _03797_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10150_ net815 net655 vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__and2_1
XANTENNA__06794__B1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10081_ net864 net704 vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__and2_1
XFILLER_58_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_58_Left_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08535__A1 top.cb_syn.char_path_n\[41\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09406__A net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11444__Q top.findLeastValue.histo_index\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10983_ clknet_leaf_5_clk _01531_ _00338_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11604_ clknet_leaf_56_clk _02152_ _00959_ vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_67_Left_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11535_ clknet_leaf_1_clk _02083_ _00890_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05668__X _02745_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11466_ clknet_leaf_95_clk _02014_ _00821_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[6\]
+ sky130_fd_sc_hd__dfstp_2
X_10417_ net870 net710 vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__and2_1
XANTENNA__08223__B1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11397_ clknet_leaf_93_clk _01945_ _00752_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[3\]
+ sky130_fd_sc_hd__dfstp_1
X_10348_ net870 net710 vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__and2_1
XANTENNA__06785__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_76_Left_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10279_ net726 net566 vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__and2_1
XANTENNA__06537__B1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07490_ top.cb_syn.char_path_n\[8\] top.cb_syn.char_path_n\[7\] top.cb_syn.char_path_n\[6\]
+ top.cb_syn.char_path_n\[5\] net399 net350 vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__mux4_1
XANTENNA__05760__B2 top.WB.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06510_ _03308_ _03310_ vssd1 vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__nor2_1
X_06441_ top.header_synthesis.count\[0\] _03245_ top.header_synthesis.count\[1\] vssd1
+ vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__a21o_1
XANTENNA__06304__A3 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05512__A1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09160_ net449 net295 top.histogram.state\[0\] vssd1 vssd1 vccd1 vccd1 _05163_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_64_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06372_ _03185_ _03219_ net301 vssd1 vssd1 vccd1 vccd1 _03220_ sky130_fd_sc_hd__and3b_1
X_09091_ net459 net468 vssd1 vssd1 vccd1 vccd1 _05111_ sky130_fd_sc_hd__or2_1
X_08111_ top.cb_syn.char_path_n\[114\] net375 net335 top.cb_syn.char_path_n\[112\]
+ net180 vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__a221o_1
X_05323_ top.compVal\[18\] vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__inv_2
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08042_ net535 _04535_ vssd1 vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_116_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09993_ net848 net688 vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__and2_1
XFILLER_103_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08944_ top.WB.CPU_DAT_O\[29\] top.cb_syn.h_element\[61\] net369 vssd1 vssd1 vccd1
+ vccd1 _01366_ sky130_fd_sc_hd__mux2_1
XANTENNA__06776__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08875_ net437 _05047_ _05051_ vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout473_A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07826_ net485 _04365_ vssd1 vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout640_A net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07757_ net429 _04310_ _04311_ net260 vssd1 vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout261_X net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout359_X net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06708_ _03494_ _03495_ vssd1 vssd1 vccd1 vccd1 _03496_ sky130_fd_sc_hd__nand2_1
XANTENNA__05751__B2 top.WB.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07688_ _02476_ net396 _04255_ vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__o21a_1
XFILLER_52_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09427_ net1013 net245 _05294_ vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__o21a_1
X_06639_ top.compVal\[3\] top.compVal\[2\] top.compVal\[1\] top.compVal\[0\] vssd1
+ vssd1 vccd1 vccd1 _03428_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout526_X net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09358_ net1532 net239 net216 _04354_ vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__a22o_1
X_08309_ top.cb_syn.char_path_n\[15\] net374 net334 top.cb_syn.char_path_n\[13\] net178
+ vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__a221o_1
X_09289_ _04006_ _05232_ _04019_ vssd1 vssd1 vccd1 vccd1 top.dut.bit_buf_next\[5\]
+ sky130_fd_sc_hd__o21a_1
X_11320_ clknet_leaf_75_clk _01868_ _00675_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_119_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11251_ clknet_leaf_49_clk _01799_ _00606_ vssd1 vssd1 vccd1 vccd1 top.hTree.nullSumIndex\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11182_ clknet_leaf_20_clk _01730_ _00537_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[84\]
+ sky130_fd_sc_hd__dfrtp_1
X_10202_ net831 net671 vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__and2_1
XANTENNA__08756__A1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10133_ net836 net676 vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__and2_1
XFILLER_0_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA_input34_A en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10064_ net860 net700 vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__and2_1
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10966_ clknet_leaf_40_clk _01514_ _00321_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_index\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06298__A2 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08692__B1 _04875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10897_ clknet_leaf_52_clk top.header_synthesis.next_header\[2\] _00252_ vssd1 vssd1
+ vccd1 vccd1 top.header_synthesis.header\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_43_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08914__S _05072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11518_ clknet_leaf_67_clk _02066_ _00873_ vssd1 vssd1 vccd1 vccd1 top.cw1\[1\] sky130_fd_sc_hd__dfrtp_2
Xhold208 top.cb_syn.char_path\[89\] vssd1 vssd1 vccd1 vccd1 net1161 sky130_fd_sc_hd__dlygate4sd3_1
X_11449_ clknet_leaf_69_clk _01997_ _00804_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.histo_index\[8\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold219 top.path\[29\] vssd1 vssd1 vccd1 vccd1 net1172 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_84_Left_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08747__A1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11349__Q top.findLeastValue.sum\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06990_ top.findLeastValue.val1\[46\] top.findLeastValue.val1\[45\] top.findLeastValue.val1\[44\]
+ top.findLeastValue.val1\[43\] vssd1 vssd1 vccd1 vccd1 _03648_ sky130_fd_sc_hd__and4_1
X_05941_ top.WB.CPU_DAT_O\[14\] net1380 net306 vssd1 vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__mux2_1
X_05872_ top.sram_interface.init_counter\[11\] _02847_ _02848_ _02850_ vssd1 vssd1
+ vccd1 vccd1 _02851_ sky130_fd_sc_hd__and4bb_1
X_08660_ net530 net529 _02858_ _04480_ vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__or4_1
XFILLER_93_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07611_ net445 top.WorR _04192_ _04193_ vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__a211o_1
X_08591_ _04814_ top.cb_syn.char_index\[1\] _04807_ vssd1 vssd1 vccd1 vccd1 _01511_
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_93_Left_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07542_ net535 net540 vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__nor2_1
XANTENNA__08683__B1 _04875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07473_ _04044_ _04063_ vssd1 vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__or2_1
X_06424_ net1644 _03249_ _03250_ vssd1 vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__o21a_1
X_09212_ top.controller.fin_reg\[1\] top.controller.fin_reg\[4\] top.controller.fin_reg\[3\]
+ top.controller.fin_reg\[2\] vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__or4bb_1
XANTENNA__08824__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_09143_ _05152_ _05151_ _05088_ vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__or3b_1
X_06355_ _03190_ _03208_ vssd1 vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__nor2_1
XANTENNA__06852__B net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout221_A net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout319_A net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05306_ top.compVal\[34\] vssd1 vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__inv_2
X_09074_ net474 _04130_ _04866_ vssd1 vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__and3_1
X_06286_ top.cw2\[1\] top.cw2\[0\] vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__or2_1
X_08025_ top.cb_syn.count\[3\] _04511_ vssd1 vssd1 vccd1 vccd1 _04524_ sky130_fd_sc_hd__or2_1
XANTENNA__05468__B _02555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold720 top.compVal\[23\] vssd1 vssd1 vccd1 vccd1 net1673 sky130_fd_sc_hd__dlygate4sd3_1
Xhold764 top.sram_interface.init_counter\[2\] vssd1 vssd1 vccd1 vccd1 net1717 sky130_fd_sc_hd__dlygate4sd3_1
Xhold742 _01895_ vssd1 vssd1 vccd1 vccd1 net1695 sky130_fd_sc_hd__dlygate4sd3_1
Xhold753 top.cb_syn.char_path_n\[90\] vssd1 vssd1 vccd1 vccd1 net1706 sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 top.findLeastValue.sum\[0\] vssd1 vssd1 vccd1 vccd1 net1684 sky130_fd_sc_hd__dlygate4sd3_1
Xhold775 top.sram_interface.init_counter\[10\] vssd1 vssd1 vccd1 vccd1 net1728 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout688_A net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout590_A net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09976_ net780 net620 vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__and2_1
XANTENNA__10390__A net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout855_A net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08927_ top.WB.CPU_DAT_O\[27\] net1340 net372 vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout476_X net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09163__A1 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08858_ _02786_ _04925_ _02785_ vssd1 vssd1 vccd1 vccd1 _05040_ sky130_fd_sc_hd__o21bai_2
X_07809_ top.findLeastValue.sum\[26\] top.hTree.tree_reg\[26\] net278 vssd1 vssd1
+ vccd1 vccd1 _04353_ sky130_fd_sc_hd__mux2_1
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08789_ top.translation.index\[2\] _04959_ _04962_ top.translation.index\[4\] vssd1
+ vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_43_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10820_ clknet_leaf_109_clk _01406_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10751_ clknet_leaf_2_clk _01350_ _00170_ vssd1 vssd1 vccd1 vccd1 top.path\[127\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05488__B1 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10682_ clknet_leaf_120_clk _01281_ _00101_ vssd1 vssd1 vccd1 vccd1 top.path\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08426__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11303_ clknet_leaf_77_clk _01851_ _00658_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[46\]
+ sky130_fd_sc_hd__dfrtp_1
X_11234_ clknet_leaf_38_clk _01782_ _00589_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.left
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05660__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11165_ clknet_leaf_17_clk _01713_ _00520_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[67\]
+ sky130_fd_sc_hd__dfrtp_1
X_11096_ clknet_leaf_28_clk _01644_ _00451_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[126\]
+ sky130_fd_sc_hd__dfrtp_1
X_10116_ net820 net660 vssd1 vssd1 vccd1 vccd1 _00730_ sky130_fd_sc_hd__and2_1
X_10047_ net858 net698 vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__and2_1
XFILLER_48_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold91 net54 vssd1 vssd1 vccd1 vccd1 net1044 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08901__A1 _03325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold80 top.hTree.node_reg\[42\] vssd1 vssd1 vccd1 vccd1 net1033 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05715__B2 top.WB.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10949_ clknet_leaf_37_clk _01504_ _00304_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.num_lefts\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_70_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__10475__A net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05494__A3 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06140_ net503 net504 vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__nand2_1
X_06071_ top.sram_interface.init_counter\[6\] _02945_ vssd1 vssd1 vccd1 vccd1 _02946_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_113_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08599__B top.CB_read_complete vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout518 net519 vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__clkbuf_4
Xfanout529 top.cb_syn.curr_state\[8\] vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__buf_2
Xfanout507 net508 vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__buf_2
X_09830_ net770 net610 vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__and2_1
XFILLER_112_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09761_ net773 net613 vssd1 vssd1 vccd1 vccd1 _00375_ sky130_fd_sc_hd__and2_1
X_06973_ top.findLeastValue.val2\[26\] top.findLeastValue.val2\[25\] top.findLeastValue.val2\[24\]
+ top.findLeastValue.val2\[23\] vssd1 vssd1 vccd1 vccd1 _03631_ sky130_fd_sc_hd__and4_1
X_08712_ net538 _04903_ _04898_ vssd1 vssd1 vccd1 vccd1 _04904_ sky130_fd_sc_hd__o21bai_1
X_05924_ top.WB.CPU_DAT_O\[31\] net1237 net304 vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__mux2_1
X_09692_ net799 net639 vssd1 vssd1 vccd1 vccd1 _00306_ sky130_fd_sc_hd__and2_1
XANTENNA__05591__X _02681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08353__C1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08643_ net1645 _04853_ vssd1 vssd1 vccd1 vccd1 _01498_ sky130_fd_sc_hd__xor2_1
XANTENNA__05706__B2 top.WB.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05855_ top.compVal\[12\] net168 net154 top.WB.CPU_DAT_O\[12\] vssd1 vssd1 vccd1
+ vccd1 _02287_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout171_A _02845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06903__B1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06339__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05786_ top.sram_interface.counter_HTREE\[0\] _02804_ vssd1 vssd1 vccd1 vccd1 _02806_
+ sky130_fd_sc_hd__nor2_1
X_08574_ net1153 top.cb_syn.char_path_n\[2\] net234 vssd1 vssd1 vccd1 vccd1 _01520_
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout269_A _03864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07525_ top.cb_syn.char_path_n\[108\] top.cb_syn.char_path_n\[107\] top.cb_syn.char_path_n\[106\]
+ top.cb_syn.char_path_n\[105\] net400 net351 vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__mux4_1
XFILLER_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_61_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08751__S0 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout436_A _02523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08120__A2 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07456_ top.cb_syn.cb_length\[4\] top.cb_syn.i\[4\] vssd1 vssd1 vccd1 vccd1 _04047_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07387_ top.dut.bit_buf\[9\] top.dut.bit_buf\[2\] net721 vssd1 vssd1 vccd1 vccd1
+ _03989_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout224_X net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout603_A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06407_ _03174_ _03241_ net300 vssd1 vssd1 vccd1 vccd1 _03242_ sky130_fd_sc_hd__and3b_1
X_09126_ net450 top.sram_interface.word_cnt\[9\] _05111_ _05140_ vssd1 vssd1 vccd1
+ vccd1 _00049_ sky130_fd_sc_hd__a31o_1
X_06338_ top.hist_data_o\[30\] _03199_ _03194_ vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__o21ba_1
X_06269_ top.cw1\[1\] top.cw1\[0\] top.cw1\[2\] vssd1 vssd1 vccd1 vccd1 _03135_ sky130_fd_sc_hd__a21o_1
X_09057_ net1201 top.WB.CPU_DAT_O\[0\] net294 vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__mux2_1
X_08008_ top.cb_syn.count\[2\] top.cb_syn.count\[1\] top.cb_syn.count\[0\] vssd1 vssd1
+ vccd1 vccd1 _04511_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_75_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05642__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold572 top.hTree.tree_reg\[45\] vssd1 vssd1 vccd1 vccd1 net1525 sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 _03301_ vssd1 vssd1 vccd1 vccd1 net1514 sky130_fd_sc_hd__dlygate4sd3_1
Xhold550 top.histogram.total\[5\] vssd1 vssd1 vccd1 vccd1 net1503 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold594 top.hTree.nullSumIndex\[6\] vssd1 vssd1 vccd1 vccd1 net1547 sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 top.hTree.tree_reg\[30\] vssd1 vssd1 vccd1 vccd1 net1536 sky130_fd_sc_hd__dlygate4sd3_1
X_09959_ net771 net611 vssd1 vssd1 vccd1 vccd1 _00573_ sky130_fd_sc_hd__and2_1
XANTENNA__08344__C1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ clknet_leaf_17_clk _02368_ _01207_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[30\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08647__B1 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10803_ clknet_leaf_48_clk _01389_ _00222_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.max_index\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_56_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_52_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_clk sky130_fd_sc_hd__clkbuf_8
X_11783_ clknet_leaf_73_clk _00017_ _01138_ vssd1 vssd1 vccd1 vccd1 top.hTree.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_10734_ clknet_leaf_119_clk _01333_ _00153_ vssd1 vssd1 vccd1 vccd1 top.path\[110\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05476__A3 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10665_ clknet_leaf_118_clk _01264_ _00084_ vssd1 vssd1 vccd1 vccd1 top.path\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07622__A1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10596_ net808 net648 vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__and2_1
XANTENNA__07622__B2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05676__X _02752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 ADR_O[8] sky130_fd_sc_hd__buf_2
X_11217_ clknet_leaf_24_clk _01765_ _00572_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[119\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08178__A2 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput92 net92 vssd1 vssd1 vccd1 vccd1 DAT_O[27] sky130_fd_sc_hd__buf_2
X_11148_ clknet_leaf_22_clk _01696_ _00503_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[50\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 DAT_O[17] sky130_fd_sc_hd__buf_2
XFILLER_0_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08335__C1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11079_ clknet_leaf_5_clk _01627_ _00434_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[109\]
+ sky130_fd_sc_hd__dfrtp_1
X_05640_ top.histogram.sram_out\[7\] net363 net419 top.hTree.node_reg\[7\] _02721_
+ vssd1 vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__a221o_1
XFILLER_63_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05571_ _02662_ _02663_ net472 vssd1 vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__o21a_1
XFILLER_51_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_43_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_clk sky130_fd_sc_hd__clkbuf_8
X_07310_ top.findLeastValue.val1\[16\] top.findLeastValue.val2\[16\] _03920_ vssd1
+ vssd1 vccd1 vccd1 _03940_ sky130_fd_sc_hd__a21o_1
XFILLER_17_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08290_ top.cb_syn.char_path_n\[24\] net204 _04672_ vssd1 vssd1 vccd1 vccd1 _01670_
+ sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_9_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07241_ _03824_ _03888_ vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__nand2_1
X_07172_ top.findLeastValue.val1\[33\] top.findLeastValue.val2\[33\] vssd1 vssd1 vccd1
+ vccd1 _03830_ sky130_fd_sc_hd__xnor2_1
X_06123_ top.cw1\[5\] top.cw1\[4\] _02993_ vssd1 vssd1 vccd1 vccd1 _02995_ sky130_fd_sc_hd__and3_1
XFILLER_8_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05624__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06054_ net454 net466 net461 _02939_ vssd1 vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__or4_1
XANTENNA__08169__A2 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout304 net305 vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__clkbuf_4
Xfanout315 net316 vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__buf_2
Xfanout348 net349 vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__clkbuf_2
Xfanout337 net349 vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__buf_2
X_09813_ net760 net600 vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__and2_1
Xfanout326 net329 vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout386_A net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout359 net360 vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08549__S net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06858__A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09744_ net788 net628 vssd1 vssd1 vccd1 vccd1 _00358_ sky130_fd_sc_hd__and2_1
X_06956_ top.compVal\[5\] top.findLeastValue.val1\[5\] net166 vssd1 vssd1 vccd1 vccd1
+ _03620_ sky130_fd_sc_hd__mux2_1
X_09675_ net797 net637 vssd1 vssd1 vccd1 vccd1 _00289_ sky130_fd_sc_hd__and2_1
X_05907_ _02529_ net478 _02562_ _02857_ _02875_ vssd1 vssd1 vccd1 vccd1 _02880_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout553_A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout174_X net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06887_ top.findLeastValue.val2\[40\] net150 net123 _03585_ vssd1 vssd1 vccd1 vccd1
+ _01982_ sky130_fd_sc_hd__o22a_1
X_08626_ top.cb_syn.num_lefts\[2\] top.cb_syn.num_lefts\[1\] top.cb_syn.num_lefts\[0\]
+ top.cb_syn.num_lefts\[3\] vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__a31o_1
XANTENNA__08341__A2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05838_ top.compVal\[29\] net169 net155 top.WB.CPU_DAT_O\[29\] vssd1 vssd1 vccd1
+ vccd1 _02304_ sky130_fd_sc_hd__a22o_1
XFILLER_54_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08629__B1 _04826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout439_X net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_34_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout341_X net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08557_ net1179 top.cb_syn.char_path_n\[19\] net222 vssd1 vssd1 vccd1 vccd1 _01537_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05769_ top.translation.index\[6\] top.translation.index\[5\] _02789_ vssd1 vssd1
+ vccd1 vccd1 _02790_ sky130_fd_sc_hd__nor3_1
X_08488_ net1236 top.cb_syn.char_path_n\[88\] net230 vssd1 vssd1 vccd1 vccd1 _01606_
+ sky130_fd_sc_hd__mux2_1
X_07508_ top.cb_syn.char_path_n\[88\] top.cb_syn.char_path_n\[87\] top.cb_syn.char_path_n\[86\]
+ top.cb_syn.char_path_n\[85\] net401 net353 vssd1 vssd1 vccd1 vccd1 _04099_ sky130_fd_sc_hd__mux4_1
XANTENNA__07527__S1 _04071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07439_ top.dut.bit_buf\[2\] net40 net721 vssd1 vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10450_ net746 net586 vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__and2_1
XANTENNA__05863__B1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09109_ net463 _05112_ top.sram_interface.word_cnt\[2\] vssd1 vssd1 vccd1 vccd1 _05128_
+ sky130_fd_sc_hd__o21ai_1
X_10381_ net855 net695 vssd1 vssd1 vccd1 vccd1 _00995_ sky130_fd_sc_hd__and2_1
XFILLER_108_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__09409__A net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07628__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold380 top.hTree.nulls\[49\] vssd1 vssd1 vccd1 vccd1 net1333 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07368__B1 _03553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08032__B top.CB_write_complete vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11002_ clknet_leaf_18_clk _01550_ _00357_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[32\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold391 top.path\[80\] vssd1 vssd1 vccd1 vccd1 net1344 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout860 net877 vssd1 vssd1 vccd1 vccd1 net860 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11447__Q top.findLeastValue.histo_index\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout871 net872 vssd1 vssd1 vccd1 vccd1 net871 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_88_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_25_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_60_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_11835_ clknet_leaf_121_clk _02351_ _01190_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07518__S1 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11766_ clknet_leaf_98_clk _02299_ _01121_ vssd1 vssd1 vccd1 vccd1 top.compVal\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07843__A1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10717_ clknet_leaf_3_clk _01316_ _00136_ vssd1 vssd1 vccd1 vccd1 top.path\[93\]
+ sky130_fd_sc_hd__dfrtp_1
X_11697_ clknet_leaf_61_clk _02230_ _01052_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_99_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05854__B1 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10648_ clknet_leaf_74_clk _00043_ _00067_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.word_cnt\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10579_ net729 net569 vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_11_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05606__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11357__Q top.findLeastValue.sum\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07790_ top.hTree.tree_reg\[30\] top.findLeastValue.sum\[30\] net248 vssd1 vssd1
+ vccd1 vccd1 _04338_ sky130_fd_sc_hd__mux2_1
X_06810_ top.findLeastValue.val1\[20\] net128 net112 top.compVal\[20\] vssd1 vssd1
+ vccd1 vccd1 _02028_ sky130_fd_sc_hd__o22a_1
X_06741_ _02414_ top.findLeastValue.val2\[34\] vssd1 vssd1 vccd1 vccd1 _03529_ sky130_fd_sc_hd__and2_1
X_09460_ net869 net709 vssd1 vssd1 vccd1 vccd1 _00074_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_108_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08411_ top.cb_syn.char_path_n\[23\] top.cb_syn.char_path_n\[24\] net515 vssd1 vssd1
+ vccd1 vccd1 _04770_ sky130_fd_sc_hd__mux2_1
X_06672_ top.compVal\[2\] top.findLeastValue.val2\[2\] vssd1 vssd1 vccd1 vccd1 _03460_
+ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_16_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_8
X_09391_ net980 net240 _05270_ _05271_ vssd1 vssd1 vccd1 vccd1 _01444_ sky130_fd_sc_hd__a22o_1
X_05623_ net1191 net140 _02707_ net174 vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__a22o_1
XANTENNA__06885__A2 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07509__S1 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08342_ top.cb_syn.char_path_n\[94\] net332 _04700_ vssd1 vssd1 vccd1 vccd1 _04701_
+ sky130_fd_sc_hd__a21oi_1
X_05554_ net456 top.hTree.node_reg\[53\] net361 net420 top.hTree.node_reg\[21\] vssd1
+ vssd1 vccd1 vccd1 _02650_ sky130_fd_sc_hd__a32o_1
XFILLER_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05485_ top.WB.curr_state\[0\] _02590_ vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__and2_1
X_08273_ top.cb_syn.char_path_n\[33\] net387 net346 top.cb_syn.char_path_n\[31\] net191
+ vssd1 vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout134_A net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07224_ net1627 net276 _03875_ _03876_ vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__a22o_1
XANTENNA__05845__B1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout301_A net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07155_ _03786_ _03789_ _03791_ _03812_ vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__o211a_1
X_06106_ _02973_ _02978_ top.TRN_char_index\[6\] _02566_ vssd1 vssd1 vccd1 vccd1 _02979_
+ sky130_fd_sc_hd__o211a_1
X_07086_ top.findLeastValue.val1\[4\] top.findLeastValue.val2\[4\] vssd1 vssd1 vccd1
+ vccd1 _03744_ sky130_fd_sc_hd__nand2_1
XANTENNA__08795__C1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06037_ top.cb_syn.cb_length\[4\] top.cb_syn.cb_length\[3\] top.cb_syn.cb_length\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02928_ sky130_fd_sc_hd__or3_1
Xfanout112 net113 vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__clkbuf_4
Xfanout145 _02595_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__clkbuf_8
Xfanout134 net136 vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__buf_2
Xfanout156 net157 vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__buf_2
Xfanout123 net124 vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__buf_2
X_07988_ _02513_ top.cb_syn.zero_count\[3\] vssd1 vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__or2_1
Xfanout189 net190 vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__buf_2
XANTENNA_fanout389_X net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout167 _03423_ vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__clkbuf_4
XFILLER_47_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout178 net179 vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_114_Right_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09727_ net739 net579 vssd1 vssd1 vccd1 vccd1 _00341_ sky130_fd_sc_hd__and2_1
X_06939_ top.findLeastValue.val2\[14\] net146 net121 _03611_ vssd1 vssd1 vccd1 vccd1
+ _01956_ sky130_fd_sc_hd__o22a_1
X_09658_ net803 net643 vssd1 vssd1 vccd1 vccd1 _00272_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_38_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08609_ top.cb_syn.num_lefts\[2\] top.cb_syn.num_lefts\[1\] top.cb_syn.num_lefts\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04828_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_83_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09589_ net822 net662 vssd1 vssd1 vccd1 vccd1 _00203_ sky130_fd_sc_hd__and2_1
X_11620_ clknet_leaf_62_clk _02168_ _00975_ vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__dfrtp_1
XFILLER_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07825__A1 top.findLeastValue.sum\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11551_ clknet_leaf_123_clk _02099_ _00906_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10502_ net753 net593 vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__and2_1
XFILLER_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05836__B1 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11482_ clknet_leaf_101_clk _02030_ _00837_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[22\]
+ sky130_fd_sc_hd__dfstp_1
X_10433_ net875 net715 vssd1 vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__and2_1
X_10364_ net865 net705 vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__and2_1
XFILLER_12_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10295_ net724 net564 vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__and2_1
XANTENNA__06800__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_05_951 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] team_05_951/LO sky130_fd_sc_hd__conb_1
Xteam_05_940 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] team_05_940/LO sky130_fd_sc_hd__conb_1
Xfanout690 net697 vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__clkbuf_2
XFILLER_93_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08917__S _05072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09602__A net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11818_ clknet_leaf_56_clk _02334_ _01173_ vssd1 vssd1 vccd1 vccd1 top.TRN_char_index\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_16_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11749_ clknet_leaf_95_clk _02282_ _01104_ vssd1 vssd1 vccd1 vccd1 top.compVal\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09018__A0 top.WB.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08960_ top.sram_interface.TRN_counter\[2\] _02889_ top.sram_interface.TRN_counter\[1\]
+ top.sram_interface.TRN_counter\[0\] vssd1 vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__or4b_4
Xclkbuf_leaf_5_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_8
X_08891_ net458 _02802_ _05060_ vssd1 vssd1 vccd1 vccd1 _05061_ sky130_fd_sc_hd__and3_1
XANTENNA__06900__S net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07911_ net483 _04433_ vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__or2_1
XFILLER_110_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07842_ net428 _04378_ _04379_ net262 vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__o211a_1
XFILLER_69_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09215__C top.controller.fin_reg\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07773_ net446 net1441 net254 net1727 _04324_ vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__a221o_1
X_09512_ net736 net576 vssd1 vssd1 vccd1 vccd1 _00126_ sky130_fd_sc_hd__and2_1
XANTENNA__06307__B2 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06724_ net494 _02487_ vssd1 vssd1 vccd1 vccd1 _03512_ sky130_fd_sc_hd__nand2_1
X_09443_ net856 net696 vssd1 vssd1 vccd1 vccd1 _00057_ sky130_fd_sc_hd__and2_1
X_06655_ net288 _03442_ vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_35_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09257__B1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06347__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09374_ net1033 net237 net214 _04290_ vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__a22o_1
X_05606_ top.cb_syn.char_path\[76\] net551 net542 top.cb_syn.char_path\[44\] vssd1
+ vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__a22o_1
X_08325_ top.cb_syn.char_path_n\[7\] net378 net337 top.cb_syn.char_path_n\[5\] net182
+ vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__a221o_1
X_06586_ _02437_ top.findLeastValue.val1\[12\] vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout137_X net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout516_A top.cb_syn.end_cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05537_ top.histogram.sram_out\[24\] net365 _02634_ _02635_ vssd1 vssd1 vccd1 vccd1
+ _02636_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_104_Left_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05468_ _02536_ _02555_ vssd1 vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__nor2_1
XFILLER_20_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09009__A0 top.WB.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07283__A2 _03658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08256_ top.cb_syn.char_path_n\[41\] net200 _04655_ vssd1 vssd1 vccd1 vccd1 _01687_
+ sky130_fd_sc_hd__o21a_1
X_07207_ _03862_ _03863_ net271 net276 net1548 vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__a32o_1
X_08187_ top.cb_syn.char_path_n\[76\] net378 net337 top.cb_syn.char_path_n\[74\] net182
+ vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__a221o_1
X_05399_ top.cb_syn.char_index\[3\] vssd1 vssd1 vccd1 vccd1 _02507_ sky130_fd_sc_hd__inv_2
X_07138_ top.findLeastValue.val1\[21\] top.findLeastValue.val2\[21\] vssd1 vssd1 vccd1
+ vccd1 _03796_ sky130_fd_sc_hd__nand2_1
XANTENNA__08768__C1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_81_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07069_ top.findLeastValue.val1\[10\] top.findLeastValue.val2\[10\] vssd1 vssd1 vccd1
+ vccd1 _03727_ sky130_fd_sc_hd__nand2_1
X_10080_ net852 net692 vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__and2_1
XFILLER_99_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_96_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Left_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold728_A top.findLeastValue.sum\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10982_ clknet_leaf_5_clk _01530_ _00337_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09141__B net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_34_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11603_ clknet_leaf_63_clk _02151_ _00958_ vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__dfrtp_1
XANTENNA__05521__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11534_ clknet_leaf_1_clk _02082_ _00889_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_49_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11465_ clknet_leaf_94_clk _02013_ _00820_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[5\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_11_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_10416_ net870 net710 vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__and2_1
XFILLER_99_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05397__A net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11396_ clknet_leaf_93_clk _01944_ _00751_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[2\]
+ sky130_fd_sc_hd__dfstp_1
X_10347_ net871 net711 vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__and2_1
XANTENNA__05588__A2 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05684__X _02758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10278_ net726 net566 vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_107_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_81_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06440_ _03257_ _03265_ vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__nor2_1
XANTENNA__10478__A net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06371_ top.hist_data_o\[15\] top.hist_data_o\[14\] _03184_ top.hist_data_o\[16\]
+ vssd1 vssd1 vccd1 vccd1 _03219_ sky130_fd_sc_hd__a31o_1
XFILLER_119_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_09090_ net459 net468 vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__nor2_1
X_08110_ top.cb_syn.char_path_n\[114\] net197 _04582_ vssd1 vssd1 vccd1 vccd1 _01760_
+ sky130_fd_sc_hd__o21a_1
X_05322_ top.compVal\[19\] vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__inv_2
X_08041_ _02862_ _04534_ vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_116_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_6_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09992_ net847 net687 vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__and2_1
XANTENNA__06776__A1 top.findLeastValue.least1\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05579__A2 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08943_ top.WB.CPU_DAT_O\[30\] net1476 net370 vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__mux2_1
XANTENNA__06776__B2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_15_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_15_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_69_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout299_A _03172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_08874_ net437 _05047_ _05043_ vssd1 vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout466_A top.controller.state_reg\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_07825_ top.hTree.tree_reg\[23\] top.findLeastValue.sum\[23\] net248 vssd1 vssd1
+ vccd1 vccd1 _04366_ sky130_fd_sc_hd__mux2_1
X_07756_ net493 _04309_ vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__or2_1
X_06707_ top.compVal\[21\] _02491_ _02492_ top.compVal\[20\] vssd1 vssd1 vccd1 vccd1
+ _03495_ sky130_fd_sc_hd__o22a_1
X_09426_ top.hTree.nulls\[63\] _02809_ net243 _05293_ vssd1 vssd1 vccd1 vccd1 _05294_
+ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout633_A net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07687_ net396 _04254_ vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__nand2_1
XFILLER_44_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10388__A net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_52_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06638_ top.compVal\[7\] top.compVal\[6\] top.compVal\[5\] top.compVal\[4\] vssd1
+ vssd1 vccd1 vccd1 _03427_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout800_A net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout421_X net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09357_ net1592 net239 net219 _04358_ vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__a22o_1
X_06569_ _02448_ top.findLeastValue.val1\[0\] _03355_ _03356_ _03357_ vssd1 vssd1
+ vccd1 vccd1 _03358_ sky130_fd_sc_hd__a311o_1
XANTENNA_fanout519_X net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09288_ top.dut.bits_in_buf_next\[1\] top.dut.bits_in_buf_next\[0\] top.dut.bits_in_buf_next\[2\]
+ net297 vssd1 vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__a31o_1
XFILLER_100_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08308_ top.cb_syn.char_path_n\[15\] net195 _04681_ vssd1 vssd1 vccd1 vccd1 _01661_
+ sky130_fd_sc_hd__o21a_1
X_08239_ top.cb_syn.char_path_n\[50\] net375 net336 top.cb_syn.char_path_n\[48\] net180
+ vssd1 vssd1 vccd1 vccd1 _04647_ sky130_fd_sc_hd__a221o_1
XFILLER_60_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_11250_ clknet_leaf_49_clk _01798_ _00605_ vssd1 vssd1 vccd1 vccd1 top.hTree.nullSumIndex\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_106_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11181_ clknet_leaf_20_clk _01729_ _00536_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[83\]
+ sky130_fd_sc_hd__dfrtp_1
X_10201_ net831 net671 vssd1 vssd1 vccd1 vccd1 _00815_ sky130_fd_sc_hd__and2_1
X_10132_ net836 net676 vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__and2_1
XFILLER_0_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10063_ net848 net688 vssd1 vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__and2_1
XANTENNA_input27_A DAT_I[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10965_ clknet_leaf_52_clk _01513_ _00320_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_index\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_55_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10896_ clknet_leaf_40_clk top.header_synthesis.next_header\[1\] _00251_ vssd1 vssd1
+ vccd1 vccd1 top.header_synthesis.header\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_26_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09298__S top.translation.index\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11517_ clknet_leaf_66_clk _02065_ _00872_ vssd1 vssd1 vccd1 vccd1 top.cw1\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__05398__Y _02506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11448_ clknet_leaf_68_clk _01996_ _00803_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.histo_index\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08930__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold209 top.cb_syn.char_path\[44\] vssd1 vssd1 vccd1 vccd1 net1162 sky130_fd_sc_hd__dlygate4sd3_1
X_11379_ clknet_leaf_81_clk _01927_ _00734_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_111_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05940_ top.WB.CPU_DAT_O\[15\] net1337 net306 vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__mux2_1
X_05871_ top.sram_interface.init_counter\[23\] top.sram_interface.init_counter\[22\]
+ _02849_ vssd1 vssd1 vccd1 vccd1 _02850_ sky130_fd_sc_hd__nor3_1
XANTENNA__11365__Q top.findLeastValue.sum\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08590_ top.cb_syn.h_element\[56\] top.cb_syn.h_element\[47\] net533 vssd1 vssd1
+ vccd1 vccd1 _04814_ sky130_fd_sc_hd__mux2_1
X_07610_ top.hTree.state\[2\] top.hTree.state\[5\] net264 vssd1 vssd1 vccd1 vccd1
+ _04193_ sky130_fd_sc_hd__o21a_1
X_07541_ top.cb_syn.pulse_first net536 _02868_ vssd1 vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_66_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08683__A1 _04134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07472_ top.cb_syn.cb_length\[5\] _02518_ _04062_ vssd1 vssd1 vccd1 vccd1 _04063_
+ sky130_fd_sc_hd__a21o_1
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06423_ _03253_ _03250_ net1519 vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__mux2_1
X_09211_ net529 net474 _04528_ _05186_ vssd1 vssd1 vccd1 vccd1 _00010_ sky130_fd_sc_hd__a31o_1
X_09142_ net450 net459 net555 top.sram_interface.word_cnt\[6\] _02774_ vssd1 vssd1
+ vccd1 vccd1 _05152_ sky130_fd_sc_hd__a32o_1
X_06354_ top.hist_data_o\[22\] _03189_ vssd1 vssd1 vccd1 vccd1 _03208_ sky130_fd_sc_hd__nor2_1
XANTENNA__08435__A1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05589__X _02679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05305_ top.compVal\[35\] vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__inv_2
X_09073_ top.cb_syn.pulse_first _02530_ _02869_ vssd1 vssd1 vccd1 vccd1 _05096_ sky130_fd_sc_hd__or3_1
X_06285_ net414 _03011_ _03149_ _02546_ vssd1 vssd1 vccd1 vccd1 _03150_ sky130_fd_sc_hd__a2bb2o_1
Xhold710 top.cb_syn.count\[2\] vssd1 vssd1 vccd1 vccd1 net1663 sky130_fd_sc_hd__dlygate4sd3_1
X_08024_ _04515_ _04520_ _04523_ _04509_ net1677 vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__a32o_1
Xhold721 top.findLeastValue.sum\[39\] vssd1 vssd1 vccd1 vccd1 net1674 sky130_fd_sc_hd__dlygate4sd3_1
Xhold743 top.cb_syn.curr_state\[0\] vssd1 vssd1 vccd1 vccd1 net1696 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_77_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold732 top.findLeastValue.sum\[10\] vssd1 vssd1 vccd1 vccd1 net1685 sky130_fd_sc_hd__dlygate4sd3_1
Xhold754 top.hist_data_o\[6\] vssd1 vssd1 vccd1 vccd1 net1707 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07946__A0 top.findLeastValue.least1\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold765 top.compVal\[10\] vssd1 vssd1 vccd1 vccd1 net1718 sky130_fd_sc_hd__dlygate4sd3_1
Xhold776 top.histogram.total\[4\] vssd1 vssd1 vccd1 vccd1 net1729 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09975_ net803 net643 vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout583_A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10390__B net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08926_ top.WB.CPU_DAT_O\[28\] net1245 net372 vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__mux2_1
XANTENNA__07174__A1 _03817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout750_A net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08857_ net1046 _05039_ _05037_ vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout848_A net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07808_ net441 net1555 net253 top.findLeastValue.sum\[27\] _04352_ vssd1 vssd1 vccd1
+ vccd1 _01832_ sky130_fd_sc_hd__a221o_1
X_08788_ net520 _04952_ _04955_ _04956_ top.translation.index\[4\] vssd1 vssd1 vccd1
+ vccd1 _04971_ sky130_fd_sc_hd__o311a_1
X_07739_ top.findLeastValue.sum\[40\] top.hTree.tree_reg\[40\] net282 vssd1 vssd1
+ vccd1 vccd1 _04297_ sky130_fd_sc_hd__mux2_1
XFILLER_25_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08123__B1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10750_ clknet_leaf_2_clk _01349_ _00169_ vssd1 vssd1 vccd1 vccd1 top.path\[126\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_25_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09409_ net406 _04226_ vssd1 vssd1 vccd1 vccd1 _05283_ sky130_fd_sc_hd__nand2_1
XFILLER_13_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10681_ clknet_leaf_120_clk _01280_ _00100_ vssd1 vssd1 vccd1 vccd1 top.path\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11302_ clknet_leaf_85_clk net1526 _00657_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[45\]
+ sky130_fd_sc_hd__dfrtp_1
X_11233_ clknet_leaf_42_clk _01781_ _00588_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.end_cnt\[6\]
+ sky130_fd_sc_hd__dfstp_1
X_11164_ clknet_leaf_17_clk _01712_ _00519_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[66\]
+ sky130_fd_sc_hd__dfrtp_1
X_11095_ clknet_leaf_30_clk _01643_ _00450_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[125\]
+ sky130_fd_sc_hd__dfrtp_1
X_10115_ net822 net662 vssd1 vssd1 vccd1 vccd1 _00729_ sky130_fd_sc_hd__and2_1
X_10046_ net858 net698 vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__and2_1
Xhold81 top.sram_interface.check vssd1 vssd1 vccd1 vccd1 net1034 sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 top.hTree.tree_reg\[48\] vssd1 vssd1 vccd1 vccd1 net1023 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 top.hTree.node_reg\[41\] vssd1 vssd1 vccd1 vccd1 net1045 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05715__A2 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10948_ clknet_leaf_33_clk _01503_ _00303_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.num_lefts\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08925__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10879_ clknet_leaf_35_clk _00010_ _00234_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.curr_state\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10475__B net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06070_ top.sram_interface.init_counter\[5\] top.sram_interface.init_counter\[4\]
+ _02944_ vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__and3_1
XANTENNA_1 _02725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05651__B2 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_TAPCELL_ROW_113_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07928__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout519 top.cb_syn.char_found vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__buf_2
Xfanout508 top.cb_syn.end_cnt\[2\] vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__clkbuf_4
X_09760_ net773 net613 vssd1 vssd1 vccd1 vccd1 _00374_ sky130_fd_sc_hd__and2_1
X_06972_ _03626_ _03627_ _03628_ _03629_ vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__and4_1
X_09691_ net799 net639 vssd1 vssd1 vccd1 vccd1 _00305_ sky130_fd_sc_hd__and2_1
X_08711_ _02518_ _04902_ vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__nor2_1
X_05923_ _02892_ vssd1 vssd1 vccd1 vccd1 _02893_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_72_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08642_ net210 _04849_ _04851_ _04852_ vssd1 vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__and4_1
XFILLER_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08353__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05706__A2 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05854_ top.compVal\[13\] net169 net155 top.WB.CPU_DAT_O\[13\] vssd1 vssd1 vccd1
+ vccd1 _02288_ sky130_fd_sc_hd__a22o_1
X_05785_ _02804_ vssd1 vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__inv_2
XANTENNA__08105__B1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08573_ net1134 top.cb_syn.char_path_n\[3\] net227 vssd1 vssd1 vccd1 vccd1 _01521_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__11823__Q top.WB.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout164_A net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07524_ top.cb_syn.char_path_n\[104\] top.cb_syn.char_path_n\[103\] top.cb_syn.char_path_n\[102\]
+ top.cb_syn.char_path_n\[101\] net399 net350 vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__mux4_1
X_07455_ top.cb_syn.i\[4\] top.cb_syn.cb_length\[4\] vssd1 vssd1 vccd1 vccd1 _04046_
+ sky130_fd_sc_hd__nand2b_1
XANTENNA__08751__S1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout429_A net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06406_ top.hist_data_o\[2\] top.hist_data_o\[1\] top.hist_data_o\[0\] top.hist_data_o\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03241_ sky130_fd_sc_hd__a31o_1
X_07386_ top.dut.bit_buf\[10\] top.dut.bit_buf\[3\] net721 vssd1 vssd1 vccd1 vccd1
+ _03988_ sky130_fd_sc_hd__mux2_1
XANTENNA__08408__A1 top.cb_syn.char_path_n\[32\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09125_ _02937_ _05110_ _05130_ top.sram_interface.word_cnt\[6\] vssd1 vssd1 vccd1
+ vccd1 _05140_ sky130_fd_sc_hd__o31a_1
X_06337_ top.hist_data_o\[29\] top.hist_data_o\[28\] _03198_ vssd1 vssd1 vccd1 vccd1
+ _03199_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout217_X net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06268_ _03000_ _03133_ _02572_ vssd1 vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__and3b_1
X_09056_ net1252 top.WB.CPU_DAT_O\[1\] net293 vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__mux2_1
X_08007_ top.cb_syn.count\[1\] top.cb_syn.count\[0\] vssd1 vssd1 vccd1 vccd1 _04510_
+ sky130_fd_sc_hd__nand2_1
X_06199_ _02995_ _03067_ vssd1 vssd1 vccd1 vccd1 _03068_ sky130_fd_sc_hd__nor2_1
Xhold562 top.hTree.state\[1\] vssd1 vssd1 vccd1 vccd1 net1515 sky130_fd_sc_hd__dlygate4sd3_1
Xhold540 _03309_ vssd1 vssd1 vccd1 vccd1 net1493 sky130_fd_sc_hd__dlygate4sd3_1
Xhold551 top.histogram.total\[6\] vssd1 vssd1 vccd1 vccd1 net1504 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07919__A0 top.findLeastValue.sum\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold573 _01850_ vssd1 vssd1 vccd1 vccd1 net1526 sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 top.findLeastValue.sum\[45\] vssd1 vssd1 vccd1 vccd1 net1548 sky130_fd_sc_hd__dlygate4sd3_1
Xhold584 top.hTree.tree_reg\[44\] vssd1 vssd1 vccd1 vccd1 net1537 sky130_fd_sc_hd__dlygate4sd3_1
X_09958_ net770 net610 vssd1 vssd1 vccd1 vccd1 _00572_ sky130_fd_sc_hd__and2_1
X_08909_ _04162_ _04187_ _05066_ _05076_ vssd1 vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__a22o_1
XANTENNA__07490__S1 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08344__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09889_ net772 net612 vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__and2_1
XFILLER_18_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ clknet_leaf_116_clk _02367_ _01206_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[29\]
+ sky130_fd_sc_hd__dfrtp_4
X_10802_ clknet_leaf_48_clk _01388_ _00221_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.max_index\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_11782_ clknet_leaf_73_clk _02315_ _01137_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.counter_HTREE\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_56_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08745__S net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10733_ clknet_leaf_119_clk _01332_ _00152_ vssd1 vssd1 vccd1 vccd1 top.path\[109\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08046__A net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_14_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10664_ clknet_leaf_118_clk _01263_ _00083_ vssd1 vssd1 vccd1 vccd1 top.path\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10595_ net841 net681 vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__and2_1
XANTENNA__08480__S net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput60 net60 vssd1 vssd1 vccd1 vccd1 ADR_O[25] sky130_fd_sc_hd__buf_2
X_11216_ clknet_leaf_24_clk _01764_ _00571_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[118\]
+ sky130_fd_sc_hd__dfrtp_2
Xoutput93 net93 vssd1 vssd1 vccd1 vccd1 DAT_O[28] sky130_fd_sc_hd__buf_2
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 ADR_O[9] sky130_fd_sc_hd__buf_2
X_11147_ clknet_leaf_22_clk _01695_ _00502_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[49\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput82 net82 vssd1 vssd1 vccd1 vccd1 DAT_O[18] sky130_fd_sc_hd__buf_2
XANTENNA__07824__S net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08335__B1 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11078_ clknet_leaf_5_clk _01626_ _00433_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[108\]
+ sky130_fd_sc_hd__dfrtp_1
X_10029_ net837 net677 vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__and2_1
XFILLER_56_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06897__B1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05570_ top.cb_syn.char_path\[18\] net557 net312 top.cb_syn.char_path\[114\] vssd1
+ vssd1 vccd1 vccd1 _02663_ sky130_fd_sc_hd__a22o_1
XFILLER_32_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10486__A net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07240_ top.findLeastValue.val1\[33\] top.findLeastValue.val2\[33\] _03833_ _03887_
+ vssd1 vssd1 vccd1 vccd1 _03888_ sky130_fd_sc_hd__o22a_1
XFILLER_118_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07171_ top.findLeastValue.val1\[32\] top.findLeastValue.val2\[32\] vssd1 vssd1 vccd1
+ vccd1 _03829_ sky130_fd_sc_hd__xnor2_1
X_06122_ _02993_ vssd1 vssd1 vccd1 vccd1 _02994_ sky130_fd_sc_hd__inv_2
XANTENNA__08390__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06053_ _02767_ _02835_ _02937_ _02938_ vssd1 vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__or4_1
XANTENNA__09366__A2 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout305 net306 vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__buf_2
XFILLER_99_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout316 _02576_ vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout338 net349 vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__clkbuf_2
X_09812_ net765 net605 vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__and2_1
Xfanout327 net329 vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__clkbuf_2
XFILLER_101_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout349 _04567_ vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__buf_2
XANTENNA__07734__S _04197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06858__B net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09743_ net789 net629 vssd1 vssd1 vccd1 vccd1 _00357_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout281_A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout379_A net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06955_ top.findLeastValue.val2\[6\] net149 net122 _03619_ vssd1 vssd1 vccd1 vccd1
+ _01948_ sky130_fd_sc_hd__o22a_1
X_09674_ net784 net624 vssd1 vssd1 vccd1 vccd1 _00288_ sky130_fd_sc_hd__and2_1
X_05906_ top.CB_read_complete _02879_ _02877_ vssd1 vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__o21a_1
XFILLER_55_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06886_ top.compVal\[40\] top.findLeastValue.val1\[40\] net165 vssd1 vssd1 vccd1
+ vccd1 _03585_ sky130_fd_sc_hd__mux2_1
X_08625_ _04831_ _04835_ _04840_ _04826_ top.cb_syn.num_lefts\[4\] vssd1 vssd1 vccd1
+ vccd1 _01503_ sky130_fd_sc_hd__a32o_1
XFILLER_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05837_ top.compVal\[30\] net169 net155 top.WB.CPU_DAT_O\[30\] vssd1 vssd1 vccd1
+ vccd1 _02305_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout546_A net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_08556_ net1248 top.cb_syn.char_path_n\[20\] net229 vssd1 vssd1 vccd1 vccd1 _01538_
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout167_X net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07507_ top.cb_syn.char_path_n\[84\] top.cb_syn.char_path_n\[83\] top.cb_syn.char_path_n\[82\]
+ top.cb_syn.char_path_n\[81\] net400 net350 vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_53_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05768_ top.translation.index\[4\] net520 net522 net411 vssd1 vssd1 vccd1 vccd1 _02789_
+ sky130_fd_sc_hd__or4_2
X_08487_ net1161 top.cb_syn.char_path_n\[89\] net232 vssd1 vssd1 vccd1 vccd1 _01607_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07689__B _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07837__C1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout334_X net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05699_ net15 net417 net359 top.WB.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 _02359_
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07438_ top.dut.out\[2\] net297 vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__and2_1
X_07369_ top.cw2\[4\] net135 _03547_ net127 _03977_ vssd1 vssd1 vccd1 vccd1 _01892_
+ sky130_fd_sc_hd__a32o_1
XANTENNA__09054__A1 top.WB.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05863__B2 top.WB.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09108_ net479 net469 top.sram_interface.word_cnt\[14\] vssd1 vssd1 vccd1 vccd1 _05127_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__07909__S net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10380_ net854 net694 vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__and2_1
XFILLER_108_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06812__B1 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09039_ net1241 top.WB.CPU_DAT_O\[18\] net291 vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__mux2_1
XANTENNA__09357__A2 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold381 top.path\[32\] vssd1 vssd1 vccd1 vccd1 net1334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold370 top.cb_syn.char_path\[108\] vssd1 vssd1 vccd1 vccd1 net1323 sky130_fd_sc_hd__dlygate4sd3_1
X_11001_ clknet_leaf_34_clk _01549_ _00356_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold392 top.path\[71\] vssd1 vssd1 vccd1 vccd1 net1345 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout850 net857 vssd1 vssd1 vccd1 vccd1 net850 sky130_fd_sc_hd__clkbuf_2
Xfanout861 net877 vssd1 vssd1 vccd1 vccd1 net861 sky130_fd_sc_hd__buf_1
Xfanout872 net876 vssd1 vssd1 vccd1 vccd1 net872 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08317__B1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05551__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08475__S net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11834_ clknet_leaf_100_clk _02350_ _01189_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[12\]
+ sky130_fd_sc_hd__dfrtp_4
X_11765_ clknet_leaf_113_clk _02298_ _01120_ vssd1 vssd1 vccd1 vccd1 top.compVal\[23\]
+ sky130_fd_sc_hd__dfrtp_2
X_11696_ clknet_leaf_62_clk _02229_ _01051_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10716_ clknet_leaf_3_clk _01315_ _00135_ vssd1 vssd1 vccd1 vccd1 top.path\[92\]
+ sky130_fd_sc_hd__dfrtp_1
X_10647_ clknet_leaf_50_clk _00042_ _00066_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.word_cnt\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__05854__B2 top.WB.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09045__A1 top.WB.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05687__X _02761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07819__S net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10578_ net751 net591 vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_11_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06803__B1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07359__B2 top.findLeastValue.sum\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06031__A1 top.WB.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06740_ _02415_ top.findLeastValue.val2\[33\] top.findLeastValue.val2\[32\] _02416_
+ vssd1 vssd1 vccd1 vccd1 _03528_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_108_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06671_ top.findLeastValue.val2\[1\] top.compVal\[1\] vssd1 vssd1 vccd1 vccd1 _03459_
+ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_108_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08410_ top.cb_syn.char_path_n\[30\] net331 _04768_ vssd1 vssd1 vccd1 vccd1 _04769_
+ sky130_fd_sc_hd__a21oi_1
X_05622_ top.hTree.node_reg\[42\] net310 _02705_ _02706_ vssd1 vssd1 vccd1 vccd1 _02707_
+ sky130_fd_sc_hd__a211o_1
X_09390_ top.hTree.nulls\[50\] net405 net244 vssd1 vssd1 vccd1 vccd1 _05271_ sky130_fd_sc_hd__o21a_1
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08341_ top.cb_syn.char_path_n\[93\] net393 _04699_ net512 net438 vssd1 vssd1 vccd1
+ vccd1 _04700_ sky130_fd_sc_hd__a221o_1
X_05553_ _02647_ _02648_ net472 vssd1 vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__o21a_1
XFILLER_51_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05484_ _02541_ _02544_ _02591_ vssd1 vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__or3b_1
X_08272_ top.cb_syn.char_path_n\[33\] net209 _04663_ vssd1 vssd1 vccd1 vccd1 _01679_
+ sky130_fd_sc_hd__o21a_1
XFILLER_20_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07223_ _03839_ _03842_ net271 vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__o21a_1
XANTENNA__05845__B2 top.WB.CPU_DAT_O\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09036__A1 top.WB.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05597__X _02686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07729__S net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08414__A _02505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07154_ _03783_ _03793_ _03811_ vssd1 vssd1 vccd1 vccd1 _03812_ sky130_fd_sc_hd__or3b_1
X_06105_ net561 _02977_ vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__and2_1
X_07085_ top.findLeastValue.val1\[5\] top.findLeastValue.val2\[5\] vssd1 vssd1 vccd1
+ vccd1 _03743_ sky130_fd_sc_hd__or2_1
X_06036_ top.cb_syn.cb_length\[1\] top.cb_syn.cb_length\[0\] vssd1 vssd1 vccd1 vccd1
+ _02927_ sky130_fd_sc_hd__or2_1
Xfanout113 net116 vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__clkbuf_4
Xfanout135 net136 vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06869__A net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout146 net148 vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__buf_2
Xfanout124 net125 vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__buf_2
XANTENNA__06022__A1 top.WB.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input1_A ACK_I vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07987_ _02515_ top.cb_syn.zero_count\[1\] vssd1 vssd1 vccd1 vccd1 _04490_ sky130_fd_sc_hd__nand2_1
XFILLER_87_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout663_A net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout179 net181 vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__buf_2
Xfanout168 net169 vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__clkbuf_4
Xfanout157 _02846_ vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout284_X net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09726_ net738 net578 vssd1 vssd1 vccd1 vccd1 _00340_ sky130_fd_sc_hd__and2_1
X_06938_ top.compVal\[14\] top.findLeastValue.val1\[14\] net162 vssd1 vssd1 vccd1
+ vccd1 _03611_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout451_X net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout549_X net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06869_ net500 _03109_ vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__or2_1
X_09657_ net859 net699 vssd1 vssd1 vccd1 vccd1 _00271_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_38_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08608_ top.cb_syn.num_lefts\[1\] top.cb_syn.num_lefts\[0\] vssd1 vssd1 vccd1 vccd1
+ _04827_ sky130_fd_sc_hd__nand2_1
XANTENNA__05533__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09588_ net846 net686 vssd1 vssd1 vccd1 vccd1 _00202_ sky130_fd_sc_hd__and2_1
X_08539_ net1256 top.cb_syn.char_path_n\[37\] net227 vssd1 vssd1 vccd1 vccd1 _01555_
+ sky130_fd_sc_hd__mux2_1
X_11550_ clknet_leaf_123_clk _02098_ _00905_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10501_ net809 net649 vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__and2_1
XANTENNA__05836__B2 top.WB.CPU_DAT_O\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11481_ clknet_leaf_101_clk _02029_ _00836_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[21\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__09027__A1 top.WB.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10432_ net875 net715 vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__and2_1
X_10363_ net853 net693 vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__and2_1
Xteam_05_930 vssd1 vssd1 vccd1 vccd1 gpio_oeb[10] team_05_930/LO sky130_fd_sc_hd__conb_1
X_10294_ net724 net564 vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__and2_1
Xteam_05_952 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] team_05_952/LO sky130_fd_sc_hd__conb_1
Xteam_05_941 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] team_05_941/LO sky130_fd_sc_hd__conb_1
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06013__A1 top.WB.CPU_DAT_O\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_8_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout691 net697 vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__clkbuf_2
XFILLER_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout680 net681 vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09602__B net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11817_ clknet_leaf_56_clk _02333_ _01172_ vssd1 vssd1 vccd1 vccd1 top.TRN_char_index\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07277__B1 _03864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11748_ clknet_leaf_95_clk _02281_ _01103_ vssd1 vssd1 vccd1 vccd1 top.compVal\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11679_ clknet_leaf_62_clk _02212_ _01034_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_58_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08890_ _05058_ _05059_ vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__nand2_1
X_07910_ top.hTree.tree_reg\[6\] top.findLeastValue.sum\[6\] net247 vssd1 vssd1 vccd1
+ vccd1 _04434_ sky130_fd_sc_hd__mux2_1
XANTENNA__06004__A1 top.WB.CPU_DAT_O\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07841_ net485 _04377_ vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__or2_1
X_07772_ net430 _04322_ _04323_ net263 vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__o211a_1
XANTENNA__07752__A1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09511_ net736 net576 vssd1 vssd1 vccd1 vccd1 _00125_ sky130_fd_sc_hd__and2_1
X_06723_ net494 _02487_ vssd1 vssd1 vccd1 vccd1 _03511_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_69_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05515__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09442_ net847 net687 vssd1 vssd1 vccd1 vccd1 _00056_ sky130_fd_sc_hd__and2_1
X_06654_ net288 _03442_ vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_4_2_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06585_ _02436_ top.findLeastValue.val1\[13\] top.findLeastValue.val1\[12\] _02437_
+ vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__o22a_1
XANTENNA__11831__Q top.WB.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05605_ net1264 net145 _02692_ net177 vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__a22o_1
XANTENNA__05835__A_N net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09373_ net1045 net237 net215 _04294_ vssd1 vssd1 vccd1 vccd1 _01435_ sky130_fd_sc_hd__a22o_1
XANTENNA__05530__A3 _02583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05536_ net458 top.hTree.node_reg\[56\] net361 net422 top.hTree.node_reg\[24\] vssd1
+ vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__a32o_1
X_08324_ top.cb_syn.char_path_n\[7\] net199 _04689_ vssd1 vssd1 vccd1 vccd1 _01653_
+ sky130_fd_sc_hd__o21a_1
XFILLER_20_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_05467_ _02572_ _02574_ net470 vssd1 vssd1 vccd1 vccd1 _02575_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout509_A net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout411_A _02788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08255_ top.cb_syn.char_path_n\[42\] net379 net338 top.cb_syn.char_path_n\[40\] net183
+ vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__a221o_1
XANTENNA__08217__C1 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07206_ net288 _03657_ vssd1 vssd1 vccd1 vccd1 _03864_ sky130_fd_sc_hd__nor2_1
X_05398_ net513 vssd1 vssd1 vccd1 vccd1 _02506_ sky130_fd_sc_hd__inv_2
XANTENNA__05768__A top.translation.index\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08186_ top.cb_syn.char_path_n\[76\] net196 _04620_ vssd1 vssd1 vccd1 vccd1 _01722_
+ sky130_fd_sc_hd__o21a_1
X_07137_ top.findLeastValue.val1\[21\] top.findLeastValue.val2\[21\] vssd1 vssd1 vccd1
+ vccd1 _03795_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout878_A net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout780_A net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07068_ _03716_ _03725_ _03715_ vssd1 vssd1 vccd1 vccd1 _03726_ sky130_fd_sc_hd__or3b_1
XANTENNA__06794__A2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06019_ net1464 top.WB.CPU_DAT_O\[16\] net356 vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__mux2_1
XFILLER_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08940__A0 top.WB.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09709_ net801 net641 vssd1 vssd1 vccd1 vccd1 _00323_ sky130_fd_sc_hd__and2_1
XFILLER_55_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10981_ clknet_leaf_5_clk _01529_ _00336_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05506__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09248__A1 top.cb_syn.char_index\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11602_ clknet_leaf_56_clk _02150_ _00957_ vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11533_ clknet_leaf_1_clk _02081_ _00888_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_96_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08054__A net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11464_ clknet_leaf_94_clk _02012_ _00819_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[4\]
+ sky130_fd_sc_hd__dfstp_1
X_10415_ net859 net699 vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__and2_1
XFILLER_109_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11395_ clknet_leaf_93_clk _01943_ _00750_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_10346_ net871 net711 vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__and2_1
XANTENNA__06785__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10277_ net726 net566 vssd1 vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__and2_1
XFILLER_66_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08931__A0 top.WB.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05745__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_105_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10478__B net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05512__A3 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06370_ net1317 net301 _03218_ vssd1 vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__o21a_1
XANTENNA__08998__A0 top.WB.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05321_ top.compVal\[20\] vssd1 vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__inv_2
XFILLER_119_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08040_ net439 _02861_ _04533_ _04138_ net474 vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__o311ai_4
XANTENNA__07670__A0 top.findLeastValue.least2\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09991_ net847 net687 vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__and2_1
X_08942_ top.WB.CPU_DAT_O\[31\] top.cb_syn.h_element\[63\] net370 vssd1 vssd1 vccd1
+ vccd1 _01368_ sky130_fd_sc_hd__mux2_1
XANTENNA__06776__A2 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07973__A1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11826__Q top.WB.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08873_ _05043_ _05049_ _05050_ vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__nand3b_1
XFILLER_84_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07824_ top.findLeastValue.sum\[23\] top.hTree.tree_reg\[23\] net285 vssd1 vssd1
+ vccd1 vccd1 _04365_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout361_A net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07755_ top.hTree.tree_reg\[37\] top.findLeastValue.sum\[37\] net250 vssd1 vssd1
+ vccd1 vccd1 _04310_ sky130_fd_sc_hd__mux2_1
X_07686_ top.findLeastValue.least2\[4\] top.hTree.tree_reg\[50\] net280 vssd1 vssd1
+ vccd1 vccd1 _04254_ sky130_fd_sc_hd__mux2_1
X_06706_ _02426_ top.findLeastValue.val2\[23\] _02490_ top.compVal\[22\] vssd1 vssd1
+ vccd1 vccd1 _03494_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_37_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09425_ _02809_ _04200_ vssd1 vssd1 vccd1 vccd1 _05293_ sky130_fd_sc_hd__nor2_1
X_06637_ top.compVal\[15\] top.compVal\[14\] top.compVal\[13\] top.compVal\[12\] vssd1
+ vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout626_A net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_09356_ net1004 net242 net218 _04362_ vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__a22o_1
X_06568_ top.compVal\[1\] top.findLeastValue.val1\[1\] vssd1 vssd1 vccd1 vccd1 _03357_
+ sky130_fd_sc_hd__and2b_1
XANTENNA__08989__A0 top.WB.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09287_ net298 _05231_ _04026_ vssd1 vssd1 vccd1 vccd1 top.dut.bit_buf_next\[4\]
+ sky130_fd_sc_hd__o21a_1
X_05519_ top.histogram.sram_out\[27\] net365 _02619_ _02620_ vssd1 vssd1 vccd1 vccd1
+ _02621_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout414_X net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08307_ top.cb_syn.char_path_n\[16\] net374 net333 top.cb_syn.char_path_n\[14\] net179
+ vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__a221o_1
X_06499_ _03283_ _03305_ vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__nor2_1
X_08238_ top.cb_syn.char_path_n\[50\] net198 _04646_ vssd1 vssd1 vccd1 vccd1 _01696_
+ sky130_fd_sc_hd__o21a_1
XFILLER_109_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10200_ net860 net700 vssd1 vssd1 vccd1 vccd1 _00814_ sky130_fd_sc_hd__and2_1
X_08169_ top.cb_syn.char_path_n\[85\] net382 net346 top.cb_syn.char_path_n\[83\] net186
+ vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__a221o_1
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11180_ clknet_leaf_21_clk _01728_ _00535_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[82\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_91_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10131_ net836 net676 vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__and2_1
XANTENNA__08684__A_N _04875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10062_ net863 net703 vssd1 vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__and2_1
XANTENNA__11736__Q top.CB_read_complete vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08748__S net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10964_ clknet_leaf_52_clk _01512_ _00319_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_index\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_10895_ clknet_leaf_40_clk top.header_synthesis.next_header\[0\] _00250_ vssd1 vssd1
+ vccd1 vccd1 top.header_synthesis.header\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_31_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08483__S net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08429__C1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11516_ clknet_leaf_71_clk _02064_ _00871_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least1\[8\]
+ sky130_fd_sc_hd__dfstp_1
X_11447_ clknet_leaf_69_clk _01995_ _00802_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.histo_index\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08827__S0 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11378_ clknet_leaf_81_clk _01926_ _00733_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10329_ net793 net633 vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_111_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05870_ top.sram_interface.init_counter\[21\] top.sram_interface.init_counter\[20\]
+ top.sram_interface.init_counter\[19\] top.sram_interface.init_counter\[18\] vssd1
+ vssd1 vccd1 vccd1 _02849_ sky130_fd_sc_hd__or4_1
XANTENNA__05718__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08380__A1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07540_ _02867_ _02871_ vssd1 vssd1 vccd1 vccd1 _04131_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_80_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07471_ _04046_ _04061_ _04045_ vssd1 vssd1 vccd1 vccd1 _04062_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06221__A2_N _02767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06143__B1 _02767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06422_ top.header_synthesis.count\[6\] top.header_synthesis.count\[5\] _03248_ _03252_
+ vssd1 vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__and4_1
X_09210_ _05184_ _05185_ net530 vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__o21a_1
XANTENNA__08393__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09141_ net479 net541 _02882_ vssd1 vssd1 vccd1 vccd1 _05151_ sky130_fd_sc_hd__and3_1
X_06353_ net1151 _03207_ net302 vssd1 vssd1 vccd1 vccd1 _02138_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_95_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09072_ net539 _04479_ _05095_ _05093_ vssd1 vssd1 vccd1 vccd1 _00006_ sky130_fd_sc_hd__a31o_1
X_05304_ top.compVal\[36\] vssd1 vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__inv_2
X_08023_ top.cb_syn.count\[4\] _04513_ vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__or2_1
X_06284_ net504 _02767_ net503 vssd1 vssd1 vccd1 vccd1 _03149_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08840__C1 top.translation.index\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout207_A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold700 top.sram_interface.TRN_counter\[1\] vssd1 vssd1 vccd1 vccd1 net1653 sky130_fd_sc_hd__dlygate4sd3_1
Xhold711 top.compVal\[0\] vssd1 vssd1 vccd1 vccd1 net1664 sky130_fd_sc_hd__dlygate4sd3_1
Xhold722 top.cb_syn.zeroes\[5\] vssd1 vssd1 vccd1 vccd1 net1675 sky130_fd_sc_hd__dlygate4sd3_1
Xhold733 top.WB.curr_state\[1\] vssd1 vssd1 vccd1 vccd1 net1686 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_77_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold755 top.cb_syn.char_path_n\[85\] vssd1 vssd1 vccd1 vccd1 net1708 sky130_fd_sc_hd__dlygate4sd3_1
Xhold744 top.findLeastValue.sum\[15\] vssd1 vssd1 vccd1 vccd1 net1697 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_103_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold777 top.findLeastValue.sum\[29\] vssd1 vssd1 vccd1 vccd1 net1730 sky130_fd_sc_hd__dlygate4sd3_1
Xhold766 top.compVal\[39\] vssd1 vssd1 vccd1 vccd1 net1719 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_33_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09974_ net797 net637 vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__and2_1
X_08925_ top.WB.CPU_DAT_O\[29\] net1195 net372 vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__mux2_1
XANTENNA__05709__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08856_ _02519_ _05038_ net473 vssd1 vssd1 vccd1 vccd1 _05039_ sky130_fd_sc_hd__a21o_1
X_07807_ net428 _04350_ _04351_ net259 vssd1 vssd1 vccd1 vccd1 _04352_ sky130_fd_sc_hd__o211a_1
X_05999_ _02904_ _02924_ vssd1 vssd1 vccd1 vccd1 _02209_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_48_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout364_X net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout743_A net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08787_ _02521_ _04935_ _04936_ vssd1 vssd1 vccd1 vccd1 _04970_ sky130_fd_sc_hd__and3_1
X_07738_ net444 net1509 net255 top.findLeastValue.sum\[41\] _04296_ vssd1 vssd1 vccd1
+ vccd1 _01846_ sky130_fd_sc_hd__a221o_1
XFILLER_37_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07669_ net257 _04239_ _04240_ top.hTree.tree_reg\[54\] net456 vssd1 vssd1 vccd1
+ vccd1 _01859_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_43_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05488__A2 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09408_ net1002 net242 _05281_ _05282_ vssd1 vssd1 vccd1 vccd1 _01450_ sky130_fd_sc_hd__a22o_1
X_10680_ clknet_leaf_119_clk _01279_ _00099_ vssd1 vssd1 vccd1 vccd1 top.path\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09339_ net983 net236 net215 _04430_ vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_109_Right_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08426__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_106_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08831__C1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11301_ clknet_leaf_104_clk _01849_ _00656_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_107_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_11232_ clknet_leaf_42_clk _01780_ _00587_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.end_cnt\[5\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__05956__A net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05660__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_11163_ clknet_leaf_18_clk _01711_ _00518_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[65\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__05948__A0 top.WB.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10114_ net820 net660 vssd1 vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__and2_1
X_11094_ clknet_leaf_29_clk _01642_ _00449_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[124\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08478__S net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10045_ net839 net679 vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_4_10_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold60 top.hTree.node_reg\[63\] vssd1 vssd1 vccd1 vccd1 net1013 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 top.hTree.node_reg\[21\] vssd1 vssd1 vccd1 vccd1 net1024 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 top.hTree.node_reg\[5\] vssd1 vssd1 vccd1 vccd1 net1035 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_36_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold93 top.translation.writeEn vssd1 vssd1 vccd1 vccd1 net1046 sky130_fd_sc_hd__dlygate4sd3_1
X_10947_ clknet_leaf_33_clk _01502_ _00302_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.num_lefts\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10878_ clknet_leaf_38_clk _00009_ _00233_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_4_14_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_14_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_61_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08822__C1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_2 _03549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07928__A1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07928__B2 top.findLeastValue.sum\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout509 net510 vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__buf_2
XANTENNA__05939__A0 top.WB.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06971_ top.findLeastValue.val2\[2\] top.findLeastValue.val2\[1\] top.findLeastValue.val2\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03629_ sky130_fd_sc_hd__and3_1
XANTENNA__06600__A1 top.compVal\[33\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09690_ net799 net639 vssd1 vssd1 vccd1 vccd1 _00304_ sky130_fd_sc_hd__and2_1
X_08710_ top.cb_syn.i\[4\] _04900_ vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__nand2_1
X_05922_ _02889_ _02891_ vssd1 vssd1 vccd1 vccd1 _02892_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_72_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08641_ top.cb_syn.cb_length\[5\] net389 vssd1 vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__nand2_1
XFILLER_94_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_05853_ top.compVal\[14\] net169 net155 top.WB.CPU_DAT_O\[14\] vssd1 vssd1 vccd1
+ vccd1 _02289_ sky130_fd_sc_hd__a22o_1
XANTENNA__06903__A2 net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05784_ net452 top.sram_interface.counter_HTREE\[3\] top.sram_interface.counter_HTREE\[2\]
+ top.sram_interface.counter_HTREE\[1\] vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__or4b_1
X_08572_ net1126 top.cb_syn.char_path_n\[4\] net227 vssd1 vssd1 vccd1 vccd1 _01522_
+ sky130_fd_sc_hd__mux2_1
X_07523_ top.cb_syn.char_path_n\[100\] top.cb_syn.char_path_n\[99\] top.cb_syn.char_path_n\[98\]
+ top.cb_syn.char_path_n\[97\] net402 net351 vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__mux4_1
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07454_ top.cb_syn.cb_length\[5\] top.cb_syn.i\[5\] vssd1 vssd1 vccd1 vccd1 _04045_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__07864__A0 top.findLeastValue.sum\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06405_ net1115 _03240_ net300 vssd1 vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__mux2_1
X_07385_ net404 vssd1 vssd1 vccd1 vccd1 top.dut.bits_in_buf_next\[0\] sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_20_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout324_A _05087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09124_ _05112_ _05130_ vssd1 vssd1 vccd1 vccd1 _05139_ sky130_fd_sc_hd__or2_1
X_06336_ top.hist_data_o\[27\] top.hist_data_o\[26\] _03197_ vssd1 vssd1 vccd1 vccd1
+ _03198_ sky130_fd_sc_hd__and3_1
X_06267_ top.cw2\[1\] top.cw2\[0\] top.cw2\[2\] vssd1 vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__a21o_1
X_09055_ net1425 top.WB.CPU_DAT_O\[2\] net293 vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout112_X net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08006_ _04507_ _04508_ net538 net476 vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__o211ai_4
XANTENNA__09369__B1 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold530 top.histogram.sram_out\[1\] vssd1 vssd1 vccd1 vccd1 net1483 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05642__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout693_A net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06198_ top.cw1\[4\] _02993_ top.cw1\[5\] vssd1 vssd1 vccd1 vccd1 _03067_ sky130_fd_sc_hd__a21oi_1
Xhold552 top.cb_syn.curr_path\[127\] vssd1 vssd1 vccd1 vccd1 net1505 sky130_fd_sc_hd__dlygate4sd3_1
Xhold563 top.histogram.total\[28\] vssd1 vssd1 vccd1 vccd1 net1516 sky130_fd_sc_hd__dlygate4sd3_1
Xhold541 top.histogram.total\[20\] vssd1 vssd1 vccd1 vccd1 net1494 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold596 top.cb_syn.curr_index\[5\] vssd1 vssd1 vccd1 vccd1 net1549 sky130_fd_sc_hd__dlygate4sd3_1
Xhold585 top.cb_syn.cb_length\[3\] vssd1 vssd1 vccd1 vccd1 net1538 sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 top.sram_interface.write_counter_FLV\[2\] vssd1 vssd1 vccd1 vccd1 net1527
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout481_X net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout860_A net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09957_ net770 net610 vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__and2_1
X_08908_ top.cb_syn.max_index\[5\] _05065_ _04188_ vssd1 vssd1 vccd1 vccd1 _05076_
+ sky130_fd_sc_hd__o21a_1
XFILLER_66_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09888_ net773 net613 vssd1 vssd1 vccd1 vccd1 _00502_ sky130_fd_sc_hd__and2_1
X_08839_ _04987_ _04988_ net520 _04985_ vssd1 vssd1 vccd1 vccd1 _05022_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_28_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ clknet_leaf_116_clk _02366_ _01205_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[28\]
+ sky130_fd_sc_hd__dfrtp_4
X_10801_ clknet_leaf_48_clk _01387_ _00220_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.max_index\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_11781_ clknet_leaf_67_clk _02314_ _01136_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.counter_HTREE\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_56_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07930__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07855__A0 top.findLeastValue.sum\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10732_ clknet_leaf_118_clk _01331_ _00151_ vssd1 vssd1 vccd1 vccd1 top.path\[108\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10663_ clknet_leaf_114_clk _01262_ _00082_ vssd1 vssd1 vccd1 vccd1 top.path\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10594_ net747 net587 vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__and2_1
XANTENNA__05686__A net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput50 net50 vssd1 vssd1 vccd1 vccd1 ADR_O[15] sky130_fd_sc_hd__buf_2
Xoutput61 net61 vssd1 vssd1 vccd1 vccd1 ADR_O[26] sky130_fd_sc_hd__buf_2
X_11215_ clknet_leaf_23_clk _01763_ _00570_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[117\]
+ sky130_fd_sc_hd__dfrtp_2
Xoutput72 net454 vssd1 vssd1 vccd1 vccd1 CYC_O sky130_fd_sc_hd__buf_2
Xoutput94 net94 vssd1 vssd1 vccd1 vccd1 DAT_O[29] sky130_fd_sc_hd__buf_2
XFILLER_110_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__08583__A1 top.cb_syn.char_index\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput83 net83 vssd1 vssd1 vccd1 vccd1 DAT_O[19] sky130_fd_sc_hd__buf_2
X_11146_ clknet_leaf_21_clk _01694_ _00501_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_8_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11077_ clknet_leaf_5_clk _01625_ _00432_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[107\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08335__A1 top.cb_syn.char_path_n\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10028_ net823 net663 vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__and2_1
XFILLER_63_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08099__B1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07840__S net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06309__X _03172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10486__B net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07170_ _03824_ _03827_ vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__nand2_1
X_06121_ top.cw1\[2\] top.cw1\[1\] top.cw1\[0\] top.cw1\[3\] vssd1 vssd1 vccd1 vccd1
+ _02993_ sky130_fd_sc_hd__a31o_1
X_06052_ top.sram_interface.word_cnt\[1\] top.sram_interface.word_cnt\[12\] vssd1
+ vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_120_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_120_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__05624__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08574__A1 top.cb_syn.char_path_n\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout339 net341 vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__buf_2
X_09811_ net765 net605 vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__and2_1
Xfanout306 net307 vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__clkbuf_4
Xfanout328 net329 vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__clkbuf_4
Xfanout317 net318 vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__clkbuf_4
X_09742_ net783 net623 vssd1 vssd1 vccd1 vccd1 _00356_ sky130_fd_sc_hd__and2_1
XFILLER_86_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload11_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06954_ top.compVal\[6\] top.findLeastValue.val1\[6\] net164 vssd1 vssd1 vccd1 vccd1
+ _03619_ sky130_fd_sc_hd__mux2_1
X_09673_ net784 net624 vssd1 vssd1 vccd1 vccd1 _00287_ sky130_fd_sc_hd__and2_1
XANTENNA__06220__A net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05905_ _02451_ top.sram_interface.CB_write_counter\[0\] _02857_ top.sram_interface.CB_read_counter
+ vssd1 vssd1 vccd1 vccd1 _02879_ sky130_fd_sc_hd__o211a_1
XANTENNA__11834__Q top.WB.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout274_A _03658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06885_ top.findLeastValue.val2\[41\] net149 net123 _03584_ vssd1 vssd1 vccd1 vccd1
+ _01983_ sky130_fd_sc_hd__o22a_1
X_08624_ top.cb_syn.num_lefts\[4\] _04829_ vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__or2_1
X_05836_ top.compVal\[31\] net169 net155 top.WB.CPU_DAT_O\[31\] vssd1 vssd1 vccd1
+ vccd1 _02306_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_85_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07603__X _04187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08555_ net1217 top.cb_syn.char_path_n\[21\] net229 vssd1 vssd1 vccd1 vccd1 _01539_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07750__S net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09531__A net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05767_ net523 net524 vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__or2_2
X_07506_ _04085_ _04096_ _04067_ vssd1 vssd1 vccd1 vccd1 _04097_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout441_A net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08486_ net1135 top.cb_syn.char_path_n\[90\] net232 vssd1 vssd1 vccd1 vccd1 _01608_
+ sky130_fd_sc_hd__mux2_1
X_05698_ net16 net415 net309 top.WB.CPU_DAT_O\[22\] vssd1 vssd1 vccd1 vccd1 _02360_
+ sky130_fd_sc_hd__o22a_1
X_07437_ _03994_ _04001_ _04032_ _03999_ _04029_ vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout706_A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07368_ top.cw1\[4\] net167 _03553_ net501 vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__a22o_1
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09107_ _02529_ _02812_ _05125_ vssd1 vssd1 vccd1 vccd1 _05126_ sky130_fd_sc_hd__or3_1
X_06319_ top.hist_data_o\[12\] _03178_ _03181_ vssd1 vssd1 vccd1 vccd1 _03182_ sky130_fd_sc_hd__and3_1
XANTENNA__08801__A2 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07299_ net269 _03931_ _03932_ net274 top.findLeastValue.sum\[21\] vssd1 vssd1 vccd1
+ vccd1 _01917_ sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_111_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_111_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout696_X net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09038_ net1093 top.WB.CPU_DAT_O\[19\] net291 vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__mux2_1
XANTENNA__10913__Q top.header_synthesis.bit1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold371 net71 vssd1 vssd1 vccd1 vccd1 net1324 sky130_fd_sc_hd__dlygate4sd3_1
Xhold360 top.cb_syn.char_path\[109\] vssd1 vssd1 vccd1 vccd1 net1313 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07368__A2 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11000_ clknet_leaf_28_clk _01548_ _00355_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[30\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold382 top.cb_syn.char_path\[111\] vssd1 vssd1 vccd1 vccd1 net1335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 top.path\[120\] vssd1 vssd1 vccd1 vccd1 net1346 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07925__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout851 net857 vssd1 vssd1 vccd1 vccd1 net851 sky130_fd_sc_hd__clkbuf_2
Xfanout840 net841 vssd1 vssd1 vccd1 vccd1 net840 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout873 net876 vssd1 vssd1 vccd1 vccd1 net873 sky130_fd_sc_hd__clkbuf_2
Xfanout862 net863 vssd1 vssd1 vccd1 vccd1 net862 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11971__A net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11833_ clknet_leaf_99_clk _02349_ _01188_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07828__B1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11764_ clknet_leaf_101_clk _02297_ _01119_ vssd1 vssd1 vccd1 vccd1 top.compVal\[22\]
+ sky130_fd_sc_hd__dfrtp_2
X_11695_ clknet_leaf_61_clk _02228_ _01050_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10715_ clknet_leaf_3_clk _01314_ _00134_ vssd1 vssd1 vccd1 vccd1 top.path\[91\]
+ sky130_fd_sc_hd__dfrtp_1
X_10646_ clknet_leaf_49_clk _00041_ _00065_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.word_cnt\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08491__S net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05854__A2 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10577_ net810 net650 vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_11_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_102_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_102_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05606__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__07835__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11129_ clknet_leaf_28_clk _01677_ _00484_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[31\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_1_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_06670_ _02438_ top.findLeastValue.val2\[11\] top.findLeastValue.val2\[10\] _02439_
+ vssd1 vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_108_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07570__S _04144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05621_ top.histogram.sram_out\[10\] net363 net419 top.hTree.node_reg\[10\] vssd1
+ vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__a22o_1
X_08340_ top.cb_syn.char_path_n\[95\] top.cb_syn.char_path_n\[96\] net516 vssd1 vssd1
+ vccd1 vccd1 _04699_ sky130_fd_sc_hd__mux2_1
X_05552_ top.cb_syn.char_path\[21\] net559 net314 top.cb_syn.char_path\[117\] vssd1
+ vssd1 vccd1 vccd1 _02648_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_50_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05483_ net212 _02590_ top.WB.curr_state\[0\] vssd1 vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__or3b_1
X_08271_ top.cb_syn.char_path_n\[34\] net388 net347 top.cb_syn.char_path_n\[32\] net192
+ vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__a221o_1
XANTENNA__07295__B2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07222_ _03839_ _03842_ vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__nand2_1
XANTENNA__05845__A2 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07153_ top.findLeastValue.val1\[16\] top.findLeastValue.val2\[16\] _03784_ vssd1
+ vssd1 vccd1 vccd1 _03811_ sky130_fd_sc_hd__a21o_1
XFILLER_20_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__06914__S net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06104_ top.TRN_char_index\[5\] top.TRN_char_index\[4\] _02975_ vssd1 vssd1 vccd1
+ vccd1 _02977_ sky130_fd_sc_hd__and3_1
XFILLER_105_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11829__Q top.WB.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07084_ top.findLeastValue.val1\[5\] top.findLeastValue.val2\[5\] vssd1 vssd1 vccd1
+ vccd1 _03742_ sky130_fd_sc_hd__and2_1
X_06035_ top.hist_data_o\[0\] top.WB.CPU_DAT_O\[0\] net355 vssd1 vssd1 vccd1 vccd1
+ _02175_ sky130_fd_sc_hd__mux2_1
XANTENNA__07745__S net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout136 _03443_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__buf_2
XANTENNA_fanout391_A net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout125 _03550_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__clkbuf_4
Xfanout114 net115 vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__clkbuf_4
Xfanout147 net148 vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__clkbuf_2
X_07986_ _02509_ top.cb_syn.zero_count\[7\] vssd1 vssd1 vccd1 vccd1 _04489_ sky130_fd_sc_hd__and2_1
XANTENNA__05773__B top.findLeastValue.least1\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout158 _02783_ vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__buf_2
Xfanout169 _02845_ vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__clkbuf_4
XFILLER_74_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09725_ net735 net575 vssd1 vssd1 vccd1 vccd1 _00339_ sky130_fd_sc_hd__and2_1
X_06937_ top.findLeastValue.val2\[15\] net146 net120 _03610_ vssd1 vssd1 vccd1 vccd1
+ _01957_ sky130_fd_sc_hd__o22a_1
X_09656_ net784 net624 vssd1 vssd1 vccd1 vccd1 _00270_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout277_X net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08607_ _04556_ _04561_ _04825_ vssd1 vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__or3b_4
X_06868_ net498 _03570_ _03578_ vssd1 vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_38_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05819_ net478 top.sram_interface.word_cnt\[9\] net960 vssd1 vssd1 vccd1 vccd1 _02311_
+ sky130_fd_sc_hd__a21o_1
X_09587_ net843 net683 vssd1 vssd1 vccd1 vccd1 _00201_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout823_A net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout444_X net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06799_ top.findLeastValue.val1\[31\] net132 net116 net1641 vssd1 vssd1 vccd1 vccd1
+ _02039_ sky130_fd_sc_hd__o22a_1
X_08538_ net1069 top.cb_syn.char_path_n\[38\] net226 vssd1 vssd1 vccd1 vccd1 _01556_
+ sky130_fd_sc_hd__mux2_1
X_08469_ net1426 top.cb_syn.char_path_n\[107\] net220 vssd1 vssd1 vccd1 vccd1 _01625_
+ sky130_fd_sc_hd__mux2_1
X_10500_ net808 net648 vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__and2_1
XANTENNA__05836__A2 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11480_ clknet_leaf_101_clk _02028_ _00835_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[20\]
+ sky130_fd_sc_hd__dfstp_2
X_10431_ net875 net715 vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__and2_1
XFILLER_10_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10362_ net871 net711 vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__and2_1
X_10293_ net724 net564 vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__and2_1
XANTENNA__06797__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xteam_05_942 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] team_05_942/LO sky130_fd_sc_hd__conb_1
Xteam_05_931 vssd1 vssd1 vccd1 vccd1 gpio_oeb[11] team_05_931/LO sky130_fd_sc_hd__conb_1
Xteam_05_953 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] team_05_953/LO sky130_fd_sc_hd__conb_1
Xhold190 top.cb_syn.char_path\[12\] vssd1 vssd1 vccd1 vccd1 net1143 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout692 net693 vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__clkbuf_2
Xfanout681 net682 vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__buf_1
Xfanout670 net671 vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08171__C1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11816_ clknet_leaf_56_clk _02332_ _01171_ vssd1 vssd1 vccd1 vccd1 top.TRN_char_index\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_11747_ clknet_leaf_94_clk _02280_ _01102_ vssd1 vssd1 vccd1 vccd1 top.compVal\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11678_ clknet_leaf_61_clk _02211_ _01033_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10629_ net798 net638 vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06788__B1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07840_ top.hTree.tree_reg\[20\] top.findLeastValue.sum\[20\] net249 vssd1 vssd1
+ vccd1 vccd1 _04378_ sky130_fd_sc_hd__mux2_1
X_07771_ net490 _04321_ vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__or2_1
XANTENNA__07752__A2 _04306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09510_ net725 net565 vssd1 vssd1 vccd1 vccd1 _00124_ sky130_fd_sc_hd__and2_1
X_06722_ top.compVal\[25\] _02488_ vssd1 vssd1 vccd1 vccd1 _03510_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09441_ net860 net700 vssd1 vssd1 vccd1 vccd1 _00055_ sky130_fd_sc_hd__and2_1
X_06653_ _03424_ _03441_ vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_35_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09372_ net1058 net238 net215 _04298_ vssd1 vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__a22o_1
X_06584_ _02435_ top.findLeastValue.val1\[14\] top.findLeastValue.val1\[13\] _02436_
+ _03372_ vssd1 vssd1 vccd1 vccd1 _03373_ sky130_fd_sc_hd__a221o_1
X_05604_ top.histogram.sram_out\[13\] net363 net421 top.hTree.node_reg\[13\] _02691_
+ vssd1 vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__a221o_1
X_05535_ _02632_ _02633_ net476 vssd1 vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__o21a_1
X_08323_ top.cb_syn.char_path_n\[8\] net378 net337 top.cb_syn.char_path_n\[6\] net182
+ vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__a221o_1
XFILLER_20_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_fanout237_A net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05466_ _02536_ _02573_ vssd1 vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_08254_ top.cb_syn.char_path_n\[42\] net195 _04654_ vssd1 vssd1 vccd1 vccd1 _01688_
+ sky130_fd_sc_hd__o21a_1
X_05397_ net508 vssd1 vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__inv_2
XANTENNA__05768__B net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08185_ top.cb_syn.char_path_n\[77\] net374 net334 top.cb_syn.char_path_n\[75\] net179
+ vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__a221o_1
X_07205_ _03659_ _03860_ _03861_ vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__nand3_1
XFILLER_4_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07136_ top.findLeastValue.val1\[20\] top.findLeastValue.val2\[20\] vssd1 vssd1 vccd1
+ vccd1 _03794_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06779__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07067_ _03717_ _03719_ vssd1 vssd1 vccd1 vccd1 _03725_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_18_Left_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05784__A net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06018_ net1625 top.WB.CPU_DAT_O\[17\] net357 vssd1 vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__mux2_1
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout394_X net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09708_ net801 net641 vssd1 vssd1 vccd1 vccd1 _00322_ sky130_fd_sc_hd__and2_1
X_07969_ top.findLeastValue.alternator_timer\[1\] top.findLeastValue.alternator_timer\[0\]
+ _04473_ vssd1 vssd1 vccd1 vccd1 _04476_ sky130_fd_sc_hd__a21boi_1
XANTENNA__06951__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05754__B2 top.WB.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08153__C1 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_27_Left_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10980_ clknet_leaf_10_clk _01528_ _00335_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_09639_ net804 net644 vssd1 vssd1 vccd1 vccd1 _00253_ sky130_fd_sc_hd__and2_1
XFILLER_28_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11601_ clknet_leaf_63_clk _02149_ _00956_ vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05959__A net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11532_ clknet_leaf_5_clk _02080_ _00887_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_99_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06781__C _03545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11463_ clknet_leaf_94_clk _02011_ _00818_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[3\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_7_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10414_ net794 net634 vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__and2_1
XANTENNA__05690__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_36_Left_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11394_ clknet_leaf_92_clk _01942_ _00749_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_10345_ net854 net694 vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10276_ net726 net566 vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_45_Left_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05320_ top.compVal\[21\] vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_54_Left_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05681__B1 _02755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09990_ net846 net686 vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__and2_1
X_08941_ net479 top.sram_interface.word_cnt\[2\] vssd1 vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__nand2_2
XANTENNA__07973__A2 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09175__A1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08872_ top.translation.index\[3\] _05048_ vssd1 vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__nand2_1
XFILLER_84_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_63_Left_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07823_ net442 net1465 net256 top.findLeastValue.sum\[24\] _04364_ vssd1 vssd1 vccd1
+ vccd1 _01829_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout187_A net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07754_ top.findLeastValue.sum\[37\] top.hTree.tree_reg\[37\] net284 vssd1 vssd1
+ vccd1 vccd1 _04309_ sky130_fd_sc_hd__mux2_1
XFILLER_65_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07685_ net263 _04252_ _04253_ net1021 net446 vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_48_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11842__Q top.WB.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06705_ _03491_ _03492_ vssd1 vssd1 vccd1 vccd1 _03493_ sky130_fd_sc_hd__or2_1
X_09424_ net967 _05292_ net245 vssd1 vssd1 vccd1 vccd1 _01456_ sky130_fd_sc_hd__mux2_1
X_06636_ top.compVal\[11\] top.compVal\[10\] top.compVal\[9\] top.compVal\[8\] vssd1
+ vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__or4_1
Xclkbuf_leaf_91_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_91_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout619_A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09355_ net1014 net241 net216 _04366_ vssd1 vssd1 vccd1 vccd1 _01417_ sky130_fd_sc_hd__a22o_1
XANTENNA__08438__B1 top.cb_syn.end_cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06567_ top.compVal\[2\] top.findLeastValue.val1\[2\] vssd1 vssd1 vccd1 vccd1 _03356_
+ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout521_A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09286_ _03996_ _04038_ vssd1 vssd1 vccd1 vccd1 _05231_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_72_Left_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05518_ net457 top.hTree.node_reg\[59\] net362 _02599_ top.hTree.node_reg\[27\] vssd1
+ vssd1 vccd1 vccd1 _02620_ sky130_fd_sc_hd__a32o_1
X_08306_ top.cb_syn.char_path_n\[16\] net197 _04680_ vssd1 vssd1 vccd1 vccd1 _01662_
+ sky130_fd_sc_hd__o21a_1
X_06498_ net1672 _03282_ vssd1 vssd1 vccd1 vccd1 _03305_ sky130_fd_sc_hd__nor2_1
X_05449_ net549 _02555_ top.sram_interface.word_cnt\[9\] vssd1 vssd1 vccd1 vccd1 _02557_
+ sky130_fd_sc_hd__a21o_1
X_08237_ top.cb_syn.char_path_n\[51\] net376 net335 top.cb_syn.char_path_n\[49\] net181
+ vssd1 vssd1 vccd1 vccd1 _04646_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_7_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05672__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout407_X net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_08168_ net1708 net208 _04611_ vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__o21a_1
X_08099_ top.cb_syn.char_path_n\[120\] net383 net342 top.cb_syn.char_path_n\[118\]
+ net187 vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__a221o_1
X_07119_ top.findLeastValue.val1\[8\] top.findLeastValue.val2\[8\] _03734_ _03732_
+ vssd1 vssd1 vccd1 vccd1 _03777_ sky130_fd_sc_hd__a31o_1
XANTENNA__06767__A3 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10130_ net836 net676 vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__and2_1
XANTENNA__09166__A1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout776_X net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10061_ net846 net686 vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__and2_1
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10963_ clknet_leaf_52_clk _01511_ _00318_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_index\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_16_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_82_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_clk sky130_fd_sc_hd__clkbuf_8
X_10894_ clknet_leaf_38_clk top.header_synthesis.next_start _00249_ vssd1 vssd1 vccd1
+ vccd1 top.header_synthesis.start sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_26_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11515_ clknet_leaf_69_clk _02063_ _00870_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least1\[7\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_8_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__05663__B1 _02740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11446_ clknet_leaf_69_clk _01994_ _00801_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.histo_index\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11199__Q top.cb_syn.char_path_n\[101\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11377_ clknet_leaf_80_clk _01925_ _00732_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10328_ net792 net632 vssd1 vssd1 vccd1 vccd1 _00942_ sky130_fd_sc_hd__and2_1
XFILLER_59_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10259_ net865 net705 vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__and2_1
XFILLER_94_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05718__B2 top.WB.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06915__B1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xclkbuf_leaf_73_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_66_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07470_ _04050_ _04059_ _04051_ _04048_ vssd1 vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_45_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06421_ top.header_synthesis.write_num_lefts _03251_ vssd1 vssd1 vccd1 vccd1 _03252_
+ sky130_fd_sc_hd__nor2_1
X_09140_ _05150_ _05148_ _05086_ vssd1 vssd1 vccd1 vccd1 _00052_ sky130_fd_sc_hd__or3b_1
X_06352_ top.hist_data_o\[23\] _03190_ _03196_ vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__o21ba_1
X_06283_ net1040 net141 _03148_ vssd1 vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__a21o_1
X_09071_ _02859_ _02860_ _02867_ _05094_ vssd1 vssd1 vccd1 vccd1 _05095_ sky130_fd_sc_hd__nor4_1
X_05303_ top.compVal\[38\] vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__inv_2
X_08022_ _04517_ _04520_ _04522_ _04509_ net1671 vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__a32o_1
XANTENNA__05654__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold701 top.header_synthesis.write_char_path vssd1 vssd1 vccd1 vccd1 net1654 sky130_fd_sc_hd__dlygate4sd3_1
Xhold712 top.hist_addr\[6\] vssd1 vssd1 vccd1 vccd1 net1665 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06922__S net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold723 top.header_synthesis.count\[3\] vssd1 vssd1 vccd1 vccd1 net1676 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_77_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold745 top.hTree.state\[2\] vssd1 vssd1 vccd1 vccd1 net1698 sky130_fd_sc_hd__dlygate4sd3_1
Xhold734 top.findLeastValue.sum\[7\] vssd1 vssd1 vccd1 vccd1 net1687 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold756 top.controller.fin_reg\[6\] vssd1 vssd1 vccd1 vccd1 net1709 sky130_fd_sc_hd__dlygate4sd3_1
X_09973_ net790 net630 vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__and2_1
Xhold767 top.hist_data_o\[15\] vssd1 vssd1 vccd1 vccd1 net1720 sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 top.compVal\[0\] vssd1 vssd1 vccd1 vccd1 net1731 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_89_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09148__A1 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08924_ top.WB.CPU_DAT_O\[30\] net1073 net372 vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__mux2_1
XANTENNA__11837__Q top.WB.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08356__C1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05709__B2 top.WB.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08855_ _02790_ net325 top.translation.totalEn vssd1 vssd1 vccd1 vccd1 _05038_ sky130_fd_sc_hd__o21bai_1
X_07806_ net486 _04349_ vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08786_ net436 _04965_ _04968_ vssd1 vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__or3_1
X_05998_ top.sram_interface.init_counter\[1\] _02903_ vssd1 vssd1 vccd1 vccd1 _02924_
+ sky130_fd_sc_hd__nor2_1
X_07737_ net429 _04294_ _04295_ net260 vssd1 vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_64_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout357_X net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08123__A2 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07668_ _02495_ net286 net485 vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__a21oi_1
X_07599_ net531 _02525_ top.cb_syn.h_element\[55\] net539 vssd1 vssd1 vccd1 vccd1
+ _04184_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_80_Left_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09407_ top.hTree.nulls\[56\] net407 net245 vssd1 vssd1 vccd1 vccd1 _05282_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout524_X net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06619_ top.compVal\[33\] _02468_ _03402_ vssd1 vssd1 vccd1 vccd1 _03408_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_23_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09338_ net1003 net238 net215 _04434_ vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__a22o_1
X_09269_ top.cb_syn.zero_count\[4\] _05219_ vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__nand2_1
X_11300_ clknet_leaf_104_clk _01848_ _00655_ vssd1 vssd1 vccd1 vccd1 top.hTree.tree_reg\[43\]
+ sky130_fd_sc_hd__dfrtp_1
X_11231_ clknet_leaf_19_clk _01779_ _00586_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.end_cnt\[4\]
+ sky130_fd_sc_hd__dfstp_2
X_11162_ clknet_leaf_18_clk _01710_ _00517_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[64\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07493__S0 _04072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10113_ net823 net663 vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__and2_1
X_11093_ clknet_leaf_29_clk _01641_ _00448_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[123\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_76_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08898__B1 _04187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10044_ net845 net685 vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__and2_1
XANTENNA_input32_A DAT_I[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold50 top.hTree.node_reg\[6\] vssd1 vssd1 vccd1 vccd1 net1003 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 top.histogram.init_edge vssd1 vssd1 vccd1 vccd1 net1036 sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 top.hTree.node_reg\[23\] vssd1 vssd1 vccd1 vccd1 net1014 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 top.hTree.node_reg\[17\] vssd1 vssd1 vccd1 vccd1 net1025 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 top.histogram.out_of_init vssd1 vssd1 vccd1 vccd1 net1047 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_55_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_clk sky130_fd_sc_hd__clkbuf_8
X_10946_ clknet_leaf_33_clk _01501_ _00301_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.num_lefts\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10877_ clknet_leaf_41_clk _00008_ _00232_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.curr_state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07873__A1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06308__A net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__05636__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_3 _04466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11429_ clknet_leaf_87_clk _01977_ _00784_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[35\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_6_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08050__A1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06061__B1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07484__S0 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06970_ top.findLeastValue.val2\[6\] top.findLeastValue.val2\[5\] top.findLeastValue.val2\[4\]
+ top.findLeastValue.val2\[3\] vssd1 vssd1 vccd1 vccd1 _03628_ sky130_fd_sc_hd__and4_1
XANTENNA__05882__A net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05921_ top.sram_interface.TRN_counter\[0\] _02890_ vssd1 vssd1 vccd1 vccd1 _02891_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_72_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08889__B1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09073__B _02530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08640_ top.cb_syn.cb_length\[5\] net389 vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__or2_1
XANTENNA__08353__A2 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05852_ top.compVal\[15\] net168 net154 top.WB.CPU_DAT_O\[15\] vssd1 vssd1 vccd1
+ vccd1 _02290_ sky130_fd_sc_hd__a22o_1
XANTENNA_wire325_X net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05783_ _02802_ net451 net458 vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__and3b_1
Xclkbuf_leaf_46_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_clk sky130_fd_sc_hd__clkbuf_8
X_08571_ net1086 top.cb_syn.char_path_n\[5\] net226 vssd1 vssd1 vccd1 vccd1 _01523_
+ sky130_fd_sc_hd__mux2_1
X_07522_ _04109_ _04110_ _04111_ _04112_ _04072_ _04071_ vssd1 vssd1 vccd1 vccd1 _04113_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07313__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09302__B2 _02523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_07453_ top.cb_syn.cb_length\[6\] top.cb_syn.i\[6\] vssd1 vssd1 vccd1 vccd1 _04044_
+ sky130_fd_sc_hd__xor2_1
X_06404_ _03175_ _03239_ vssd1 vssd1 vccd1 vccd1 _03240_ sky130_fd_sc_hd__nor2_1
X_07384_ net722 top.dut.bits_in_buf\[0\] vssd1 vssd1 vccd1 vccd1 _03987_ sky130_fd_sc_hd__xnor2_2
X_09123_ net550 _05136_ _05138_ _02578_ vssd1 vssd1 vccd1 vccd1 _00048_ sky130_fd_sc_hd__a211o_1
XFILLER_50_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06335_ top.hist_data_o\[25\] top.hist_data_o\[24\] _03196_ vssd1 vssd1 vccd1 vccd1
+ _03197_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_20_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06266_ net503 _03131_ net412 vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__mux2_1
X_09054_ net1212 top.WB.CPU_DAT_O\[3\] net293 vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__mux2_1
X_08005_ top.cb_syn.h_element\[63\] _04125_ vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__nand2_1
Xhold520 _00035_ vssd1 vssd1 vccd1 vccd1 net1473 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09369__B2 _04310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold542 top.header_synthesis.count\[4\] vssd1 vssd1 vccd1 vccd1 net1495 sky130_fd_sc_hd__dlygate4sd3_1
Xhold553 top.sram_interface.init_counter\[10\] vssd1 vssd1 vccd1 vccd1 net1506 sky130_fd_sc_hd__dlygate4sd3_1
X_06197_ top.cw2\[4\] _03001_ top.cw2\[5\] vssd1 vssd1 vccd1 vccd1 _03066_ sky130_fd_sc_hd__a21o_1
Xhold531 top.hTree.nullSumIndex\[1\] vssd1 vssd1 vccd1 vccd1 net1484 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout686_A net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold575 top.hTree.nulls\[54\] vssd1 vssd1 vccd1 vccd1 net1528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 top.hTree.node_reg\[29\] vssd1 vssd1 vccd1 vccd1 net1517 sky130_fd_sc_hd__dlygate4sd3_1
Xhold586 top.hTree.tree_reg\[25\] vssd1 vssd1 vccd1 vccd1 net1539 sky130_fd_sc_hd__dlygate4sd3_1
Xhold597 top.histogram.total\[3\] vssd1 vssd1 vccd1 vccd1 net1550 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11567__Q top.histogram.sram_out\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09956_ net769 net609 vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__and2_1
X_08907_ top.cb_syn.max_index\[6\] _05072_ _05075_ vssd1 vssd1 vccd1 vccd1 _01392_
+ sky130_fd_sc_hd__o21ba_1
X_09887_ net772 net612 vssd1 vssd1 vccd1 vccd1 _00501_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout853_A net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08344__A2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08838_ net520 _05003_ _05006_ _05009_ _05020_ vssd1 vssd1 vccd1 vccd1 _05021_ sky130_fd_sc_hd__o32a_1
Xclkbuf_leaf_37_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08769_ net433 _04950_ _04951_ vssd1 vssd1 vccd1 vccd1 _04952_ sky130_fd_sc_hd__o21a_1
X_10800_ clknet_leaf_39_clk _00002_ _00219_ vssd1 vssd1 vccd1 vccd1 top.WB.curr_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11780_ clknet_leaf_66_clk _02313_ _01135_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.counter_HTREE\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10731_ clknet_leaf_111_clk _01330_ _00150_ vssd1 vssd1 vccd1 vccd1 top.path\[107\]
+ sky130_fd_sc_hd__dfrtp_1
X_10662_ clknet_leaf_114_clk _01261_ _00081_ vssd1 vssd1 vccd1 vccd1 top.path\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11969__A net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10593_ net788 net628 vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__and2_1
XANTENNA__05618__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08062__B net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11214_ clknet_leaf_23_clk _01762_ _00569_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[116\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput51 net51 vssd1 vssd1 vccd1 vccd1 ADR_O[16] sky130_fd_sc_hd__buf_2
Xoutput62 net62 vssd1 vssd1 vccd1 vccd1 ADR_O[28] sky130_fd_sc_hd__buf_2
X_11145_ clknet_leaf_7_clk _01693_ _00500_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[47\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 DAT_O[0] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_8_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 DAT_O[1] sky130_fd_sc_hd__buf_2
XFILLER_110_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
XANTENNA__09127__A4 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput95 net95 vssd1 vssd1 vccd1 vccd1 DAT_O[2] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_94_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11076_ clknet_leaf_4_clk _01624_ _00431_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[106\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08335__A2 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10027_ net823 net663 vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__and2_1
XANTENNA__10113__A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_28_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_56_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06897__A2 net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10929_ clknet_leaf_32_clk _01484_ _00284_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.zeroes\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_32_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06120_ top.cw1\[2\] top.cw1\[1\] top.cw1\[0\] vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__nand3_1
XANTENNA__05609__B1 _02695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06282__B1 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06051_ net481 net464 vssd1 vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__or2_2
XANTENNA__08271__B2 top.cb_syn.char_path_n\[32\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_47_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07377__A3 _03547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09810_ net787 net627 vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__and2_1
Xfanout329 _04926_ vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__buf_2
Xfanout307 _02892_ vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__buf_2
Xfanout318 net319 vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__buf_2
XANTENNA__08700__B net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09741_ net778 net618 vssd1 vssd1 vccd1 vccd1 _00355_ sky130_fd_sc_hd__and2_1
X_06953_ top.findLeastValue.val2\[7\] net149 net122 _03618_ vssd1 vssd1 vccd1 vccd1
+ _01949_ sky130_fd_sc_hd__o22a_1
X_05904_ _02877_ _02878_ vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_105_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09672_ net785 net625 vssd1 vssd1 vccd1 vccd1 _00286_ sky130_fd_sc_hd__and2_1
X_06884_ top.compVal\[41\] top.findLeastValue.val1\[41\] net164 vssd1 vssd1 vccd1
+ vccd1 _03584_ sky130_fd_sc_hd__mux2_1
X_08623_ _04833_ _04835_ _04839_ _04826_ net1651 vssd1 vssd1 vccd1 vccd1 _01504_ sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_19_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_8
X_05835_ net171 _02843_ vssd1 vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__and2b_1
X_08554_ net1156 top.cb_syn.char_path_n\[22\] net229 vssd1 vssd1 vccd1 vccd1 _01540_
+ sky130_fd_sc_hd__mux2_1
X_05766_ net473 _02784_ _02786_ top.TRN_sram_complete vssd1 vssd1 vccd1 vccd1 _02787_
+ sky130_fd_sc_hd__or4b_1
XFILLER_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07505_ _04090_ _04095_ _04069_ vssd1 vssd1 vccd1 vccd1 _04096_ sky130_fd_sc_hd__mux2_1
XANTENNA__08428__A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09023__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08485_ net1288 top.cb_syn.char_path_n\[91\] net232 vssd1 vssd1 vccd1 vccd1 _01609_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__05848__B1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11850__Q top.WB.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05697_ net17 net415 net308 top.WB.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 _02361_
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout434_A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07436_ _04020_ _04031_ _03986_ vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__mux2_1
XFILLER_23_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07367_ net1657 net134 _03547_ net126 _03976_ vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_33_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09106_ net458 _02814_ _02803_ vssd1 vssd1 vccd1 vccd1 _05125_ sky130_fd_sc_hd__a21oi_1
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08798__C1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06318_ top.hist_data_o\[11\] top.hist_data_o\[10\] top.hist_data_o\[9\] top.hist_data_o\[8\]
+ vssd1 vssd1 vccd1 vccd1 _03181_ sky130_fd_sc_hd__and4_1
X_09037_ net1176 top.WB.CPU_DAT_O\[20\] net291 vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__mux2_1
X_07298_ _03797_ _03930_ vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__or2_1
X_06249_ _02994_ _03115_ _02574_ vssd1 vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__o21a_1
XANTENNA__06812__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold361 top.hTree.nulls\[56\] vssd1 vssd1 vccd1 vccd1 net1314 sky130_fd_sc_hd__dlygate4sd3_1
Xhold350 top.hTree.nulls\[48\] vssd1 vssd1 vccd1 vccd1 net1303 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout689_X net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold372 net91 vssd1 vssd1 vccd1 vccd1 net1325 sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 top.hTree.nulls\[51\] vssd1 vssd1 vccd1 vccd1 net1347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 top.path\[124\] vssd1 vssd1 vccd1 vccd1 net1336 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout852 net853 vssd1 vssd1 vccd1 vccd1 net852 sky130_fd_sc_hd__clkbuf_2
XFILLER_77_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout841 net842 vssd1 vssd1 vccd1 vccd1 net841 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_5_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout830 net831 vssd1 vssd1 vccd1 vccd1 net830 sky130_fd_sc_hd__clkbuf_2
Xfanout874 net876 vssd1 vssd1 vccd1 vccd1 net874 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout856_X net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_13_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_13_0_clk sky130_fd_sc_hd__clkbuf_8
Xfanout863 net866 vssd1 vssd1 vccd1 vccd1 net863 sky130_fd_sc_hd__clkbuf_2
X_09939_ net787 net627 vssd1 vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__and2_1
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06879__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11832_ clknet_leaf_100_clk _02348_ _01187_ vssd1 vssd1 vccd1 vccd1 top.WB.CPU_DAT_O\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__05551__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07828__A1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07828__B2 top.findLeastValue.sum\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11763_ clknet_leaf_113_clk _02296_ _01118_ vssd1 vssd1 vccd1 vccd1 top.compVal\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__05839__B1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11694_ clknet_leaf_62_clk _02227_ _01049_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10714_ clknet_leaf_3_clk _01313_ _00133_ vssd1 vssd1 vccd1 vccd1 top.path\[90\]
+ sky130_fd_sc_hd__dfrtp_1
X_10645_ clknet_leaf_65_clk _00040_ _00064_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.word_cnt\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10576_ net729 net569 vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_11_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08253__B2 top.cb_syn.char_path_n\[41\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06803__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11128_ clknet_leaf_28_clk _01676_ _00483_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[30\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_3_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11059_ clknet_leaf_26_clk _01607_ _00414_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[89\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_05620_ _02703_ _02704_ net472 vssd1 vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__o21a_1
XANTENNA__09070__C _02530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05551_ top.cb_syn.char_path\[85\] net553 net544 top.cb_syn.char_path\[53\] vssd1
+ vssd1 vccd1 vccd1 _02647_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_50_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05482_ _02552_ _02558_ _02571_ _02586_ vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__o31a_1
X_08270_ top.cb_syn.char_path_n\[34\] net202 _04662_ vssd1 vssd1 vccd1 vccd1 _01680_
+ sky130_fd_sc_hd__o21a_1
X_07221_ net271 _03873_ _03874_ net276 net1570 vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__a32o_1
X_07152_ top.findLeastValue.val1\[21\] top.findLeastValue.val2\[21\] top.findLeastValue.val2\[20\]
+ top.findLeastValue.val1\[20\] vssd1 vssd1 vccd1 vccd1 _03810_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_30_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06103_ top.TRN_char_index\[4\] top.TRN_char_index\[3\] _02974_ vssd1 vssd1 vccd1
+ vccd1 _02976_ sky130_fd_sc_hd__and3_1
XANTENNA__05400__A top.cb_syn.char_index\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_8_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__10018__A net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07083_ _03739_ _03740_ vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__nand2_1
XANTENNA__08795__A2 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09807__A net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06930__S net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06034_ top.hist_data_o\[1\] top.WB.CPU_DAT_O\[1\] net355 vssd1 vssd1 vccd1 vccd1
+ _02176_ sky130_fd_sc_hd__mux2_1
Xfanout137 _02941_ vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__buf_2
Xfanout126 _03549_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__buf_2
XFILLER_59_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09018__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout115 net116 vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__clkbuf_4
Xfanout159 net160 vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__clkbuf_4
X_07985_ _02510_ top.cb_syn.zero_count\[6\] top.cb_syn.zero_count\[5\] _02511_ vssd1
+ vssd1 vccd1 vccd1 _04488_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout384_A net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11845__Q top.WB.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout148 net153 vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__buf_2
X_06936_ top.compVal\[15\] top.findLeastValue.val1\[15\] net161 vssd1 vssd1 vccd1
+ vccd1 _03610_ sky130_fd_sc_hd__mux2_1
X_09724_ net735 net575 vssd1 vssd1 vccd1 vccd1 _00338_ sky130_fd_sc_hd__and2_1
X_09655_ net798 net638 vssd1 vssd1 vccd1 vccd1 _00269_ sky130_fd_sc_hd__and2_1
XFILLER_103_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06867_ net498 _03570_ _03568_ vssd1 vssd1 vccd1 vccd1 _03578_ sky130_fd_sc_hd__a21bo_1
X_08606_ _04138_ _04142_ _04531_ _04824_ vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__and4_1
X_05818_ _02827_ _02834_ vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout551_A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__05533__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09586_ net843 net683 vssd1 vssd1 vccd1 vccd1 _00200_ sky130_fd_sc_hd__and2_1
XFILLER_63_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06798_ top.findLeastValue.val1\[32\] net133 net117 top.compVal\[32\] vssd1 vssd1
+ vccd1 vccd1 _02040_ sky130_fd_sc_hd__o22a_1
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08537_ net1085 top.cb_syn.char_path_n\[39\] net226 vssd1 vssd1 vccd1 vccd1 _01557_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout437_X net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05749_ top.compVal\[45\] net172 net158 top.WB.CPU_DAT_O\[13\] vssd1 vssd1 vccd1
+ vccd1 _02330_ sky130_fd_sc_hd__a22o_1
XFILLER_23_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08468_ net1323 top.cb_syn.char_path_n\[108\] net220 vssd1 vssd1 vccd1 vccd1 _01626_
+ sky130_fd_sc_hd__mux2_1
X_07419_ top.dut.out\[6\] net297 _03999_ _04017_ vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__a22o_1
XFILLER_11_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_10430_ net875 net715 vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_98_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08399_ net517 top.cb_syn.char_path_n\[2\] top.cb_syn.char_path_n\[3\] top.cb_syn.char_path_n\[4\]
+ net513 net509 vssd1 vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__mux4_1
XANTENNA__05310__A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10361_ net874 net714 vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__and2_1
X_10292_ net724 net564 vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__and2_1
XANTENNA__06797__B2 top.compVal\[33\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold180 net97 vssd1 vssd1 vccd1 vccd1 net1133 sky130_fd_sc_hd__dlygate4sd3_1
Xteam_05_910 vssd1 vssd1 vccd1 vccd1 team_05_910/HI gpio_out[25] sky130_fd_sc_hd__conb_1
Xteam_05_921 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] team_05_921/LO sky130_fd_sc_hd__conb_1
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xteam_05_932 vssd1 vssd1 vccd1 vccd1 gpio_oeb[12] team_05_932/LO sky130_fd_sc_hd__conb_1
Xteam_05_943 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] team_05_943/LO sky130_fd_sc_hd__conb_1
Xhold191 top.cb_syn.char_path\[73\] vssd1 vssd1 vccd1 vccd1 net1144 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout660 net663 vssd1 vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__clkbuf_2
Xfanout693 net697 vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__clkbuf_2
Xfanout682 net719 vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__clkbuf_2
Xfanout671 net675 vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__clkbuf_2
XFILLER_19_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08767__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07671__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08171__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11815_ clknet_leaf_56_clk _02331_ _01170_ vssd1 vssd1 vccd1 vccd1 top.TRN_char_index\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_11746_ clknet_leaf_94_clk _02279_ _01101_ vssd1 vssd1 vccd1 vccd1 top.compVal\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11677_ clknet_leaf_61_clk _02210_ _01032_ vssd1 vssd1 vccd1 vccd1 top.sram_interface.init_counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10628_ net805 net645 vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__and2_1
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10559_ net855 net695 vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_58_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06051__A net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07770_ top.findLeastValue.sum\[34\] _04321_ net396 vssd1 vssd1 vccd1 vccd1 _04322_
+ sky130_fd_sc_hd__mux2_1
X_06721_ _02424_ top.findLeastValue.val2\[26\] vssd1 vssd1 vccd1 vccd1 _03509_ sky130_fd_sc_hd__or2_1
X_09440_ net860 net700 vssd1 vssd1 vccd1 vccd1 _00054_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_69_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05515__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06652_ top.controller.fin_FLV top.findLeastValue.histo_index\[8\] net423 _03440_
+ vssd1 vssd1 vccd1 vccd1 _03441_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_35_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09371_ net993 net238 net215 _04302_ vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__a22o_1
X_06583_ _03371_ _03370_ vssd1 vssd1 vccd1 vccd1 _03372_ sky130_fd_sc_hd__nand2b_1
X_05603_ net480 _02689_ net310 top.hTree.node_reg\[45\] vssd1 vssd1 vccd1 vccd1 _02691_
+ sky130_fd_sc_hd__a22o_1
X_05534_ top.cb_syn.char_path\[24\] net559 net314 top.cb_syn.char_path\[120\] vssd1
+ vssd1 vccd1 vccd1 _02633_ sky130_fd_sc_hd__a22o_1
X_08322_ top.cb_syn.char_path_n\[8\] net199 _04688_ vssd1 vssd1 vccd1 vccd1 _01654_
+ sky130_fd_sc_hd__o21a_1
X_08253_ top.cb_syn.char_path_n\[43\] net373 net333 top.cb_syn.char_path_n\[41\] net178
+ vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__a221o_1
X_05465_ top.findLeastValue.wipe_the_char_1 _02548_ vssd1 vssd1 vccd1 vccd1 _02573_
+ sky130_fd_sc_hd__nand2_2
X_07204_ _03659_ _03860_ _03861_ vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout132_A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05396_ net505 vssd1 vssd1 vccd1 vccd1 _02504_ sky130_fd_sc_hd__clkinv_4
X_08184_ top.cb_syn.char_path_n\[77\] net196 _04619_ vssd1 vssd1 vccd1 vccd1 _01723_
+ sky130_fd_sc_hd__o21a_1
XFILLER_20_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05768__C net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07135_ _03788_ _03789_ _03790_ vssd1 vssd1 vccd1 vccd1 _03793_ sky130_fd_sc_hd__or3_1
XFILLER_3_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07066_ _03710_ _03712_ _03709_ vssd1 vssd1 vccd1 vccd1 _03724_ sky130_fd_sc_hd__a21o_1
X_06017_ net1482 top.WB.CPU_DAT_O\[18\] net357 vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_93_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_07968_ net423 _04475_ _04472_ net287 vssd1 vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__o211a_1
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout766_A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09707_ net801 net641 vssd1 vssd1 vccd1 vccd1 _00321_ sky130_fd_sc_hd__and2_1
X_06919_ top.findLeastValue.val2\[24\] net148 net124 _03601_ vssd1 vssd1 vccd1 vccd1
+ _01966_ sky130_fd_sc_hd__o22a_1
X_07899_ top.findLeastValue.sum\[8\] top.hTree.tree_reg\[8\] net278 vssd1 vssd1 vccd1
+ vccd1 _04425_ sky130_fd_sc_hd__mux2_1
X_09638_ net850 net690 vssd1 vssd1 vccd1 vccd1 _00252_ sky130_fd_sc_hd__and2_1
XANTENNA__07900__A0 top.findLeastValue.sum\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09569_ net843 net683 vssd1 vssd1 vccd1 vccd1 _00183_ sky130_fd_sc_hd__and2_1
X_11600_ clknet_leaf_61_clk _02148_ _00955_ vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11531_ clknet_leaf_5_clk _02079_ _00886_ vssd1 vssd1 vccd1 vccd1 top.histogram.total\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06781__D net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11462_ clknet_leaf_93_clk _02010_ _00817_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val1\[2\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_11_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10413_ net796 net636 vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__and2_1
XANTENNA__05690__A1 net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05690__B2 top.WB.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11393_ clknet_leaf_83_clk _01941_ _00748_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_99_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10344_ net871 net711 vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__and2_1
XANTENNA__08351__A net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10275_ net726 net566 vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__and2_1
Xfanout490 net491 vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_100_Left_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_105_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload8_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_11729_ clknet_leaf_122_clk _02262_ _01084_ vssd1 vssd1 vccd1 vccd1 top.path\[60\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_40_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05681__B2 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07576__S _04144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07958__A0 top.findLeastValue.least1\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09076__B net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08940_ top.WB.CPU_DAT_O\[14\] net1084 net372 vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__mux2_1
X_08871_ top.translation.index\[4\] _05049_ _05045_ vssd1 vssd1 vccd1 vccd1 _01466_
+ sky130_fd_sc_hd__a21o_1
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07822_ net427 _04362_ _04363_ net259 vssd1 vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__o211a_1
XFILLER_29_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07605__A net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07753_ net443 net1606 net255 net1732 _04308_ vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__a221o_1
X_07684_ net491 _04249_ vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__or2_1
XANTENNA__07489__A2 top.cb_syn.char_path_n\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06704_ _02431_ top.findLeastValue.val2\[18\] top.findLeastValue.val2\[17\] _02432_
+ vssd1 vssd1 vccd1 vccd1 _03492_ sky130_fd_sc_hd__a22o_1
XFILLER_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09423_ top.hTree.nulls\[62\] _04204_ net407 vssd1 vssd1 vccd1 vccd1 _05292_ sky130_fd_sc_hd__mux2_1
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06635_ _03388_ _03413_ _03422_ vssd1 vssd1 vccd1 vccd1 _03424_ sky130_fd_sc_hd__a21o_4
X_09354_ net1009 net241 net217 _04370_ vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__a22o_1
XANTENNA__08438__A1 _02504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08305_ top.cb_syn.char_path_n\[17\] net375 net335 top.cb_syn.char_path_n\[15\] net180
+ vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__a221o_1
X_06566_ top.findLeastValue.val1\[1\] top.compVal\[1\] vssd1 vssd1 vccd1 vccd1 _03355_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_21_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09285_ _04000_ _04030_ vssd1 vssd1 vccd1 vccd1 top.dut.bit_buf_next\[3\] sky130_fd_sc_hd__and2_1
X_05517_ _02617_ _02618_ net476 vssd1 vssd1 vccd1 vccd1 _02619_ sky130_fd_sc_hd__o21a_1
XANTENNA__07379__A2_N net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout514_A top.cb_syn.end_cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06497_ _03284_ _03304_ vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__nor2_1
X_05448_ net479 net548 _02555_ vssd1 vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__and3_1
X_08236_ top.cb_syn.char_path_n\[51\] net198 _04645_ vssd1 vssd1 vccd1 vccd1 _01697_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_95_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08167_ top.cb_syn.char_path_n\[86\] net387 net346 top.cb_syn.char_path_n\[84\] net191
+ vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout302_X net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07118_ _03770_ _03772_ _03774_ _03736_ vssd1 vssd1 vccd1 vccd1 _03776_ sky130_fd_sc_hd__a211o_1
X_05379_ top.findLeastValue.val2\[27\] vssd1 vssd1 vccd1 vccd1 _02487_ sky130_fd_sc_hd__inv_2
XFILLER_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08098_ top.cb_syn.char_path_n\[120\] net204 _04576_ vssd1 vssd1 vccd1 vccd1 _01766_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07049_ _03679_ _03676_ vssd1 vssd1 vccd1 vccd1 _03707_ sky130_fd_sc_hd__nand2b_1
X_10060_ net849 net689 vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__and2_1
XANTENNA__08913__A2 _04187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10962_ clknet_leaf_52_clk _01510_ _00317_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_index\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_90_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10893_ clknet_leaf_12_clk _01470_ _00248_ vssd1 vssd1 vccd1 vccd1 top.translation.writeEn
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08429__A1 _02506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11514_ clknet_leaf_69_clk _02062_ _00869_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.least1\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_11_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08780__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11445_ clknet_leaf_69_clk _01993_ _00800_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.histo_index\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05663__B2 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11376_ clknet_leaf_81_clk _01924_ _00731_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10327_ net792 net632 vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__and2_1
X_10258_ net865 net705 vssd1 vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__and2_1
XFILLER_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10189_ net864 net704 vssd1 vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__and2_1
XFILLER_66_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05718__A2 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06420_ top.header_synthesis.write_char_path top.header_synthesis.start vssd1 vssd1
+ vccd1 vccd1 _03251_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_45_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09093__A1 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06351_ net1177 _03206_ net302 vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__mux2_1
X_09070_ top.cb_syn.wait_cycle _02553_ _02530_ top.cb_syn.h_element\[54\] vssd1 vssd1
+ vccd1 vccd1 _05094_ sky130_fd_sc_hd__or4b_1
X_06282_ _03138_ _03142_ _03147_ net159 vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__o31a_1
X_05302_ top.compVal\[39\] vssd1 vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__inv_2
X_08021_ _02501_ _04515_ vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__nand2_1
Xhold702 top.sram_interface.zero_cnt\[1\] vssd1 vssd1 vccd1 vccd1 net1655 sky130_fd_sc_hd__dlygate4sd3_1
Xhold735 top.cb_syn.num_lefts\[3\] vssd1 vssd1 vccd1 vccd1 net1688 sky130_fd_sc_hd__dlygate4sd3_1
Xhold724 top.cb_syn.count\[4\] vssd1 vssd1 vccd1 vccd1 net1677 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_77_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold746 top.compVal\[28\] vssd1 vssd1 vccd1 vccd1 net1699 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07159__X _03817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold713 top.hist_data_o\[13\] vssd1 vssd1 vccd1 vccd1 net1666 sky130_fd_sc_hd__dlygate4sd3_1
X_09972_ net776 net616 vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__and2_1
Xhold757 top.findLeastValue.sum\[32\] vssd1 vssd1 vccd1 vccd1 net1710 sky130_fd_sc_hd__dlygate4sd3_1
Xhold779 top.findLeastValue.sum\[38\] vssd1 vssd1 vccd1 vccd1 net1732 sky130_fd_sc_hd__dlygate4sd3_1
Xhold768 top.histogram.total\[26\] vssd1 vssd1 vccd1 vccd1 net1721 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10026__A net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09148__A2 _02530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08923_ top.WB.CPU_DAT_O\[31\] net1439 net372 vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__mux2_1
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07606__Y _04190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08854_ net431 top.header_synthesis.enable _05036_ top.controller.state_reg\[5\]
+ net36 vssd1 vssd1 vccd1 vccd1 _05037_ sky130_fd_sc_hd__o2111a_1
XANTENNA__05709__A2 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05997_ _02905_ _02923_ vssd1 vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__nor2_1
XFILLER_84_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07805_ top.hTree.tree_reg\[27\] top.findLeastValue.sum\[27\] net249 vssd1 vssd1
+ vccd1 vccd1 _04350_ sky130_fd_sc_hd__mux2_1
XANTENNA__11853__Q top.WB.CPU_DAT_O\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08785_ net433 _04966_ _04967_ vssd1 vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout464_A net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09305__C1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07736_ net488 _04293_ vssd1 vssd1 vccd1 vccd1 _04295_ sky130_fd_sc_hd__or2_1
XFILLER_111_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06134__A2 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout631_A net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07667_ top.findLeastValue.least2\[8\] net394 net248 top.hTree.tree_reg\[54\] net485
+ vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__o221a_1
XFILLER_52_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07867__C1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07598_ top.cb_syn.h_element\[55\] top.cb_syn.h_element\[46\] _04145_ vssd1 vssd1
+ vccd1 vccd1 _04183_ sky130_fd_sc_hd__mux2_1
X_09406_ net407 _04231_ vssd1 vssd1 vccd1 vccd1 _05281_ sky130_fd_sc_hd__nand2_1
X_06618_ _03393_ _03405_ _03406_ _03395_ vssd1 vssd1 vccd1 vccd1 _03407_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_23_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06549_ _03329_ _03337_ _03328_ vssd1 vssd1 vccd1 vccd1 _03338_ sky130_fd_sc_hd__o21a_1
X_09337_ net1035 net236 net214 _04438_ vssd1 vssd1 vccd1 vccd1 _01399_ sky130_fd_sc_hd__a22o_1
X_09268_ _05213_ _05220_ _05221_ _05214_ net1632 vssd1 vssd1 vccd1 vccd1 top.header_synthesis.next_zero_count\[3\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout517_X net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08219_ top.cb_syn.char_path_n\[60\] net386 net345 top.cb_syn.char_path_n\[58\] net190
+ vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__a221o_1
XANTENNA__08831__B2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09199_ top.hTree.state\[4\] _05062_ net264 vssd1 vssd1 vccd1 vccd1 _00022_ sky130_fd_sc_hd__mux2_1
XANTENNA__06842__B1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_40_12
X_11230_ clknet_leaf_35_clk _01778_ _00585_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.end_cnt\[3\]
+ sky130_fd_sc_hd__dfstp_1
X_11161_ clknet_leaf_18_clk _01709_ _00516_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_96_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07493__S1 _04071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10112_ net812 net652 vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__and2_1
X_11092_ clknet_leaf_29_clk _01640_ _00447_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_88_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10043_ net839 net679 vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__and2_1
Xhold40 top.hTree.node_reg\[39\] vssd1 vssd1 vccd1 vccd1 net993 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 net50 vssd1 vssd1 vccd1 vccd1 net1026 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input25_A DAT_I[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold62 top.hTree.tree_reg\[47\] vssd1 vssd1 vccd1 vccd1 net1015 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 top.hTree.node_reg\[24\] vssd1 vssd1 vccd1 vccd1 net1004 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 net58 vssd1 vssd1 vccd1 vccd1 net1037 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06373__A2 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold95 top.histogram.sram_out\[12\] vssd1 vssd1 vccd1 vccd1 net1048 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05581__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10945_ clknet_leaf_33_clk _01500_ _00300_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.num_lefts\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_10876_ clknet_leaf_36_clk _00007_ _00231_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.curr_state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08076__A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08822__B2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06833__B1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08035__C1 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11428_ clknet_leaf_86_clk _01976_ _00783_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.val2\[34\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_4 top.WB.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11359_ clknet_leaf_97_clk _01907_ _00714_ vssd1 vssd1 vccd1 vccd1 top.findLeastValue.sum\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_98_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__07484__S1 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07854__S net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05920_ top.sram_interface.TRN_counter\[2\] top.sram_interface.TRN_counter\[1\] vssd1
+ vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_72_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05851_ top.compVal\[16\] net168 net154 top.WB.CPU_DAT_O\[16\] vssd1 vssd1 vccd1
+ vccd1 _02291_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_6_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07561__B2 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07561__A1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08570_ net1147 top.cb_syn.char_path_n\[6\] net226 vssd1 vssd1 vccd1 vccd1 _01524_
+ sky130_fd_sc_hd__mux2_1
X_07521_ top.cb_syn.curr_path\[127\] top.cb_syn.char_path_n\[127\] top.cb_syn.char_path_n\[126\]
+ top.cb_syn.char_path_n\[125\] net401 net352 vssd1 vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__mux4_1
X_05782_ top.hTree.write_HT_fin net430 _02801_ vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__or3_1
XANTENNA__07313__B2 top.findLeastValue.sum\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07313__A1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07452_ top.findLeastValue.startup net423 net288 vssd1 vssd1 vccd1 vccd1 _01879_
+ sky130_fd_sc_hd__a21o_1
XFILLER_50_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07383_ net354 vssd1 vssd1 vccd1 vccd1 top.dut.bits_in_buf_next\[1\] sky130_fd_sc_hd__inv_2
X_06403_ top.hist_data_o\[4\] _03174_ vssd1 vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__nor2_1
X_09122_ net451 net548 net463 _05137_ vssd1 vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__a31o_1
X_06334_ top.hist_data_o\[23\] top.hist_data_o\[22\] _03189_ vssd1 vssd1 vccd1 vccd1
+ _03196_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_20_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06265_ net502 _03011_ vssd1 vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__xnor2_1
X_09053_ net1221 top.WB.CPU_DAT_O\[4\] net293 vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__mux2_1
X_08004_ _04503_ _04506_ _04504_ _04496_ vssd1 vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__o211a_2
X_06196_ net500 _02767_ _03014_ _03064_ vssd1 vssd1 vccd1 vccd1 _03065_ sky130_fd_sc_hd__o2bb2a_1
Xhold510 top.hTree.tree_reg\[1\] vssd1 vssd1 vccd1 vccd1 net1463 sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 top.cb_syn.left vssd1 vssd1 vccd1 vccd1 net1507 sky130_fd_sc_hd__dlygate4sd3_1
Xhold521 top.cb_syn.curr_index\[6\] vssd1 vssd1 vccd1 vccd1 net1474 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11848__Q top.WB.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold543 top.hist_data_o\[5\] vssd1 vssd1 vccd1 vccd1 net1496 sky130_fd_sc_hd__dlygate4sd3_1
Xhold532 top.hist_data_o\[7\] vssd1 vssd1 vccd1 vccd1 net1485 sky130_fd_sc_hd__dlygate4sd3_1
Xhold576 top.cb_syn.cb_enable vssd1 vssd1 vccd1 vccd1 net1529 sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 top.cb_syn.char_path\[127\] vssd1 vssd1 vccd1 vccd1 net1518 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07617__X _04198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold587 _01830_ vssd1 vssd1 vccd1 vccd1 net1540 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_106_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09955_ net769 net609 vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__and2_1
Xhold598 top.hTree.tree_reg\[23\] vssd1 vssd1 vccd1 vccd1 net1551 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout581_A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08906_ _04187_ _05067_ _05074_ _05073_ _05072_ vssd1 vssd1 vccd1 vccd1 _05075_ sky130_fd_sc_hd__o311a_1
X_09886_ net745 net585 vssd1 vssd1 vccd1 vccd1 _00500_ sky130_fd_sc_hd__and2_1
X_08837_ net522 _05010_ _02522_ vssd1 vssd1 vccd1 vccd1 _05020_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout846_A net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06760__C1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05563__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08768_ top.path\[80\] net409 net327 top.path\[81\] net436 vssd1 vssd1 vccd1 vccd1
+ _04951_ sky130_fd_sc_hd__o221a_1
X_08699_ _04875_ _04885_ _02516_ vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07719_ top.findLeastValue.sum\[44\] top.hTree.tree_reg\[44\] net283 vssd1 vssd1
+ vccd1 vccd1 _04281_ sky130_fd_sc_hd__mux2_1
X_10730_ clknet_leaf_112_clk _01329_ _00149_ vssd1 vssd1 vccd1 vccd1 top.path\[106\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09057__A1 top.WB.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05866__B2 top.WB.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10661_ clknet_leaf_118_clk _01260_ _00080_ vssd1 vssd1 vccd1 vccd1 top.path\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07939__S net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06843__S _03424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10592_ net747 net587 vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__and2_1
XANTENNA__05967__B _02581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06815__B1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06144__A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11213_ clknet_leaf_23_clk _01761_ _00568_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[115\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput52 net52 vssd1 vssd1 vccd1 vccd1 ADR_O[17] sky130_fd_sc_hd__buf_2
Xoutput63 net63 vssd1 vssd1 vccd1 vccd1 ADR_O[29] sky130_fd_sc_hd__buf_2
Xoutput85 net85 vssd1 vssd1 vccd1 vccd1 DAT_O[20] sky130_fd_sc_hd__buf_2
X_11144_ clknet_leaf_8_clk _01692_ _00499_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path_n\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_8_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 DAT_O[10] sky130_fd_sc_hd__buf_2
Xoutput96 net96 vssd1 vssd1 vccd1 vccd1 DAT_O[30] sky130_fd_sc_hd__buf_2
XFILLER_110_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__09174__B net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11075_ clknet_leaf_10_clk _01623_ _00430_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.char_path\[105\]
+ sky130_fd_sc_hd__dfrtp_1
X_10026_ net822 net662 vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__and2_1
XFILLER_36_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10928_ clknet_leaf_31_clk _01483_ _00283_ vssd1 vssd1 vccd1 vccd1 top.cb_syn.zeroes\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05857__B2 top.WB.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10859_ clknet_leaf_77_clk _01445_ vssd1 vssd1 vccd1 vccd1 top.hTree.node_reg\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09048__A1 top.WB.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07849__S net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06806__B1 net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06050_ net1043 _02592_ net160 vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__a21o_1
XANTENNA__06054__A net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06034__A1 top.WB.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout308 net309 vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__buf_2
Xfanout319 net320 vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__clkbuf_4
X_09740_ net778 net618 vssd1 vssd1 vccd1 vccd1 _00354_ sky130_fd_sc_hd__and2_1
XFILLER_98_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07782__A1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06952_ top.compVal\[7\] top.findLeastValue.val1\[7\] net164 vssd1 vssd1 vccd1 vccd1
+ _03618_ sky130_fd_sc_hd__mux2_1
.ends

