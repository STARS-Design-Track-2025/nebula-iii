* NGSPICE file created from team_02.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

.subckt team_02 clk en gpio_in[0] gpio_in[10] gpio_in[11] gpio_in[12] gpio_in[13]
+ gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17] gpio_in[18] gpio_in[19] gpio_in[1]
+ gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23] gpio_in[24] gpio_in[25] gpio_in[26]
+ gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2] gpio_in[30] gpio_in[31] gpio_in[32]
+ gpio_in[33] gpio_in[3] gpio_in[4] gpio_in[5] gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9]
+ gpio_oeb[0] gpio_oeb[10] gpio_oeb[11] gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15]
+ gpio_oeb[16] gpio_oeb[17] gpio_oeb[18] gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21]
+ gpio_oeb[22] gpio_oeb[23] gpio_oeb[24] gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28]
+ gpio_oeb[29] gpio_oeb[2] gpio_oeb[30] gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[3]
+ gpio_oeb[4] gpio_oeb[5] gpio_oeb[6] gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0]
+ gpio_out[10] gpio_out[11] gpio_out[12] gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16]
+ gpio_out[17] gpio_out[18] gpio_out[19] gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22]
+ gpio_out[23] gpio_out[24] gpio_out[25] gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29]
+ gpio_out[2] gpio_out[30] gpio_out[31] gpio_out[32] gpio_out[33] gpio_out[3] gpio_out[4]
+ gpio_out[5] gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9] nrst vccd1 vssd1
X_2106_ dut.data_in\[3\] _0515_ vssd1 vssd1 vccd1 vccd1 _0523_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_37_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2037_ _0973_ _0474_ _0475_ vssd1 vssd1 vccd1 vccd1 _0012_ sky130_fd_sc_hd__and3_1
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout75_A net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1606_ _0913_ _1187_ _1189_ _1191_ _1194_ vssd1 vssd1 vccd1 vccd1 _1195_ sky130_fd_sc_hd__a311o_1
X_2724_ clknet_leaf_4_clk _0094_ net67 vssd1 vssd1 vccd1 vccd1 dut.microstep_y.ctr\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_2655_ clknet_leaf_25_clk _0126_ net60 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.bit_count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1399_ dut.lcd1602.cnt_200ms\[5\] dut.lcd1602.cnt_200ms\[4\] _1002_ vssd1 vssd1 vccd1
+ vccd1 _1003_ sky130_fd_sc_hd__and3_1
X_1537_ _1119_ _1125_ vssd1 vssd1 vccd1 vccd1 _1126_ sky130_fd_sc_hd__nand2_1
X_1468_ dut.actual_duty_y\[3\] _1046_ _1056_ vssd1 vssd1 vccd1 vccd1 _1057_ sky130_fd_sc_hd__nand3_1
X_2586_ dut.ir_sensor_array.final_sensor_data\[30\] _0883_ dut.ir_sensor_array.final_sensor_data\[29\]
+ vssd1 vssd1 vccd1 vccd1 _0884_ sky130_fd_sc_hd__o21ba_1
XFILLER_27_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xteam_02_95 vssd1 vssd1 vccd1 vccd1 team_02_95/HI gpio_oeb[11] sky130_fd_sc_hd__conb_1
XFILLER_50_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold170 dut.lcd1602.cnt_200ms\[13\] vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2440_ _0775_ _0785_ vssd1 vssd1 vccd1 vccd1 _0792_ sky130_fd_sc_hd__nand2_1
X_2371_ net300 _1003_ vssd1 vssd1 vccd1 vccd1 _0745_ sky130_fd_sc_hd__nor2_1
X_1322_ _0940_ net32 vssd1 vssd1 vccd1 vccd1 _0944_ sky130_fd_sc_hd__nand2_1
XFILLER_64_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2638_ clknet_leaf_15_clk _0109_ net83 vssd1 vssd1 vccd1 vccd1 dut.sdo_lcd sky130_fd_sc_hd__dfrtp_1
X_2569_ net274 dut.ir_sensor_array.final_sensor_data\[34\] net34 vssd1 vssd1 vccd1
+ vccd1 _0217_ sky130_fd_sc_hd__mux2_1
X_2707_ clknet_2_2__leaf_clk dut.pwm_a_inst_x.count_d\[10\] net78 vssd1 vssd1 vccd1
+ vccd1 dut.pwm_a_inst_x.count_q\[10\] sky130_fd_sc_hd__dfrtp_4
XFILLER_55_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1940_ net280 _0417_ vssd1 vssd1 vccd1 vccd1 _0418_ sky130_fd_sc_hd__nor2_1
XFILLER_9_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1871_ _0376_ net26 _0375_ vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_x.count_d\[11\]
+ sky130_fd_sc_hd__and3b_1
X_2423_ _0766_ _0772_ vssd1 vssd1 vccd1 vccd1 _0775_ sky130_fd_sc_hd__or2_1
X_2354_ _0705_ _0720_ dut.microstep_x.clk_en vssd1 vssd1 vccd1 vccd1 _0737_ sky130_fd_sc_hd__o21ai_1
X_1305_ net2 vssd1 vssd1 vccd1 vccd1 _0929_ sky130_fd_sc_hd__inv_2
X_2285_ _0666_ _0512_ vssd1 vssd1 vccd1 vccd1 _0673_ sky130_fd_sc_hd__and2b_1
XFILLER_37_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2070_ _0976_ _0494_ vssd1 vssd1 vccd1 vccd1 dut.cs_n_lcd sky130_fd_sc_hd__nor2_1
XFILLER_38_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1923_ net17 _0407_ vssd1 vssd1 vccd1 vccd1 _0408_ sky130_fd_sc_hd__nor2_1
X_1785_ _1257_ _0287_ _0289_ vssd1 vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__nor3_1
X_1854_ _0327_ _0361_ vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__and2_1
X_2406_ _0764_ net214 vssd1 vssd1 vccd1 vccd1 _0160_ sky130_fd_sc_hd__nor2_1
X_2199_ _0581_ _0600_ vssd1 vssd1 vccd1 vccd1 _0602_ sky130_fd_sc_hd__nand2_1
XFILLER_29_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2268_ _0939_ _0653_ dut.ir_sensor_array.bit_count\[3\] vssd1 vssd1 vccd1 vccd1 _0659_
+ sky130_fd_sc_hd__a21o_1
X_2337_ dut.actual_duty_x\[0\] _0724_ dut.microstep_x.clk_en vssd1 vssd1 vccd1 vccd1
+ _0132_ sky130_fd_sc_hd__mux2_1
XFILLER_52_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold52 dut.lcd1602.cnt_200ms\[14\] vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 dut.lcd1602.cnt_200ms\[7\] vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 dut.microstep_x.ctr\[26\] vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 dut.clkdiv_inst.counter\[1\] vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 dut.ir_sensor_array.bit_count\[5\] vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 dut.pwm_a_inst_y.count_q\[7\] vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 dut.ir_sensor_array.final_sensor_data\[33\] vssd1 vssd1 vccd1 vccd1 net248
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1570_ _1073_ _1087_ _1140_ vssd1 vssd1 vccd1 vccd1 _1159_ sky130_fd_sc_hd__or3_1
XFILLER_6_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2122_ dut.lcd1602.out_valid _0514_ _0529_ _0531_ _0984_ vssd1 vssd1 vccd1 vccd1
+ _0532_ sky130_fd_sc_hd__o2111a_1
X_2053_ net276 _0484_ vssd1 vssd1 vccd1 vccd1 _0003_ sky130_fd_sc_hd__xor2_1
XFILLER_13_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1906_ _0910_ _0389_ _0397_ vssd1 vssd1 vccd1 vccd1 _0095_ sky130_fd_sc_hd__a21oi_1
X_2886_ clknet_leaf_5_clk _0007_ net62 vssd1 vssd1 vccd1 vccd1 dut.clkdiv_inst.counter\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1837_ dut.pwm_a_inst_x.count_q\[18\] dut.pwm_a_inst_x.count_q\[19\] _0354_ vssd1
+ vssd1 vccd1 vccd1 _0355_ sky130_fd_sc_hd__nor3_1
X_1768_ _0235_ _0285_ _1273_ vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__a21o_1
X_1699_ _1243_ _1244_ _1252_ vssd1 vssd1 vccd1 vccd1 _1269_ sky130_fd_sc_hd__o21ai_1
XFILLER_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput7 net7 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__buf_2
XFILLER_16_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2671_ clknet_leaf_9_clk _0034_ net70 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_500hz\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_1622_ dut.pwm_a_inst_y.count_q\[14\] _1209_ _1210_ dut.pwm_a_inst_y.count_q\[19\]
+ dut.pwm_a_inst_y.count_q\[18\] vssd1 vssd1 vccd1 vccd1 _1211_ sky130_fd_sc_hd__a2111o_1
X_2740_ clknet_leaf_6_clk _0082_ net62 vssd1 vssd1 vccd1 vccd1 dut.microstep_y.ctr\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2812__RESET_B net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1553_ _1050_ _1052_ _1053_ _1058_ vssd1 vssd1 vccd1 vccd1 _1142_ sky130_fd_sc_hd__a211oi_1
X_1484_ _1062_ _1071_ vssd1 vssd1 vccd1 vccd1 _1073_ sky130_fd_sc_hd__xnor2_1
XFILLER_39_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2105_ dut.spi.shift_reg_q\[1\] net20 _0520_ net246 _0522_ vssd1 vssd1 vccd1 vccd1
+ _0102_ sky130_fd_sc_hd__o221a_1
XFILLER_39_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2036_ dut.clkdiv_inst.counter\[3\] _0969_ vssd1 vssd1 vccd1 vccd1 _0475_ sky130_fd_sc_hd__or2_1
XFILLER_22_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2869_ clknet_leaf_12_clk _0222_ net79 vssd1 vssd1 vccd1 vccd1 dut.ball_pos_x\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout68_A net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_5_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2723_ clknet_leaf_4_clk _0093_ net67 vssd1 vssd1 vccd1 vccd1 dut.microstep_y.ctr\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_2654_ clknet_leaf_14_clk _0125_ vssd1 vssd1 vccd1 vccd1 dut.data_in\[9\] sky130_fd_sc_hd__dfxtp_1
X_1536_ _1120_ _1124_ vssd1 vssd1 vccd1 vccd1 _1125_ sky130_fd_sc_hd__and2_1
X_1605_ dut.pwm_a_inst_y.count_q\[2\] _1185_ _1193_ dut.pwm_a_inst_y.count_q\[3\]
+ vssd1 vssd1 vccd1 vccd1 _1194_ sky130_fd_sc_hd__o22ai_1
X_2585_ dut.ir_sensor_array.final_sensor_data\[16\] _0882_ dut.ir_sensor_array.final_sensor_data\[31\]
+ vssd1 vssd1 vccd1 vccd1 _0883_ sky130_fd_sc_hd__o21ba_1
X_1398_ dut.lcd1602.cnt_200ms\[3\] _1001_ vssd1 vssd1 vccd1 vccd1 _1002_ sky130_fd_sc_hd__and2_1
X_1467_ net36 net37 vssd1 vssd1 vccd1 vccd1 _1056_ sky130_fd_sc_hd__or2_2
Xteam_02_96 vssd1 vssd1 vccd1 vccd1 team_02_96/HI gpio_oeb[12] sky130_fd_sc_hd__conb_1
XFILLER_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2019_ _0464_ _0465_ vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_19_Left_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold160 dut.lcd1602.cnt_500hz\[11\] vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 dut.ir_sensor_array.final_sensor_data\[25\] vssd1 vssd1 vccd1 vccd1 net323
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_56_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2370_ _1003_ _0744_ net13 vssd1 vssd1 vccd1 vccd1 _0145_ sky130_fd_sc_hd__o21ai_1
X_1321_ net35 dut.ir_sensor_array.state\[1\] vssd1 vssd1 vccd1 vccd1 _0943_ sky130_fd_sc_hd__nand2_2
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_19_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2706_ clknet_leaf_21_clk dut.pwm_a_inst_x.count_d\[9\] net78 vssd1 vssd1 vccd1 vccd1
+ dut.pwm_a_inst_x.count_q\[9\] sky130_fd_sc_hd__dfrtp_2
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2637_ clknet_leaf_13_clk net178 net82 vssd1 vssd1 vccd1 vccd1 dut.spi.shift_reg_q\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_1519_ dut.actual_duty_y\[3\] net41 vssd1 vssd1 vccd1 vccd1 _1108_ sky130_fd_sc_hd__and2_1
X_2568_ net301 net248 net34 vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__mux2_1
X_2499_ _0817_ _0830_ net44 vssd1 vssd1 vccd1 vccd1 _0845_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1870_ dut.pwm_a_inst_x.count_q\[10\] dut.pwm_a_inst_x.count_q\[11\] _0372_ vssd1
+ vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__and3_1
XFILLER_43_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2422_ _0769_ _0773_ dut.pid_y.y_pid.last_error\[3\] vssd1 vssd1 vccd1 vccd1 _0774_
+ sky130_fd_sc_hd__o21ai_1
X_2353_ _0696_ _0722_ _0728_ vssd1 vssd1 vccd1 vccd1 _0736_ sky130_fd_sc_hd__a21oi_1
XFILLER_49_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1304_ dut.ir_sensor_array.final_sensor_data\[1\] vssd1 vssd1 vccd1 vccd1 _0928_
+ sky130_fd_sc_hd__inv_2
X_2284_ _0669_ _0670_ vssd1 vssd1 vccd1 vccd1 _0672_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1999_ _0453_ vssd1 vssd1 vccd1 vccd1 _0454_ sky130_fd_sc_hd__inv_2
XFILLER_55_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1922_ dut.microstep_y.ctr\[15\] _0405_ vssd1 vssd1 vccd1 vccd1 _0407_ sky130_fd_sc_hd__and2_1
X_1853_ dut.pwm_a_inst_x.count_q\[5\] _0363_ vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__or2_1
X_1784_ _0295_ _0301_ _0297_ vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__a21bo_1
X_2405_ dut.lcd1602.cnt_200ms\[19\] _0762_ net213 vssd1 vssd1 vccd1 vccd1 _0765_ sky130_fd_sc_hd__a21oi_1
X_2336_ _0922_ _0672_ _0723_ vssd1 vssd1 vccd1 vccd1 _0724_ sky130_fd_sc_hd__mux2_1
XFILLER_52_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2198_ net12 _0571_ vssd1 vssd1 vccd1 vccd1 _0601_ sky130_fd_sc_hd__nand2_1
X_2267_ net210 _0656_ _0658_ vssd1 vssd1 vccd1 vccd1 _0128_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_35_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold75 dut.lcd1602.cnt_200ms\[5\] vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 dut.lcd1602.cnt_200ms\[13\] vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 dut.lcd1602.cnt_200ms\[0\] vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 dut.microstep_y.ctr\[24\] vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 dut.spi.shift_reg_q\[4\] vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 dut.microstep_y.ctr\[20\] vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 dut.microstep_y.ctr\[14\] vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 _0385_ vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_43_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2121_ dut.spi.bit_counter_q\[0\] dut.spi.bit_counter_q\[3\] _0530_ _0977_ vssd1
+ vssd1 vccd1 vccd1 _0531_ sky130_fd_sc_hd__a31o_1
XFILLER_34_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2052_ _0019_ _0483_ _0484_ vssd1 vssd1 vccd1 vccd1 _0018_ sky130_fd_sc_hd__nor3_1
XFILLER_19_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1905_ _0066_ _0396_ vssd1 vssd1 vccd1 vccd1 _0397_ sky130_fd_sc_hd__or2_1
XFILLER_34_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2885_ clknet_leaf_5_clk _0006_ net53 vssd1 vssd1 vccd1 vccd1 dut.clkdiv_inst.counter\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_1698_ _1265_ _1267_ vssd1 vssd1 vccd1 vccd1 _1268_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1767_ _0237_ _0284_ vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__or2_1
X_1836_ _0301_ _0352_ _0353_ dut.pwm_a_inst_x.count_q\[16\] dut.pwm_a_inst_x.count_q\[17\]
+ vssd1 vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__o311a_1
X_2319_ _0921_ _0687_ vssd1 vssd1 vccd1 vccd1 _0707_ sky130_fd_sc_hd__or2_1
XFILLER_25_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput8 net8 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_33_Left_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput10 net10 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__buf_2
XFILLER_0_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2670_ clknet_leaf_10_clk _0033_ net71 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_500hz\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_1621_ dut.pwm_a_inst_y.count_q\[17\] dut.pwm_a_inst_y.count_q\[16\] dut.pwm_a_inst_y.count_q\[15\]
+ vssd1 vssd1 vccd1 vccd1 _1210_ sky130_fd_sc_hd__or3_1
X_1552_ _1087_ _1140_ _1073_ vssd1 vssd1 vccd1 vccd1 _1141_ sky130_fd_sc_hd__o21ai_1
XFILLER_8_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2104_ dut.data_in\[2\] _0515_ vssd1 vssd1 vccd1 vccd1 _0522_ sky130_fd_sc_hd__or2_1
X_1483_ _1071_ _1062_ vssd1 vssd1 vccd1 vccd1 _1072_ sky130_fd_sc_hd__nand2b_1
X_2035_ dut.clkdiv_inst.counter\[3\] _0969_ vssd1 vssd1 vccd1 vccd1 _0474_ sky130_fd_sc_hd__nand2_1
X_2868_ clknet_leaf_4_clk _0221_ net68 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[39\]
+ sky130_fd_sc_hd__dfrtp_1
X_2799_ clknet_leaf_8_clk _0153_ net64 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_200ms\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_1819_ _0275_ _0336_ _0335_ dut.pwm_a_inst_x.count_q\[3\] vssd1 vssd1 vccd1 vccd1
+ _0337_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_43_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_51_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2722_ clknet_leaf_4_clk _0092_ net67 vssd1 vssd1 vccd1 vccd1 dut.microstep_y.ctr\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2653_ clknet_leaf_13_clk _0124_ vssd1 vssd1 vccd1 vccd1 dut.data_in\[7\] sky130_fd_sc_hd__dfxtp_1
X_1535_ dut.actual_duty_y\[1\] _1108_ _1109_ vssd1 vssd1 vccd1 vccd1 _1124_ sky130_fd_sc_hd__o21a_1
X_1604_ dut.actual_duty_y\[3\] _1192_ vssd1 vssd1 vccd1 vccd1 _1193_ sky130_fd_sc_hd__xnor2_1
X_2584_ dut.ir_sensor_array.final_sensor_data\[18\] _0881_ dut.ir_sensor_array.final_sensor_data\[17\]
+ vssd1 vssd1 vccd1 vccd1 _0882_ sky130_fd_sc_hd__o21ba_1
X_1397_ dut.lcd1602.cnt_200ms\[0\] dut.lcd1602.cnt_200ms\[1\] dut.lcd1602.cnt_200ms\[2\]
+ vssd1 vssd1 vccd1 vccd1 _1001_ sky130_fd_sc_hd__and3_1
X_1466_ _1043_ _1054_ vssd1 vssd1 vccd1 vccd1 _1055_ sky130_fd_sc_hd__nand2_1
Xteam_02_97 vssd1 vssd1 vccd1 vccd1 team_02_97/HI gpio_oeb[13] sky130_fd_sc_hd__conb_1
X_2018_ dut.microstep_x.ctr\[23\] dut.microstep_x.ctr\[24\] _0463_ vssd1 vssd1 vccd1
+ vccd1 _0465_ sky130_fd_sc_hd__and3_1
Xhold150 dut.lcd1602.cnt_500hz\[3\] vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout80_A net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold161 dut.pwm_a_inst_x.count_q\[17\] vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_5_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1320_ net35 dut.ir_sensor_array.state\[1\] vssd1 vssd1 vccd1 vccd1 _0942_ sky130_fd_sc_hd__and2_1
XFILLER_64_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Left_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2636_ clknet_leaf_15_clk net229 net82 vssd1 vssd1 vccd1 vccd1 dut.spi.shift_reg_q\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2705_ clknet_leaf_21_clk dut.pwm_a_inst_x.count_d\[8\] net76 vssd1 vssd1 vccd1 vccd1
+ dut.pwm_a_inst_x.count_q\[8\] sky130_fd_sc_hd__dfrtp_1
X_1449_ _1036_ _1037_ dut.pwm_a_inst_y.count_q\[8\] vssd1 vssd1 vccd1 vccd1 _1038_
+ sky130_fd_sc_hd__o21a_1
X_1518_ _1101_ _1106_ vssd1 vssd1 vccd1 vccd1 _1107_ sky130_fd_sc_hd__and2_1
X_2567_ net234 net248 _0943_ vssd1 vssd1 vccd1 vccd1 _0215_ sky130_fd_sc_hd__mux2_1
X_2498_ _0838_ _0844_ net38 net44 vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_55_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_4_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2421_ _0772_ vssd1 vssd1 vccd1 vccd1 _0773_ sky130_fd_sc_hd__inv_2
X_2352_ net48 _0735_ dut.microstep_x.clk_en vssd1 vssd1 vccd1 vccd1 _0136_ sky130_fd_sc_hd__mux2_1
X_1303_ dut.ir_sensor_array.final_sensor_data\[6\] vssd1 vssd1 vccd1 vccd1 _0927_
+ sky130_fd_sc_hd__inv_2
X_2283_ _0669_ _0670_ vssd1 vssd1 vccd1 vccd1 _0671_ sky130_fd_sc_hd__and2b_1
XFILLER_64_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2619_ clknet_leaf_10_clk dut.spi.cs_low_counter_d\[5\] net69 vssd1 vssd1 vccd1 vccd1
+ dut.spi.cs_low_counter_q\[5\] sky130_fd_sc_hd__dfrtp_1
X_1998_ dut.microstep_x.ctr\[15\] dut.microstep_x.ctr\[16\] _0449_ vssd1 vssd1 vccd1
+ vccd1 _0453_ sky130_fd_sc_hd__and3_1
XFILLER_28_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1921_ _0405_ _0406_ vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__nor2_1
X_1852_ _0363_ _0364_ vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_x.count_d\[4\] sky130_fd_sc_hd__nor2_1
X_1783_ dut.pwm_a_inst_x.count_q\[10\] dut.pwm_a_inst_x.count_q\[11\] dut.pwm_a_inst_x.count_q\[9\]
+ vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__and3_1
X_2404_ dut.lcd1602.cnt_200ms\[19\] dut.lcd1602.cnt_200ms\[20\] _0762_ vssd1 vssd1
+ vccd1 vccd1 _0764_ sky130_fd_sc_hd__and3_1
X_2266_ net210 _0656_ net28 vssd1 vssd1 vccd1 vccd1 _0658_ sky130_fd_sc_hd__a21boi_1
X_2335_ _0719_ _0722_ vssd1 vssd1 vccd1 vccd1 _0723_ sky130_fd_sc_hd__nor2_1
X_2197_ net12 _0571_ vssd1 vssd1 vccd1 vccd1 _0600_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_35_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Left_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold32 dut.spi.clk_counter_q\[0\] vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 dut.lcd1602.cnt_500hz\[9\] vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 _0100_ vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 dut.spi.shift_reg_q\[7\] vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 _0104_ vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold21 dut.pid_y.y_pid.last_error\[1\] vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 dut.microstep_x.ctr\[20\] vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 dut.microstep_x.ctr\[23\] vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 dut.microstep_x.ctr\[24\] vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_51_Left_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_60_Left_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2120_ dut.spi.bit_counter_q\[1\] dut.spi.bit_counter_q\[2\] vssd1 vssd1 vccd1 vccd1
+ _0530_ sky130_fd_sc_hd__nor2_1
XFILLER_3_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2051_ dut.clkdiv_inst.counter\[9\] dut.clkdiv_inst.counter\[8\] _0480_ vssd1 vssd1
+ vccd1 vccd1 _0484_ sky130_fd_sc_hd__and3_1
X_1904_ _0910_ _0389_ vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_32_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2884_ clknet_leaf_1_clk _0005_ net53 vssd1 vssd1 vccd1 vccd1 dut.clkdiv_inst.counter\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_1835_ dut.pwm_a_inst_x.count_q\[13\] dut.pwm_a_inst_x.count_q\[15\] dut.pwm_a_inst_x.count_q\[14\]
+ dut.pwm_a_inst_x.count_q\[12\] vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__or4_1
X_1697_ _0920_ _1266_ vssd1 vssd1 vccd1 vccd1 _1267_ sky130_fd_sc_hd__nor2_1
X_1766_ _0248_ _0250_ _0283_ vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__o21ba_1
X_2249_ _0629_ _0632_ _0644_ _0647_ vssd1 vssd1 vccd1 vccd1 _0648_ sky130_fd_sc_hd__or4_1
X_2318_ net11 _0705_ vssd1 vssd1 vccd1 vccd1 _0706_ sky130_fd_sc_hd__or2_1
XFILLER_25_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput9 net9 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_46_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1620_ _1149_ _1165_ dut.pwm_a_inst_y.count_q\[13\] dut.pwm_a_inst_y.count_q\[12\]
+ vssd1 vssd1 vccd1 vccd1 _1209_ sky130_fd_sc_hd__a211o_1
X_1551_ _1103_ _1139_ _1089_ vssd1 vssd1 vccd1 vccd1 _1140_ sky130_fd_sc_hd__a21oi_1
X_1482_ _1064_ _1068_ _1070_ vssd1 vssd1 vccd1 vccd1 _1071_ sky130_fd_sc_hd__o21a_1
XFILLER_54_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2103_ net161 net20 _0520_ net252 _0521_ vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__o221a_1
XFILLER_62_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2034_ _0969_ net170 vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__nor2_1
X_2798_ clknet_leaf_8_clk _0152_ net64 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_200ms\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_2867_ clknet_leaf_3_clk _0220_ net68 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1818_ _0266_ _0270_ vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__xor2_1
X_1749_ dut.actual_duty_x\[1\] dut.actual_duty_x\[0\] vssd1 vssd1 vccd1 vccd1 _0267_
+ sky130_fd_sc_hd__or2_2
XFILLER_60_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2652_ clknet_leaf_13_clk _0123_ vssd1 vssd1 vccd1 vccd1 dut.data_in\[6\] sky130_fd_sc_hd__dfxtp_1
X_2721_ clknet_leaf_5_clk _0091_ net63 vssd1 vssd1 vccd1 vccd1 dut.microstep_y.ctr\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1534_ _1121_ _1122_ vssd1 vssd1 vccd1 vccd1 _1123_ sky130_fd_sc_hd__nor2_1
X_1465_ net40 dut.actual_duty_y\[7\] vssd1 vssd1 vccd1 vccd1 _1054_ sky130_fd_sc_hd__or2_1
X_1603_ dut.actual_duty_y\[0\] _1122_ vssd1 vssd1 vccd1 vccd1 _1192_ sky130_fd_sc_hd__nor2_1
X_2583_ dut.ir_sensor_array.final_sensor_data\[20\] _0880_ dut.ir_sensor_array.final_sensor_data\[19\]
+ vssd1 vssd1 vccd1 vccd1 _0881_ sky130_fd_sc_hd__o21ba_1
X_1396_ _0999_ _1000_ _0991_ vssd1 vssd1 vccd1 vccd1 dut.spi.cs_low_counter_d\[5\]
+ sky130_fd_sc_hd__o21a_1
X_2017_ dut.microstep_x.ctr\[23\] _0463_ net239 vssd1 vssd1 vccd1 vccd1 _0464_ sky130_fd_sc_hd__a21oi_1
XFILLER_50_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xteam_02_98 vssd1 vssd1 vccd1 vccd1 team_02_98/HI gpio_out[0] sky130_fd_sc_hd__conb_1
Xhold140 dut.clkdiv_inst.counter\[8\] vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 dut.pwm_a_inst_x.count_q\[7\] vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 dut.microstep_x.ctr\[11\] vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2635_ clknet_leaf_13_clk net243 net82 vssd1 vssd1 vccd1 vccd1 dut.spi.shift_reg_q\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_2704_ clknet_leaf_21_clk dut.pwm_a_inst_x.count_d\[7\] net76 vssd1 vssd1 vccd1 vccd1
+ dut.pwm_a_inst_x.count_q\[7\] sky130_fd_sc_hd__dfrtp_4
X_1448_ dut.pwm_a_inst_y.count_q\[7\] dut.pwm_a_inst_y.count_q\[6\] vssd1 vssd1 vccd1
+ vccd1 _1037_ sky130_fd_sc_hd__or2_1
X_1517_ _1099_ _1100_ vssd1 vssd1 vccd1 vccd1 _1106_ sky130_fd_sc_hd__or2_1
X_2566_ net234 dut.ir_sensor_array.final_sensor_data\[31\] net34 vssd1 vssd1 vccd1
+ vccd1 _0214_ sky130_fd_sc_hd__mux2_1
X_2497_ _0807_ _0813_ _0819_ _0833_ net44 vssd1 vssd1 vccd1 vccd1 _0844_ sky130_fd_sc_hd__o221a_1
X_1379_ _0908_ _0988_ _0989_ vssd1 vssd1 vccd1 vccd1 dut.spi.clk_counter_d\[5\] sky130_fd_sc_hd__a21oi_1
XFILLER_55_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_53_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2420_ _0507_ _0771_ _0770_ vssd1 vssd1 vccd1 vccd1 _0772_ sky130_fd_sc_hd__a21bo_1
X_1302_ dut.ir_sensor_array.final_sensor_data\[33\] vssd1 vssd1 vccd1 vccd1 _0926_
+ sky130_fd_sc_hd__inv_2
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2351_ _0734_ _0714_ _0719_ vssd1 vssd1 vccd1 vccd1 _0735_ sky130_fd_sc_hd__mux2_1
X_2282_ dut.pid_x.x_pid.last_error\[2\] _0925_ _0509_ vssd1 vssd1 vccd1 vccd1 _0670_
+ sky130_fd_sc_hd__o21a_1
XFILLER_64_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1997_ net309 _0449_ _0452_ vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__o21a_1
XFILLER_20_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2618_ clknet_leaf_10_clk dut.spi.cs_low_counter_d\[4\] net81 vssd1 vssd1 vccd1 vccd1
+ dut.spi.cs_low_counter_q\[4\] sky130_fd_sc_hd__dfrtp_1
X_2549_ dut.ir_sensor_array.final_sensor_data\[14\] dut.ir_sensor_array.final_sensor_data\[15\]
+ _0943_ vssd1 vssd1 vccd1 vccd1 _0197_ sky130_fd_sc_hd__mux2_1
XFILLER_18_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1920_ dut.microstep_y.ctr\[13\] _0402_ net249 vssd1 vssd1 vccd1 vccd1 _0406_ sky130_fd_sc_hd__a21oi_1
X_1851_ dut.pwm_a_inst_x.count_q\[4\] _0361_ net27 vssd1 vssd1 vccd1 vccd1 _0364_
+ sky130_fd_sc_hd__o21ai_1
X_2403_ net198 _0762_ vssd1 vssd1 vccd1 vccd1 _0159_ sky130_fd_sc_hd__xor2_1
XANTENNA_clkbuf_leaf_3_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1782_ _0298_ _0299_ vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__and2_1
X_2196_ _0547_ _0553_ vssd1 vssd1 vccd1 vccd1 _0599_ sky130_fd_sc_hd__nand2_1
X_2265_ net28 _0655_ _0657_ vssd1 vssd1 vccd1 vccd1 _0127_ sky130_fd_sc_hd__and3_1
X_2334_ _0698_ _0699_ _0721_ vssd1 vssd1 vccd1 vccd1 _0722_ sky130_fd_sc_hd__a21o_2
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold22 dut.microstep_y.ctr\[5\] vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 dut.microstep_x.ctr\[5\] vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 dut.lcd1602.cnt_200ms\[12\] vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 _0107_ vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 dut.lcd1602.cnt_500hz\[14\] vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 dut.microstep_y.ctr\[29\] vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 dut.lcd1602.cnt_200ms\[2\] vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 dut.microstep_y.ctr\[23\] vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_26_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold88 dut.pwm_a_inst_x.count_q\[1\] vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_43_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2050_ dut.clkdiv_inst.counter\[8\] _0480_ dut.clkdiv_inst.counter\[9\] vssd1 vssd1
+ vccd1 vccd1 _0483_ sky130_fd_sc_hd__a21oi_1
XFILLER_19_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1903_ _0388_ _0389_ _0395_ vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__and3_1
X_2883_ clknet_leaf_1_clk _0004_ net53 vssd1 vssd1 vccd1 vccd1 dut.clkdiv_inst.counter\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_1765_ _0261_ _0282_ _0251_ vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__a21oi_1
X_1834_ dut.pwm_a_inst_x.count_q\[7\] dut.pwm_a_inst_x.count_q\[6\] dut.pwm_a_inst_x.count_q\[10\]
+ dut.pwm_a_inst_x.count_q\[11\] dut.pwm_a_inst_x.count_q\[8\] vssd1 vssd1 vccd1 vccd1
+ _0352_ sky130_fd_sc_hd__o2111a_1
X_1696_ _1261_ _1264_ vssd1 vssd1 vccd1 vccd1 _1266_ sky130_fd_sc_hd__xor2_1
XFILLER_57_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2248_ _0598_ _0606_ _0613_ vssd1 vssd1 vccd1 vccd1 _0647_ sky130_fd_sc_hd__or3_1
X_2179_ _0577_ _0580_ vssd1 vssd1 vccd1 vccd1 _0582_ sky130_fd_sc_hd__or2_2
X_2317_ _0701_ _0704_ vssd1 vssd1 vccd1 vccd1 _0705_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_23_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_2_0__f_clk_X clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1550_ _1115_ _1138_ _1105_ vssd1 vssd1 vccd1 vccd1 _1139_ sky130_fd_sc_hd__a21o_1
X_1481_ _1044_ _1067_ _1069_ vssd1 vssd1 vccd1 vccd1 _1070_ sky130_fd_sc_hd__o21ai_1
X_2102_ dut.data_in\[1\] _0515_ vssd1 vssd1 vccd1 vccd1 _0521_ sky130_fd_sc_hd__or2_1
XFILLER_11_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2033_ dut.clkdiv_inst.counter\[1\] dut.clkdiv_inst.counter\[0\] net169 vssd1 vssd1
+ vccd1 vccd1 _0473_ sky130_fd_sc_hd__a21oi_1
X_2797_ clknet_leaf_7_clk _0151_ net64 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_200ms\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_2866_ clknet_leaf_3_clk _0219_ net68 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[37\]
+ sky130_fd_sc_hd__dfrtp_1
X_1748_ dut.actual_duty_x\[1\] _0256_ vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__xnor2_1
X_1817_ dut.pwm_a_inst_x.count_q\[2\] _0331_ _0334_ vssd1 vssd1 vccd1 vccd1 _0335_
+ sky130_fd_sc_hd__a21o_1
X_1679_ _1246_ _1248_ vssd1 vssd1 vccd1 vccd1 _1249_ sky130_fd_sc_hd__nand2_1
XFILLER_45_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2651_ clknet_leaf_12_clk _0122_ vssd1 vssd1 vccd1 vccd1 dut.data_in\[5\] sky130_fd_sc_hd__dfxtp_1
X_1602_ _0913_ _1189_ _1190_ _1187_ vssd1 vssd1 vccd1 vccd1 _1191_ sky130_fd_sc_hd__o211a_1
X_2720_ clknet_leaf_1_clk _0090_ net55 vssd1 vssd1 vccd1 vccd1 dut.microstep_y.ctr\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2582_ dut.ir_sensor_array.final_sensor_data\[22\] _0879_ dut.ir_sensor_array.final_sensor_data\[21\]
+ vssd1 vssd1 vccd1 vccd1 _0880_ sky130_fd_sc_hd__o21ba_1
X_1395_ dut.spi.cs_low_counter_q\[5\] _0998_ vssd1 vssd1 vccd1 vccd1 _1000_ sky130_fd_sc_hd__and2_1
X_1464_ net40 _1046_ vssd1 vssd1 vccd1 vccd1 _1053_ sky130_fd_sc_hd__nor2_1
X_1533_ net41 dut.actual_duty_y\[1\] vssd1 vssd1 vccd1 vccd1 _1122_ sky130_fd_sc_hd__nor2_1
XFILLER_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2016_ net195 _0463_ vssd1 vssd1 vccd1 vccd1 _0051_ sky130_fd_sc_hd__xor2_1
Xteam_02_88 vssd1 vssd1 vccd1 vccd1 team_02_88/HI gpio_oeb[3] sky130_fd_sc_hd__conb_1
Xteam_02_99 vssd1 vssd1 vccd1 vccd1 team_02_99/HI gpio_out[1] sky130_fd_sc_hd__conb_1
XFILLER_50_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold130 dut.spi.bit_counter_q\[2\] vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 dut.pwm_a_inst_y.count_q\[17\] vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 dut.microstep_y.ctr\[11\] vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 dut.ir_sensor_array.final_sensor_data\[25\] vssd1 vssd1 vccd1 vccd1 net315
+ sky130_fd_sc_hd__dlygate4sd3_1
X_2849_ clknet_leaf_2_clk _0202_ net54 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_2_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_5_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_21_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_1_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_12_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_32_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2634_ clknet_leaf_13_clk net220 net79 vssd1 vssd1 vccd1 vccd1 dut.spi.shift_reg_q\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_1516_ _1103_ _1104_ vssd1 vssd1 vccd1 vccd1 _1105_ sky130_fd_sc_hd__nand2_1
X_2565_ dut.ir_sensor_array.final_sensor_data\[31\] dut.ir_sensor_array.final_sensor_data\[30\]
+ net33 vssd1 vssd1 vccd1 vccd1 _0213_ sky130_fd_sc_hd__mux2_1
X_2703_ clknet_leaf_20_clk dut.pwm_a_inst_x.count_d\[6\] net77 vssd1 vssd1 vccd1 vccd1
+ dut.pwm_a_inst_x.count_q\[6\] sky130_fd_sc_hd__dfrtp_2
X_1378_ dut.spi.clk_counter_q\[5\] dut.spi.clk_counter_q\[4\] _0987_ _0977_ vssd1
+ vssd1 vccd1 vccd1 _0989_ sky130_fd_sc_hd__a31o_1
X_1447_ dut.pwm_a_inst_y.count_q\[5\] dut.pwm_a_inst_y.count_q\[4\] vssd1 vssd1 vccd1
+ vccd1 _1036_ sky130_fd_sc_hd__or2_2
X_2496_ _0842_ _0843_ net39 net44 vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout80 net87 vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_1_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1301_ dut.pid_x.x_pid.last_error\[3\] vssd1 vssd1 vccd1 vccd1 _0925_ sky130_fd_sc_hd__inv_2
X_2350_ _0677_ _0682_ _0722_ vssd1 vssd1 vccd1 vccd1 _0734_ sky130_fd_sc_hd__mux2_1
X_2281_ _0512_ _0668_ vssd1 vssd1 vccd1 vccd1 _0669_ sky130_fd_sc_hd__xnor2_1
XFILLER_64_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1996_ _0035_ _0451_ vssd1 vssd1 vccd1 vccd1 _0452_ sky130_fd_sc_hd__nor2_1
X_2617_ clknet_leaf_14_clk dut.spi.cs_low_counter_d\[3\] net81 vssd1 vssd1 vccd1 vccd1
+ dut.spi.cs_low_counter_q\[3\] sky130_fd_sc_hd__dfrtp_1
X_2548_ dut.ir_sensor_array.final_sensor_data\[14\] net308 net31 vssd1 vssd1 vccd1
+ vccd1 _0196_ sky130_fd_sc_hd__mux2_1
X_2479_ _0786_ _0819_ _0821_ _0802_ _0829_ vssd1 vssd1 vccd1 vccd1 _0831_ sky130_fd_sc_hd__a221o_1
XFILLER_28_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload0 clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload0/X sky130_fd_sc_hd__clkbuf_8
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1850_ dut.pwm_a_inst_x.count_q\[4\] _0361_ vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__and2_1
X_1781_ dut.pwm_a_inst_x.count_q\[12\] _0297_ vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__nand2_1
X_2402_ _0762_ _0763_ vssd1 vssd1 vccd1 vccd1 _0158_ sky130_fd_sc_hd__nor2_1
X_2333_ _1245_ _1247_ _0694_ vssd1 vssd1 vccd1 vccd1 _0721_ sky130_fd_sc_hd__mux2_1
X_2195_ _0571_ _0588_ _0597_ _0581_ vssd1 vssd1 vccd1 vccd1 _0598_ sky130_fd_sc_hd__a22o_1
X_2264_ _0656_ vssd1 vssd1 vccd1 vccd1 _0657_ sky130_fd_sc_hd__inv_2
XFILLER_52_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1979_ _0911_ _0433_ _0441_ vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__a21oi_1
Xhold56 dut.lcd1602.cnt_200ms\[17\] vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 dut.spi.clk_counter_q\[2\] vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 _0387_ vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 dut.microstep_x.ctr\[29\] vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 _0431_ vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_20_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold78 dut.lcd1602.cnt_200ms\[18\] vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 dut.spi.shift_reg_q\[5\] vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_26_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold89 dut.pwm_a_inst_x.count_d\[1\] vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_19_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1902_ _0948_ _0392_ _0394_ vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__or3_1
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2882_ clknet_leaf_1_clk _0003_ net53 vssd1 vssd1 vccd1 vccd1 dut.clkdiv_inst.counter\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_1833_ _0291_ _0348_ _0349_ _0347_ vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__a22o_1
X_1764_ _0280_ _0281_ _0263_ vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__o21ai_1
X_2316_ net48 _0700_ net47 vssd1 vssd1 vccd1 vccd1 _0704_ sky130_fd_sc_hd__a21oi_1
X_1695_ _1261_ _1264_ vssd1 vssd1 vccd1 vccd1 _1265_ sky130_fd_sc_hd__and2b_1
X_2247_ net158 net19 net79 _0646_ vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__o211a_1
X_2178_ _0577_ _0580_ vssd1 vssd1 vccd1 vccd1 _0581_ sky130_fd_sc_hd__nor2_1
XFILLER_25_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_2_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1480_ _1064_ _1068_ vssd1 vssd1 vccd1 vccd1 _1069_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2101_ dut.data_in\[0\] dut.lcd1602.out_valid _0513_ _0519_ net161 vssd1 vssd1 vccd1
+ vccd1 _0100_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2032_ net182 net155 vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__xor2_1
XFILLER_50_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2865_ clknet_leaf_3_clk _0218_ net68 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_22_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2796_ clknet_leaf_9_clk _0150_ net65 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_200ms\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1678_ net46 net45 vssd1 vssd1 vccd1 vccd1 _1248_ sky130_fd_sc_hd__or2_1
X_1747_ _0258_ _0264_ vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__nand2_1
X_1816_ dut.pwm_a_inst_x.count_q\[2\] _0331_ _0332_ dut.pwm_a_inst_x.count_q\[1\]
+ _0333_ vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_39_Left_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Left_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xteam_02_150 vssd1 vssd1 vccd1 vccd1 gpio_out[3] team_02_150/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_8_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_57_Left_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2650_ clknet_leaf_12_clk _0121_ vssd1 vssd1 vccd1 vccd1 dut.data_in\[4\] sky130_fd_sc_hd__dfxtp_1
X_1601_ _0914_ net42 _1188_ dut.pwm_a_inst_y.count_q\[1\] vssd1 vssd1 vccd1 vccd1
+ _1190_ sky130_fd_sc_hd__o22a_1
X_1532_ net41 dut.actual_duty_y\[1\] vssd1 vssd1 vccd1 vccd1 _1121_ sky130_fd_sc_hd__and2_1
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2581_ dut.ir_sensor_array.final_sensor_data\[8\] _0878_ dut.ir_sensor_array.final_sensor_data\[23\]
+ vssd1 vssd1 vccd1 vccd1 _0879_ sky130_fd_sc_hd__o21ba_1
X_1394_ dut.spi.cs_low_counter_q\[5\] _0998_ vssd1 vssd1 vccd1 vccd1 _0999_ sky130_fd_sc_hd__nor2_1
X_1463_ net40 dut.actual_duty_y\[7\] dut.actual_duty_y\[5\] vssd1 vssd1 vccd1 vccd1
+ _1052_ sky130_fd_sc_hd__a21o_1
XFILLER_27_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2015_ _0462_ _0463_ vssd1 vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__nor2_1
X_2848_ clknet_leaf_2_clk _0201_ net54 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[19\]
+ sky130_fd_sc_hd__dfrtp_1
Xteam_02_89 vssd1 vssd1 vccd1 vccd1 team_02_89/HI gpio_oeb[4] sky130_fd_sc_hd__conb_1
XFILLER_12_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold142 dut.spi.bit_counter_q\[3\] vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 dut.microstep_y.ctr\[8\] vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 dut.ball_pos_y\[0\] vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 dut.pwm_a_inst_x.count_q\[15\] vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__dlygate4sd3_1
X_2779_ clknet_leaf_29_clk _0051_ net50 vssd1 vssd1 vccd1 vccd1 dut.microstep_x.ctr\[23\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold120 dut.microstep_x.ctr\[6\] vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout59_A net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2702_ clknet_leaf_20_clk dut.pwm_a_inst_x.count_d\[5\] net77 vssd1 vssd1 vccd1 vccd1
+ dut.pwm_a_inst_x.count_q\[5\] sky130_fd_sc_hd__dfrtp_1
X_2633_ clknet_leaf_13_clk net217 net80 vssd1 vssd1 vccd1 vccd1 dut.spi.shift_reg_q\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1515_ _1091_ _1102_ vssd1 vssd1 vccd1 vccd1 _1104_ sky130_fd_sc_hd__nand2_1
X_2495_ _0821_ _0833_ _0834_ _0801_ dut.microstep_y.clk_en vssd1 vssd1 vccd1 vccd1
+ _0843_ sky130_fd_sc_hd__o221a_1
X_2564_ dut.ir_sensor_array.final_sensor_data\[30\] net320 net33 vssd1 vssd1 vccd1
+ vccd1 _0212_ sky130_fd_sc_hd__mux2_1
X_1377_ dut.spi.clk_counter_q\[4\] _0987_ _0988_ _0983_ vssd1 vssd1 vccd1 vccd1 dut.spi.clk_counter_d\[4\]
+ sky130_fd_sc_hd__o211a_1
X_1446_ net218 _1033_ _1035_ vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__o21a_1
XFILLER_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout81 net83 vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__buf_2
Xfanout70 net71 vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_24_Left_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1300_ dut.pid_y.y_pid.last_error\[3\] vssd1 vssd1 vccd1 vccd1 _0924_ sky130_fd_sc_hd__inv_2
XFILLER_1_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2280_ _0664_ _0667_ _0666_ vssd1 vssd1 vccd1 vccd1 _0668_ sky130_fd_sc_hd__o21ba_1
XFILLER_52_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2616_ clknet_leaf_14_clk dut.spi.cs_low_counter_d\[2\] net81 vssd1 vssd1 vccd1 vccd1
+ dut.spi.cs_low_counter_q\[2\] sky130_fd_sc_hd__dfrtp_1
X_1995_ dut.microstep_x.ctr\[15\] _0449_ vssd1 vssd1 vccd1 vccd1 _0451_ sky130_fd_sc_hd__and2_1
XFILLER_20_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1429_ dut.lcd1602.cnt_500hz\[7\] dut.lcd1602.cnt_500hz\[8\] _1021_ vssd1 vssd1 vccd1
+ vccd1 _1025_ sky130_fd_sc_hd__and3_1
X_2478_ _1048_ _0814_ net37 vssd1 vssd1 vccd1 vccd1 _0830_ sky130_fd_sc_hd__a21oi_1
X_2547_ net308 dut.ir_sensor_array.final_sensor_data\[12\] net31 vssd1 vssd1 vccd1
+ vccd1 _0195_ sky130_fd_sc_hd__mux2_1
XFILLER_55_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload1 clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload1/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_21_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1780_ dut.pwm_a_inst_x.count_q\[12\] _0297_ vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__or2_1
X_2401_ net230 _0760_ vssd1 vssd1 vccd1 vccd1 _0763_ sky130_fd_sc_hd__nor2_1
XFILLER_34_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2332_ _0719_ vssd1 vssd1 vccd1 vccd1 _0720_ sky130_fd_sc_hd__inv_2
X_2194_ _0595_ _0596_ vssd1 vssd1 vccd1 vccd1 _0597_ sky130_fd_sc_hd__nand2_1
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2263_ dut.ir_sensor_array.bit_count\[1\] _0653_ vssd1 vssd1 vccd1 vccd1 _0656_ sky130_fd_sc_hd__and2_1
XFILLER_1_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1978_ net15 _0440_ vssd1 vssd1 vccd1 vccd1 _0441_ sky130_fd_sc_hd__or2_1
Xhold46 dut.lcd1602.cnt_200ms\[19\] vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 _0761_ vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 dut.spi.cs_low_counter_q\[0\] vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 _0105_ vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 dut.data_in\[5\] vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 dut.clkdiv_inst.counter\[16\] vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold13 dut.pid_x.x_pid.last_error\[1\] vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1901_ _0951_ _0953_ _0954_ _0393_ vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__or4_1
XFILLER_34_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2881_ clknet_leaf_1_clk _0018_ net56 vssd1 vssd1 vccd1 vccd1 dut.clkdiv_inst.counter\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_1832_ dut.pwm_a_inst_x.count_q\[13\] _0298_ dut.pwm_a_inst_x.count_q\[14\] vssd1
+ vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__a21oi_1
X_1694_ net46 dut.actual_duty_x\[5\] _1263_ vssd1 vssd1 vccd1 vccd1 _1264_ sky130_fd_sc_hd__a21bo_1
X_1763_ _0260_ _0272_ vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__nor2_1
X_2246_ _0606_ _0629_ _0645_ _0643_ vssd1 vssd1 vccd1 vccd1 _0646_ sky130_fd_sc_hd__or4b_1
XPHY_EDGE_ROW_27_Left_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2315_ net45 _0702_ vssd1 vssd1 vccd1 vccd1 _0703_ sky130_fd_sc_hd__nor2_1
X_2177_ dut.lcd1602.currentState\[5\] _0579_ vssd1 vssd1 vccd1 vccd1 _0580_ sky130_fd_sc_hd__nor2_1
XFILLER_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Left_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2100_ _0515_ net20 vssd1 vssd1 vccd1 vccd1 _0520_ sky130_fd_sc_hd__nand2_2
XFILLER_62_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2031_ net186 _0471_ _0472_ vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__a21o_1
X_2795_ clknet_leaf_9_clk _0149_ net65 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_200ms\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_2864_ clknet_leaf_12_clk _0217_ net68 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[35\]
+ sky130_fd_sc_hd__dfrtp_1
X_1815_ dut.pwm_a_inst_x.count_q\[1\] dut.actual_duty_x\[1\] _0922_ dut.pwm_a_inst_x.count_q\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__a211o_1
X_1677_ net46 net45 vssd1 vssd1 vccd1 vccd1 _1247_ sky130_fd_sc_hd__nor2_1
X_1746_ _0253_ _0257_ vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__nand2_1
X_2229_ _0576_ _0596_ vssd1 vssd1 vccd1 vccd1 _0632_ sky130_fd_sc_hd__nor2_1
XANTENNA__2870__RESET_B net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xteam_02_140 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] team_02_140/LO sky130_fd_sc_hd__conb_1
Xteam_02_151 vssd1 vssd1 vccd1 vccd1 gpio_out[4] team_02_151/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_42_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1531_ net39 _1110_ vssd1 vssd1 vccd1 vccd1 _1120_ sky130_fd_sc_hd__xnor2_1
X_1462_ dut.actual_duty_y\[6\] _1049_ _1047_ vssd1 vssd1 vccd1 vccd1 _1051_ sky130_fd_sc_hd__o21a_1
X_1600_ _1188_ vssd1 vssd1 vccd1 vccd1 _1189_ sky130_fd_sc_hd__inv_2
X_2580_ dut.ir_sensor_array.final_sensor_data\[10\] _0877_ dut.ir_sensor_array.final_sensor_data\[9\]
+ vssd1 vssd1 vccd1 vccd1 _0878_ sky130_fd_sc_hd__o21ba_1
X_1393_ _0991_ _0997_ _0998_ vssd1 vssd1 vccd1 vccd1 dut.spi.cs_low_counter_d\[4\]
+ sky130_fd_sc_hd__and3_1
X_2014_ dut.microstep_x.ctr\[22\] _0461_ vssd1 vssd1 vccd1 vccd1 _0463_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_2_1__f_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2847_ clknet_leaf_2_clk _0200_ net59 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[18\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold110 dut.microstep_x.ctr\[14\] vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__dlygate4sd3_1
X_2778_ clknet_leaf_29_clk _0050_ net50 vssd1 vssd1 vccd1 vccd1 dut.microstep_x.ctr\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold121 dut.microstep_y.ctr\[6\] vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_1_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold143 dut.clkdiv_inst.counter\[6\] vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 dut.microstep_x.ctr\[8\] vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 dut.actual_duty_x\[3\] vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__dlygate4sd3_1
X_1729_ _0240_ _0244_ _0246_ vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__o21ba_1
Xhold165 dut.ir_sensor_array.final_sensor_data\[23\] vssd1 vssd1 vccd1 vccd1 net317
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2632_ clknet_leaf_13_clk net223 net80 vssd1 vssd1 vccd1 vccd1 dut.spi.shift_reg_q\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_2701_ clknet_leaf_20_clk dut.pwm_a_inst_x.count_d\[4\] net77 vssd1 vssd1 vccd1 vccd1
+ dut.pwm_a_inst_x.count_q\[4\] sky130_fd_sc_hd__dfrtp_2
X_1445_ net218 _1033_ _1019_ vssd1 vssd1 vccd1 vccd1 _1035_ sky130_fd_sc_hd__a21oi_1
X_1514_ _1091_ _1102_ vssd1 vssd1 vccd1 vccd1 _1103_ sky130_fd_sc_hd__or2_1
X_2494_ _0811_ _0812_ _0803_ vssd1 vssd1 vccd1 vccd1 _0842_ sky130_fd_sc_hd__o21ai_1
X_2563_ net320 dut.ir_sensor_array.final_sensor_data\[28\] net33 vssd1 vssd1 vccd1
+ vccd1 _0211_ sky130_fd_sc_hd__mux2_1
XFILLER_4_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1376_ dut.spi.clk_counter_q\[4\] _0987_ vssd1 vssd1 vccd1 vccd1 _0988_ sky130_fd_sc_hd__nand2_1
XFILLER_55_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout71_A net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout82 net83 vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__clkbuf_4
Xfanout71 net72 vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__buf_2
XFILLER_6_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout60 net61 vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_4
XFILLER_37_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1994_ _0449_ _0450_ vssd1 vssd1 vccd1 vccd1 _0041_ sky130_fd_sc_hd__nor2_1
XFILLER_20_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2615_ clknet_leaf_10_clk net232 net81 vssd1 vssd1 vccd1 vccd1 dut.spi.cs_low_counter_q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1428_ dut.lcd1602.cnt_500hz\[6\] dut.lcd1602.cnt_500hz\[7\] _0934_ dut.lcd1602.cnt_500hz\[8\]
+ vssd1 vssd1 vccd1 vccd1 _1024_ sky130_fd_sc_hd__a31o_1
X_2477_ _0802_ _0821_ _0823_ _0793_ _0828_ vssd1 vssd1 vccd1 vccd1 _0829_ sky130_fd_sc_hd__o221a_1
X_2546_ dut.ir_sensor_array.final_sensor_data\[12\] dut.ir_sensor_array.final_sensor_data\[11\]
+ net31 vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__mux2_1
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1359_ dut.spi.state_q\[0\] _0975_ vssd1 vssd1 vccd1 vccd1 _0976_ sky130_fd_sc_hd__and2_1
XFILLER_28_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload2 clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload2/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_21_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2400_ dut.lcd1602.cnt_200ms\[18\] _0760_ vssd1 vssd1 vccd1 vccd1 _0762_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_12_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2262_ dut.ir_sensor_array.bit_count\[1\] _0653_ vssd1 vssd1 vccd1 vccd1 _0655_ sky130_fd_sc_hd__or2_1
X_2331_ _1246_ _0706_ _0716_ _0718_ _0703_ vssd1 vssd1 vccd1 vccd1 _0719_ sky130_fd_sc_hd__a41o_2
XFILLER_52_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2193_ net12 _0570_ _0587_ vssd1 vssd1 vccd1 vccd1 _0596_ sky130_fd_sc_hd__or3_1
XFILLER_1_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1977_ _0911_ _0433_ vssd1 vssd1 vccd1 vccd1 _0440_ sky130_fd_sc_hd__nor2_1
X_2529_ dut.ball_pos_y\[1\] net28 _0866_ _0867_ vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__a22o_1
Xhold25 dut.spi.shift_reg_q\[8\] vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 dut.microstep_y.ctr\[4\] vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 dut.ir_sensor_array.bit_count\[2\] vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 dut.ir_sensor_array.bit_count\[0\] vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 dut.pwm_a_inst_x.count_q\[12\] vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 dut.microstep_x.ctr\[1\] vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1900_ dut.microstep_y.ctr\[12\] dut.microstep_y.ctr\[14\] dut.microstep_y.ctr\[17\]
+ dut.microstep_y.ctr\[13\] vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__or4bb_1
X_2880_ clknet_leaf_1_clk _0017_ net53 vssd1 vssd1 vccd1 vccd1 dut.clkdiv_inst.counter\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_1831_ _0292_ _0300_ _0348_ _0291_ vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__o22a_1
X_1693_ net48 _1262_ vssd1 vssd1 vccd1 vccd1 _1263_ sky130_fd_sc_hd__nand2_1
X_1762_ _0277_ _0279_ vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__nor2_1
X_2245_ _0589_ _0593_ _0616_ _0644_ vssd1 vssd1 vccd1 vccd1 _0645_ sky130_fd_sc_hd__or4_1
X_2176_ _0563_ _0578_ dut.lcd1602.currentState\[4\] vssd1 vssd1 vccd1 vccd1 _0579_
+ sky130_fd_sc_hd__a21oi_1
X_2314_ net46 _0701_ vssd1 vssd1 vccd1 vccd1 _0702_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_31_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2030_ dut.microstep_x.ctr\[29\] dut.microstep_x.ctr\[28\] _0469_ vssd1 vssd1 vccd1
+ vccd1 _0472_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_45_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2794_ clknet_leaf_8_clk _0148_ net66 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_200ms\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_2863_ clknet_leaf_3_clk _0216_ net71 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1745_ _0261_ _0262_ vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__and2_1
X_1814_ _0267_ _0268_ vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__nand2_1
X_1676_ net46 net45 vssd1 vssd1 vccd1 vccd1 _1246_ sky130_fd_sc_hd__nand2_1
XFILLER_7_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2228_ _0630_ vssd1 vssd1 vccd1 vccd1 _0631_ sky130_fd_sc_hd__inv_2
X_2159_ _0541_ _0548_ _0561_ dut.lcd1602.currentState\[3\] vssd1 vssd1 vccd1 vccd1
+ _0562_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_41_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_51_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xteam_02_152 vssd1 vssd1 vccd1 vccd1 gpio_out[5] team_02_152/LO sky130_fd_sc_hd__conb_1
Xteam_02_141 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] team_02_141/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_59_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xteam_02_130 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] team_02_130/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_8_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_24_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1392_ dut.spi.cs_low_counter_q\[4\] _0996_ vssd1 vssd1 vccd1 vccd1 _0998_ sky130_fd_sc_hd__nand2_1
X_1530_ _1114_ _1118_ vssd1 vssd1 vccd1 vccd1 _1119_ sky130_fd_sc_hd__nor2_1
X_1461_ _1049_ vssd1 vssd1 vccd1 vccd1 _1050_ sky130_fd_sc_hd__inv_2
X_2013_ net275 _0461_ vssd1 vssd1 vccd1 vccd1 _0462_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_15_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold144 dut.lcd1602.cnt_200ms\[4\] vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__dlygate4sd3_1
Xhold100 dut.spi.shift_reg_q\[1\] vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 dut.ir_sensor_array.final_sensor_data\[35\] vssd1 vssd1 vccd1 vccd1 net274
+ sky130_fd_sc_hd__dlygate4sd3_1
X_2846_ clknet_leaf_2_clk _0199_ net59 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_2777_ clknet_leaf_29_clk _0049_ net50 vssd1 vssd1 vccd1 vccd1 dut.microstep_x.ctr\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold111 dut.microstep_x.ctr\[18\] vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 dut.microstep_x.ctr\[25\] vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__dlygate4sd3_1
X_1728_ _0922_ _0245_ vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__nor2_1
XFILLER_58_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1659_ dut.pwm_a_inst_y.count_q\[12\] _1234_ net22 vssd1 vssd1 vccd1 vccd1 _1235_
+ sky130_fd_sc_hd__o21ai_1
Xhold166 dut.pwm_a_inst_y.count_q\[1\] vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 dut.ir_sensor_array.final_sensor_data\[1\] vssd1 vssd1 vccd1 vccd1 net307
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_64_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2631_ clknet_leaf_13_clk net247 net82 vssd1 vssd1 vccd1 vccd1 dut.spi.shift_reg_q\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2562_ dut.ir_sensor_array.final_sensor_data\[28\] dut.ir_sensor_array.final_sensor_data\[27\]
+ net33 vssd1 vssd1 vccd1 vccd1 _0210_ sky130_fd_sc_hd__mux2_1
X_2700_ clknet_leaf_20_clk dut.pwm_a_inst_x.count_d\[3\] net77 vssd1 vssd1 vccd1 vccd1
+ dut.pwm_a_inst_x.count_q\[3\] sky130_fd_sc_hd__dfrtp_1
X_1375_ _0987_ _0976_ _0986_ vssd1 vssd1 vccd1 vccd1 dut.spi.clk_counter_d\[3\] sky130_fd_sc_hd__and3b_1
X_1444_ net202 _1032_ _1034_ vssd1 vssd1 vccd1 vccd1 _0024_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_4_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1513_ _1093_ _1098_ _1101_ vssd1 vssd1 vccd1 vccd1 _1102_ sky130_fd_sc_hd__o21a_1
X_2493_ _0840_ _0841_ dut.actual_duty_y\[3\] net44 vssd1 vssd1 vccd1 vccd1 _0171_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2829_ clknet_leaf_25_clk _0182_ net73 vssd1 vssd1 vccd1 vccd1 dut.ball_pos_y\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_46_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout83 net87 vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__clkbuf_2
Xfanout61 net72 vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_2
Xfanout50 net52 vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_4
Xfanout72 dut.clkdiv_inst.reset_n vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__clkbuf_2
XFILLER_64_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1993_ dut.microstep_x.ctr\[13\] _0446_ net262 vssd1 vssd1 vccd1 vccd1 _0450_ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_0_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2614_ clknet_leaf_10_clk dut.spi.cs_low_counter_d\[0\] net69 vssd1 vssd1 vccd1 vccd1
+ dut.spi.cs_low_counter_q\[0\] sky130_fd_sc_hd__dfrtp_2
Xclkload20 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 clkload20/Y sky130_fd_sc_hd__inv_8
X_2545_ dut.ir_sensor_array.final_sensor_data\[11\] dut.ir_sensor_array.final_sensor_data\[10\]
+ net31 vssd1 vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__mux2_1
X_1358_ dut.spi.state_q\[2\] dut.spi.state_q\[1\] vssd1 vssd1 vccd1 vccd1 _0975_ sky130_fd_sc_hd__nor2_1
X_1427_ _1018_ _1022_ _1023_ vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__and3_1
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2476_ _0793_ _0823_ _0826_ _0827_ vssd1 vssd1 vccd1 vccd1 _0828_ sky130_fd_sc_hd__a22o_1
X_1289_ dut.pwm_a_inst_y.count_q\[1\] vssd1 vssd1 vccd1 vccd1 _0913_ sky130_fd_sc_hd__inv_2
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload3 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 clkload3/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_21_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_2_3__f_clk_X clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2192_ _0554_ _0592_ vssd1 vssd1 vccd1 vccd1 _0595_ sky130_fd_sc_hd__or2_1
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2261_ net199 net34 net28 _0654_ vssd1 vssd1 vccd1 vccd1 _0126_ sky130_fd_sc_hd__o211a_1
X_2330_ _0702_ _0717_ vssd1 vssd1 vccd1 vccd1 _0718_ sky130_fd_sc_hd__or2_1
XFILLER_33_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1976_ _0432_ _0433_ _0439_ vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__and3_1
X_2528_ _0851_ _0863_ net29 vssd1 vssd1 vccd1 vccd1 _0867_ sky130_fd_sc_hd__and3_1
Xhold37 dut.lcd1602.cnt_500hz\[0\] vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 dut.lcd1602.cnt_200ms\[15\] vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold48 dut.lcd1602.cnt_500hz\[10\] vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 _0108_ vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__dlygate4sd3_1
X_2459_ _0809_ _0810_ vssd1 vssd1 vccd1 vccd1 _0811_ sky130_fd_sc_hd__and2_1
Xhold15 dut.microstep_x.ctr\[4\] vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1830_ dut.pwm_a_inst_x.count_q\[13\] _0298_ vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__xnor2_1
X_1761_ _0260_ _0278_ vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__xor2_1
X_2313_ net48 net47 _0700_ vssd1 vssd1 vccd1 vccd1 _0701_ sky130_fd_sc_hd__and3_1
X_1692_ dut.actual_duty_x\[6\] net47 vssd1 vssd1 vccd1 vccd1 _1262_ sky130_fd_sc_hd__xor2_1
X_2244_ _0599_ _0602_ net18 vssd1 vssd1 vccd1 vccd1 _0644_ sky130_fd_sc_hd__o21ai_1
X_2175_ net43 _0544_ _0557_ vssd1 vssd1 vccd1 vccd1 _0578_ sky130_fd_sc_hd__a21bo_1
XFILLER_40_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1959_ net188 net156 vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__xor2_1
XFILLER_0_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_2793_ clknet_leaf_9_clk _0147_ net65 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_200ms\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_2862_ clknet_leaf_3_clk _0215_ net60 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1813_ dut.actual_duty_x\[2\] _0267_ vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__xnor2_2
X_1744_ _0258_ _0260_ _0252_ vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__o21ai_1
X_1675_ net46 dut.actual_duty_x\[7\] vssd1 vssd1 vccd1 vccd1 _1245_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2227_ _0938_ _0629_ vssd1 vssd1 vccd1 vccd1 _0630_ sky130_fd_sc_hd__or2_1
X_2158_ _0545_ _0555_ vssd1 vssd1 vccd1 vccd1 _0561_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2089_ dut.clk_en net165 _0509_ _0511_ vssd1 vssd1 vccd1 vccd1 _0097_ sky130_fd_sc_hd__o22a_1
X_2696__124 vssd1 vssd1 vccd1 vccd1 _2696__124/HI net124 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xteam_02_142 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] team_02_142/LO sky130_fd_sc_hd__conb_1
Xteam_02_120 vssd1 vssd1 vccd1 vccd1 team_02_120/HI gpio_out[32] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_59_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xteam_02_131 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] team_02_131/LO sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1391_ dut.spi.cs_low_counter_q\[4\] _0996_ vssd1 vssd1 vccd1 vccd1 _0997_ sky130_fd_sc_hd__or2_1
X_1460_ net38 net40 net36 vssd1 vssd1 vccd1 vccd1 _1049_ sky130_fd_sc_hd__and3_1
XFILLER_4_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_35_Left_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2012_ _0460_ _0461_ vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__nor2_1
XFILLER_35_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2845_ clknet_leaf_26_clk _0198_ net59 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold101 dut.lcd1602.cnt_200ms\[3\] vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__dlygate4sd3_1
X_1658_ _1234_ net22 _1233_ vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_y.count_d\[11\]
+ sky130_fd_sc_hd__and3b_1
Xhold167 dut.ir_sensor_array.final_sensor_data\[37\] vssd1 vssd1 vccd1 vccd1 net319
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 dut.ir_sensor_array.final_sensor_data\[39\] vssd1 vssd1 vccd1 vccd1 net286
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 dut.clkdiv_inst.counter\[7\] vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__dlygate4sd3_1
X_2776_ clknet_leaf_29_clk _0048_ net50 vssd1 vssd1 vccd1 vccd1 dut.microstep_x.ctr\[20\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold123 dut.microstep_x.ctr\[22\] vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__dlygate4sd3_1
X_1727_ _0240_ _0244_ vssd1 vssd1 vccd1 vccd1 _0245_ sky130_fd_sc_hd__xnor2_1
XFILLER_12_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold156 dut.ir_sensor_array.final_sensor_data\[13\] vssd1 vssd1 vccd1 vccd1 net308
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 dut.ir_sensor_array.bit_count\[4\] vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1589_ dut.pwm_a_inst_y.count_q\[5\] dut.pwm_a_inst_y.count_q\[4\] vssd1 vssd1 vccd1
+ vccd1 _1178_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_64_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_4_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2630_ clknet_leaf_13_clk _0101_ net82 vssd1 vssd1 vccd1 vccd1 dut.spi.shift_reg_q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1512_ _1099_ _1100_ vssd1 vssd1 vccd1 vccd1 _1101_ sky130_fd_sc_hd__nand2_1
X_2561_ dut.ir_sensor_array.final_sensor_data\[27\] dut.ir_sensor_array.final_sensor_data\[26\]
+ net33 vssd1 vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__mux2_1
X_2492_ _0823_ _0833_ _0834_ _0792_ net44 vssd1 vssd1 vccd1 vccd1 _0841_ sky130_fd_sc_hd__o221a_1
X_1374_ dut.spi.clk_counter_q\[3\] dut.spi.clk_counter_q\[2\] _0978_ vssd1 vssd1 vccd1
+ vccd1 _0987_ sky130_fd_sc_hd__and3_1
X_1443_ net14 _1033_ vssd1 vssd1 vccd1 vccd1 _1034_ sky130_fd_sc_hd__nor2_1
XFILLER_63_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2828_ clknet_leaf_3_clk _0181_ net73 vssd1 vssd1 vccd1 vccd1 dut.ball_pos_y\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2759_ clknet_leaf_0_clk _0059_ net52 vssd1 vssd1 vccd1 vccd1 dut.microstep_x.ctr\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout62 net63 vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_4
Xfanout40 dut.actual_duty_y\[4\] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__buf_1
Xfanout51 net52 vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_4
XFILLER_14_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout73 net75 vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__clkbuf_4
Xfanout84 net85 vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__clkbuf_4
XFILLER_13_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload10 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 clkload10/Y sky130_fd_sc_hd__clkinv_2
X_1992_ dut.microstep_x.ctr\[13\] dut.microstep_x.ctr\[14\] _0446_ vssd1 vssd1 vccd1
+ vccd1 _0449_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_15_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2475_ _1186_ _0786_ vssd1 vssd1 vccd1 vccd1 _0827_ sky130_fd_sc_hd__nand2_1
Xclkload21 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 clkload21/Y sky130_fd_sc_hd__inv_6
X_2613_ clknet_leaf_25_clk net299 net60 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2544_ dut.ir_sensor_array.final_sensor_data\[10\] net311 net31 vssd1 vssd1 vccd1
+ vccd1 _0192_ sky130_fd_sc_hd__mux2_1
X_1357_ dut.spi.state_q\[2\] dut.spi.state_q\[0\] vssd1 vssd1 vccd1 vccd1 _0974_ sky130_fd_sc_hd__and2b_1
XFILLER_55_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1288_ net293 vssd1 vssd1 vccd1 vccd1 _0912_ sky130_fd_sc_hd__inv_2
X_1426_ dut.lcd1602.cnt_500hz\[7\] _1021_ vssd1 vssd1 vccd1 vccd1 _1023_ sky130_fd_sc_hd__nand2_1
XFILLER_36_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload4 clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 clkload4/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_21_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2191_ _0589_ _0593_ vssd1 vssd1 vccd1 vccd1 _0594_ sky130_fd_sc_hd__nor2_1
XFILLER_37_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2260_ _0653_ vssd1 vssd1 vccd1 vccd1 _0654_ sky130_fd_sc_hd__inv_2
XFILLER_52_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1975_ _0959_ _0436_ _0438_ vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__or3_1
X_1409_ net189 net13 vssd1 vssd1 vccd1 vccd1 _0020_ sky130_fd_sc_hd__nor2_1
Xhold16 dut.data_in\[9\] vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2458_ net37 _0805_ _0808_ _0787_ net36 vssd1 vssd1 vccd1 vccd1 _0810_ sky130_fd_sc_hd__o221a_1
X_2527_ _0853_ _0855_ _0858_ _0860_ vssd1 vssd1 vccd1 vccd1 _0866_ sky130_fd_sc_hd__or4_1
Xhold38 dut.microstep_x.ctr\[3\] vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 dut.microstep_x.ctr\[2\] vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 dut.lcd1602.cnt_200ms\[16\] vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__dlygate4sd3_1
X_2389_ net205 _0754_ vssd1 vssd1 vccd1 vccd1 _0153_ sky130_fd_sc_hd__xor2_1
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1691_ _1250_ _1260_ vssd1 vssd1 vccd1 vccd1 _1261_ sky130_fd_sc_hd__or2_1
X_1760_ _0258_ _0272_ vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__nand2_1
XFILLER_15_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2312_ _0254_ _0267_ vssd1 vssd1 vccd1 vccd1 _0700_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_48_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2243_ _0553_ _0582_ _0592_ vssd1 vssd1 vccd1 vccd1 _0643_ sky130_fd_sc_hd__or3_1
X_2174_ _0542_ _0575_ _0574_ vssd1 vssd1 vccd1 vccd1 _0577_ sky130_fd_sc_hd__a21o_1
XFILLER_38_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1958_ net185 _0427_ _0428_ vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__a21o_1
X_1889_ net181 _0945_ vssd1 vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__nor2_1
XFILLER_48_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload2_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2861_ clknet_leaf_3_clk _0214_ net60 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[32\]
+ sky130_fd_sc_hd__dfrtp_1
X_2792_ clknet_leaf_9_clk _0146_ net66 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_200ms\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1674_ _0919_ net45 net48 vssd1 vssd1 vccd1 vccd1 _1244_ sky130_fd_sc_hd__and3_1
XFILLER_7_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1743_ _0252_ _0258_ _0260_ vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__or3_1
X_1812_ _0277_ _0329_ vssd1 vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__and2_1
X_2226_ _0608_ _0622_ _0627_ _0628_ vssd1 vssd1 vccd1 vccd1 _0629_ sky130_fd_sc_hd__and4_1
XFILLER_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2157_ _0559_ vssd1 vssd1 vccd1 vccd1 _0560_ sky130_fd_sc_hd__inv_2
X_2088_ net35 _0506_ vssd1 vssd1 vccd1 vccd1 _0511_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout87_A dut.clkdiv_inst.reset_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_02_121 vssd1 vssd1 vccd1 vccd1 team_02_121/HI gpio_out[33] sky130_fd_sc_hd__conb_1
Xteam_02_143 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] team_02_143/LO sky130_fd_sc_hd__conb_1
Xteam_02_110 vssd1 vssd1 vccd1 vccd1 team_02_110/HI gpio_out[22] sky130_fd_sc_hd__conb_1
XFILLER_29_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xteam_02_132 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] team_02_132/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_42_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1390_ _0996_ _0991_ _0995_ vssd1 vssd1 vccd1 vccd1 dut.spi.cs_low_counter_d\[3\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_4_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2011_ dut.microstep_x.ctr\[21\] dut.microstep_x.ctr\[20\] _0459_ vssd1 vssd1 vccd1
+ vccd1 _0461_ sky130_fd_sc_hd__and3_1
X_2844_ clknet_leaf_26_clk _0197_ net57 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_1657_ dut.pwm_a_inst_y.count_q\[10\] dut.pwm_a_inst_y.count_q\[11\] _1230_ vssd1
+ vssd1 vccd1 vccd1 _1234_ sky130_fd_sc_hd__and3_1
X_1588_ _1137_ _1176_ vssd1 vssd1 vccd1 vccd1 _1177_ sky130_fd_sc_hd__and2_1
Xhold135 dut.clkdiv_inst.counter\[14\] vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 dut.ir_sensor_array.final_sensor_data\[29\] vssd1 vssd1 vccd1 vccd1 net320
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 dut.clkdiv_inst.counter\[10\] vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 dut.ir_sensor_array.state\[2\] vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 dut.microstep_x.ctr\[21\] vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__dlygate4sd3_1
X_2775_ clknet_leaf_29_clk _0046_ net50 vssd1 vssd1 vccd1 vccd1 dut.microstep_x.ctr\[19\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold157 dut.microstep_x.ctr\[15\] vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__dlygate4sd3_1
X_1726_ _0920_ _0243_ _0241_ vssd1 vssd1 vccd1 vccd1 _0244_ sky130_fd_sc_hd__o21a_1
Xhold113 dut.clkdiv_inst.counter\[4\] vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__dlygate4sd3_1
X_2209_ _0570_ _0581_ _0611_ vssd1 vssd1 vccd1 vccd1 _0612_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_64_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_2_0__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_4_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1442_ dut.lcd1602.cnt_500hz\[13\] _1032_ vssd1 vssd1 vccd1 vccd1 _1033_ sky130_fd_sc_hd__and2_1
X_1511_ _1093_ _1098_ vssd1 vssd1 vccd1 vccd1 _1100_ sky130_fd_sc_hd__xor2_1
X_2560_ dut.ir_sensor_array.final_sensor_data\[26\] net315 net33 vssd1 vssd1 vccd1
+ vccd1 _0208_ sky130_fd_sc_hd__mux2_1
X_2491_ _0811_ _0812_ _0796_ vssd1 vssd1 vccd1 vccd1 _0840_ sky130_fd_sc_hd__o21ai_1
X_1373_ dut.spi.clk_counter_q\[1\] dut.spi.clk_counter_q\[0\] dut.spi.clk_counter_q\[2\]
+ dut.spi.clk_counter_q\[3\] vssd1 vssd1 vccd1 vccd1 _0986_ sky130_fd_sc_hd__a31o_1
XFILLER_63_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2827_ clknet_leaf_3_clk _0180_ net60 vssd1 vssd1 vccd1 vccd1 dut.ball_pos_y\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_2758_ clknet_leaf_0_clk _0058_ net54 vssd1 vssd1 vccd1 vccd1 dut.microstep_x.ctr\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2689_ clknet_leaf_17_clk dut.pwm_a_inst_y.count_d\[12\] net85 vssd1 vssd1 vccd1
+ vccd1 dut.pwm_a_inst_y.count_q\[12\] sky130_fd_sc_hd__dfrtp_2
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1709_ dut.actual_duty_x\[4\] dut.actual_duty_x\[5\] vssd1 vssd1 vccd1 vccd1 _0227_
+ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_18_Left_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_54_Left_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout85 net86 vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__clkbuf_4
Xfanout41 dut.actual_duty_y\[2\] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_2
Xfanout63 net67 vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__clkbuf_4
Xfanout52 net56 vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__clkbuf_2
Xfanout74 net75 vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_63_Left_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload11 clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 clkload11/Y sky130_fd_sc_hd__inv_6
Xclkload22 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 clkload22/Y sky130_fd_sc_hd__inv_6
X_1991_ net258 _0446_ _0448_ net16 vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__a211oi_1
XFILLER_9_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2612_ clknet_leaf_26_clk _0000_ net60 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_1425_ dut.lcd1602.cnt_500hz\[7\] _1021_ vssd1 vssd1 vccd1 vccd1 _1022_ sky130_fd_sc_hd__or2_1
X_2474_ _1185_ _0787_ _0825_ _1189_ _0824_ vssd1 vssd1 vccd1 vccd1 _0826_ sky130_fd_sc_hd__a221o_1
X_2543_ dut.ir_sensor_array.final_sensor_data\[8\] net311 _0943_ vssd1 vssd1 vccd1
+ vccd1 _0191_ sky130_fd_sc_hd__mux2_1
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1356_ net3 net1 vssd1 vssd1 vccd1 vccd1 dut.clkdiv_inst.reset_n sky130_fd_sc_hd__and2_1
X_1287_ net155 vssd1 vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__inv_2
XFILLER_63_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload5 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 clkload5/Y sky130_fd_sc_hd__inv_6
XFILLER_59_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Left_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2190_ _0582_ _0590_ _0591_ _0588_ vssd1 vssd1 vccd1 vccd1 _0593_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_37_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1974_ _0962_ _0964_ _0965_ _0437_ vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__or4_1
XFILLER_20_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1408_ _1006_ _1011_ vssd1 vssd1 vccd1 vccd1 _1012_ sky130_fd_sc_hd__or2_1
X_2388_ _0754_ _0755_ vssd1 vssd1 vccd1 vccd1 _0152_ sky130_fd_sc_hd__nor2_1
X_2526_ _0861_ _0863_ net29 net28 net316 vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__a32o_1
X_2457_ _0801_ _0803_ _0808_ _0787_ _0804_ vssd1 vssd1 vccd1 vccd1 _0809_ sky130_fd_sc_hd__a221o_1
Xhold39 dut.microstep_y.ctr\[1\] vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 dut.clkdiv_inst.counter\[2\] vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 _0429_ vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1339_ _0958_ vssd1 vssd1 vccd1 vccd1 _0959_ sky130_fd_sc_hd__inv_2
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout72_X net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_60 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1690_ _1246_ _1248_ net47 vssd1 vssd1 vccd1 vccd1 _1260_ sky130_fd_sc_hd__a21oi_1
X_2242_ _0553_ _0571_ _0582_ vssd1 vssd1 vccd1 vccd1 _0642_ sky130_fd_sc_hd__or3_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2311_ net11 _0696_ _0697_ vssd1 vssd1 vccd1 vccd1 _0699_ sky130_fd_sc_hd__a21oi_1
XFILLER_53_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2173_ _0542_ _0575_ _0574_ vssd1 vssd1 vccd1 vccd1 _0576_ sky130_fd_sc_hd__a21oi_1
XFILLER_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1957_ dut.microstep_y.ctr\[29\] dut.microstep_y.ctr\[28\] _0425_ vssd1 vssd1 vccd1
+ vccd1 _0428_ sky130_fd_sc_hd__and3b_1
XFILLER_31_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2509_ dut.ir_sensor_array.final_sensor_data\[24\] dut.ir_sensor_array.final_sensor_data\[25\]
+ vssd1 vssd1 vccd1 vccd1 _0849_ sky130_fd_sc_hd__nor2_1
X_1888_ _0945_ net172 vssd1 vssd1 vccd1 vccd1 _0089_ sky130_fd_sc_hd__nor2_1
XFILLER_0_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_6_Left_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_27_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2791_ clknet_leaf_9_clk _0145_ net65 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_200ms\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_45_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2860_ clknet_leaf_3_clk _0213_ net59 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1811_ _0274_ _0276_ vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__or2_1
X_1673_ _0919_ net45 net48 vssd1 vssd1 vccd1 vccd1 _1243_ sky130_fd_sc_hd__a21oi_1
XFILLER_7_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1742_ _0246_ _0259_ vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__or2_1
X_2225_ _0582_ _0592_ _0604_ _0624_ _0571_ vssd1 vssd1 vccd1 vccd1 _0628_ sky130_fd_sc_hd__o32a_1
X_2156_ dut.lcd1602.currentState\[5\] _0558_ vssd1 vssd1 vccd1 vccd1 _0559_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_18_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_38_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2087_ _0509_ vssd1 vssd1 vccd1 vccd1 _0510_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xteam_02_100 vssd1 vssd1 vccd1 vccd1 team_02_100/HI gpio_out[2] sky130_fd_sc_hd__conb_1
Xteam_02_133 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] team_02_133/LO sky130_fd_sc_hd__conb_1
Xteam_02_111 vssd1 vssd1 vccd1 vccd1 team_02_111/HI gpio_out[23] sky130_fd_sc_hd__conb_1
XFILLER_29_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xteam_02_144 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] team_02_144/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_42_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_32_Left_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2010_ dut.microstep_x.ctr\[20\] _0459_ net254 vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_7_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2774_ clknet_leaf_29_clk _0045_ net50 vssd1 vssd1 vccd1 vccd1 dut.microstep_x.ctr\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_1725_ _0241_ _0242_ vssd1 vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__nand2_1
X_2843_ clknet_leaf_28_clk _0196_ net57 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold136 dut.lcd1602.cnt_500hz\[5\] vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1656_ dut.pwm_a_inst_y.count_q\[10\] dut.pwm_a_inst_y.count_q\[9\] _1229_ dut.pwm_a_inst_y.count_q\[11\]
+ vssd1 vssd1 vccd1 vccd1 _1233_ sky130_fd_sc_hd__a31o_1
X_1587_ _1128_ _1136_ vssd1 vssd1 vccd1 vccd1 _1176_ sky130_fd_sc_hd__nand2_1
Xhold114 dut.microstep_y.ctr\[21\] vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__dlygate4sd3_1
Xhold125 dut.pid_y.y_pid.last_error\[3\] vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 _0001_ vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 dut.ir_sensor_array.final_sensor_data\[16\] vssd1 vssd1 vccd1 vccd1 net310
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold169 dut.ir_sensor_array.final_sensor_data\[21\] vssd1 vssd1 vccd1 vccd1 net321
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold103 dut.microstep_x.ctr\[19\] vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__dlygate4sd3_1
X_2139_ dut.lcd1602.currentState\[3\] dut.lcd1602.currentState\[5\] vssd1 vssd1 vccd1
+ vccd1 _0542_ sky130_fd_sc_hd__nor2_1
X_2208_ net12 _0599_ vssd1 vssd1 vccd1 vccd1 _0611_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_64_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1441_ _1032_ _1018_ _1031_ vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__and3b_1
X_1510_ net38 _1094_ _1095_ vssd1 vssd1 vccd1 vccd1 _1099_ sky130_fd_sc_hd__a21bo_1
X_2490_ net41 _0931_ _0838_ _0839_ vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__a22o_1
X_1372_ net197 _0978_ _0985_ vssd1 vssd1 vccd1 vccd1 dut.spi.clk_counter_d\[2\] sky130_fd_sc_hd__a21oi_1
XFILLER_63_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2826_ clknet_leaf_15_clk _0179_ net82 vssd1 vssd1 vccd1 vccd1 dut.spi.spi_clk_q
+ sky130_fd_sc_hd__dfrtp_1
X_2688_ clknet_leaf_17_clk dut.pwm_a_inst_y.count_d\[11\] net85 vssd1 vssd1 vccd1
+ vccd1 dut.pwm_a_inst_y.count_q\[11\] sky130_fd_sc_hd__dfrtp_1
X_1708_ dut.actual_duty_x\[4\] net47 vssd1 vssd1 vccd1 vccd1 _0226_ sky130_fd_sc_hd__and2_1
X_2757_ clknet_leaf_0_clk _0047_ net54 vssd1 vssd1 vccd1 vccd1 dut.microstep_x.ctr\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1639_ _1221_ _1222_ vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_y.count_d\[4\] sky130_fd_sc_hd__nor2_1
XFILLER_64_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout20 _0518_ vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__buf_2
Xfanout64 net66 vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__clkbuf_4
Xfanout86 net87 vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__clkbuf_2
Xfanout42 dut.actual_duty_y\[0\] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__buf_2
Xfanout31 _0942_ vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_4
Xfanout75 net87 vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__clkbuf_4
Xfanout53 net56 vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__clkbuf_4
XFILLER_60_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1990_ dut.microstep_x.ctr\[13\] _0446_ vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_15_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload23 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 clkload23/X sky130_fd_sc_hd__clkbuf_8
XFILLER_55_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload12 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 clkload12/Y sky130_fd_sc_hd__clkinvlp_4
X_2611_ net298 dut.ir_sensor_array.state\[0\] net35 vssd1 vssd1 vccd1 vccd1 _0225_
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2542_ dut.ir_sensor_array.final_sensor_data\[8\] dut.ir_sensor_array.final_sensor_data\[7\]
+ net32 vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__mux2_1
X_1424_ _1021_ _1018_ _1020_ vssd1 vssd1 vccd1 vccd1 _0031_ sky130_fd_sc_hd__and3b_1
X_2473_ _0780_ _0782_ _0788_ vssd1 vssd1 vccd1 vccd1 _0825_ sky130_fd_sc_hd__o21ai_1
X_1355_ _0973_ vssd1 vssd1 vccd1 vccd1 _0019_ sky130_fd_sc_hd__inv_2
X_1286_ net306 vssd1 vssd1 vccd1 vccd1 _0911_ sky130_fd_sc_hd__inv_2
XFILLER_63_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload6 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 clkload6/Y sky130_fd_sc_hd__clkinv_2
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2809_ clknet_leaf_11_clk _0162_ net68 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.currentState\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_46_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1973_ dut.microstep_x.ctr\[12\] dut.microstep_x.ctr\[14\] dut.microstep_x.ctr\[17\]
+ dut.microstep_x.ctr\[13\] vssd1 vssd1 vccd1 vccd1 _0437_ sky130_fd_sc_hd__or4bb_1
X_2525_ dut.ir_sensor_array.final_sensor_data\[39\] dut.ir_sensor_array.final_sensor_data\[38\]
+ dut.ir_sensor_array.final_sensor_data\[37\] dut.ir_sensor_array.final_sensor_data\[36\]
+ vssd1 vssd1 vccd1 vccd1 _0865_ sky130_fd_sc_hd__nor4_1
X_1407_ _1008_ _1009_ _1010_ vssd1 vssd1 vccd1 vccd1 _1011_ sky130_fd_sc_hd__or3_1
X_2387_ net207 _0752_ vssd1 vssd1 vccd1 vccd1 _0755_ sky130_fd_sc_hd__nor2_1
Xhold29 dut.microstep_y.ctr\[3\] vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__dlygate4sd3_1
X_2456_ _0807_ vssd1 vssd1 vccd1 vccd1 _0808_ sky130_fd_sc_hd__inv_2
X_1338_ dut.microstep_x.ctr\[5\] dut.microstep_x.ctr\[4\] _0957_ vssd1 vssd1 vccd1
+ vccd1 _0958_ sky130_fd_sc_hd__and3_2
Xhold18 _0473_ vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_24_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2241_ net69 _0641_ vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__and2_1
X_2172_ dut.lcd1602.currentState\[4\] _0557_ _0567_ vssd1 vssd1 vccd1 vccd1 _0575_
+ sky130_fd_sc_hd__a21oi_1
X_2310_ net45 _1249_ _0694_ vssd1 vssd1 vccd1 vccd1 _0698_ sky130_fd_sc_hd__mux2_1
XFILLER_2_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1956_ _0426_ _0427_ vssd1 vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__and2_1
X_1887_ dut.microstep_y.ctr\[1\] dut.microstep_y.ctr\[0\] net171 vssd1 vssd1 vccd1
+ vccd1 _0385_ sky130_fd_sc_hd__a21oi_1
X_2508_ dut.ir_sensor_array.final_sensor_data\[31\] dut.ir_sensor_array.final_sensor_data\[30\]
+ dut.ir_sensor_array.final_sensor_data\[29\] dut.ir_sensor_array.final_sensor_data\[28\]
+ vssd1 vssd1 vccd1 vccd1 _0848_ sky130_fd_sc_hd__or4_1
XFILLER_56_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2439_ _0786_ _0790_ vssd1 vssd1 vccd1 vccd1 _0791_ sky130_fd_sc_hd__or2_1
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2790_ clknet_leaf_9_clk _0144_ net70 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_200ms\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1741_ _0922_ _0245_ vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__and2_1
X_1810_ _0293_ _0327_ vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__nor2_1
X_1672_ _0912_ _1242_ net21 vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_y.count_d\[17\]
+ sky130_fd_sc_hd__a21boi_1
XFILLER_7_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2155_ dut.lcd1602.currentState\[3\] _0557_ _0906_ vssd1 vssd1 vccd1 vccd1 _0558_
+ sky130_fd_sc_hd__a21oi_1
X_2224_ _0623_ _0626_ vssd1 vssd1 vccd1 vccd1 _0627_ sky130_fd_sc_hd__nor2_1
XFILLER_53_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2086_ _0500_ _0508_ _0507_ vssd1 vssd1 vccd1 vccd1 _0509_ sky130_fd_sc_hd__o21ai_4
X_1939_ _0416_ _0417_ vssd1 vssd1 vccd1 vccd1 _0080_ sky130_fd_sc_hd__nor2_1
Xteam_02_134 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] team_02_134/LO sky130_fd_sc_hd__conb_1
Xteam_02_112 vssd1 vssd1 vccd1 vccd1 team_02_112/HI gpio_out[24] sky130_fd_sc_hd__conb_1
Xteam_02_101 vssd1 vssd1 vccd1 vccd1 team_02_101/HI gpio_out[6] sky130_fd_sc_hd__conb_1
Xteam_02_145 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] team_02_145/LO sky130_fd_sc_hd__conb_1
XFILLER_29_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold115 dut.clkdiv_inst.counter\[11\] vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__dlygate4sd3_1
X_2773_ clknet_leaf_29_clk _0044_ net51 vssd1 vssd1 vccd1 vccd1 dut.microstep_x.ctr\[17\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold126 dut.microstep_x.ctr\[12\] vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold104 dut.microstep_x.ctr\[9\] vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__dlygate4sd3_1
X_1724_ net48 net49 vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__or2_1
X_2842_ clknet_leaf_28_clk _0195_ net57 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold137 dut.spi.clk_counter_q\[5\] vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 dut.lcd1602.cnt_200ms\[6\] vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__dlygate4sd3_1
X_1655_ dut.pwm_a_inst_y.count_q\[10\] _1230_ _1232_ vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_y.count_d\[10\]
+ sky130_fd_sc_hd__o21a_1
X_1586_ dut.pwm_a_inst_y.count_q\[6\] _1036_ vssd1 vssd1 vccd1 vccd1 _1175_ sky130_fd_sc_hd__xor2_1
Xhold159 dut.ir_sensor_array.final_sensor_data\[9\] vssd1 vssd1 vccd1 vccd1 net311
+ sky130_fd_sc_hd__dlygate4sd3_1
X_2069_ dut.spi.state_q\[1\] _0974_ _0493_ dut.spi.state_q\[2\] vssd1 vssd1 vccd1
+ vccd1 _0494_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_56_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2138_ dut.lcd1602.currentState\[3\] net43 _0906_ vssd1 vssd1 vccd1 vccd1 _0541_
+ sky130_fd_sc_hd__o21a_1
X_2207_ _0585_ _0590_ vssd1 vssd1 vccd1 vccd1 _0610_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_64_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1371_ dut.spi.clk_counter_q\[2\] _0978_ _0983_ vssd1 vssd1 vccd1 vccd1 _0985_ sky130_fd_sc_hd__o21ai_1
X_1440_ dut.lcd1602.cnt_500hz\[11\] dut.lcd1602.cnt_500hz\[12\] _1028_ vssd1 vssd1
+ vccd1 vccd1 _1032_ sky130_fd_sc_hd__and3_1
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2825_ clknet_leaf_24_clk _0178_ net73 vssd1 vssd1 vccd1 vccd1 dut.pid_y.y_pid.last_error\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2687_ clknet_leaf_17_clk dut.pwm_a_inst_y.count_d\[10\] net86 vssd1 vssd1 vccd1
+ vccd1 dut.pwm_a_inst_y.count_q\[10\] sky130_fd_sc_hd__dfrtp_4
X_1638_ dut.pwm_a_inst_y.count_q\[4\] _1219_ net21 vssd1 vssd1 vccd1 vccd1 _1222_
+ sky130_fd_sc_hd__o21ai_1
X_1707_ _1263_ _1276_ vssd1 vssd1 vccd1 vccd1 _1277_ sky130_fd_sc_hd__nand2_1
X_2756_ clknet_leaf_0_clk _0036_ net54 vssd1 vssd1 vccd1 vccd1 dut.microstep_x.ctr\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1569_ dut.pwm_a_inst_y.count_q\[10\] _1039_ vssd1 vssd1 vccd1 vccd1 _1158_ sky130_fd_sc_hd__xor2_1
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout21 _1215_ vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_2
XFILLER_39_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout65 net66 vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_4
Xfanout43 dut.lcd1602.currentState\[2\] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__buf_2
Xfanout87 dut.clkdiv_inst.reset_n vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__buf_2
Xfanout54 net56 vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_4
Xfanout76 net77 vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__clkbuf_4
Xfanout32 _0942_ vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__buf_2
XFILLER_1_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload24 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 clkload24/X sky130_fd_sc_hd__clkbuf_4
Xclkload13 clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 clkload13/Y sky130_fd_sc_hd__inv_6
X_2472_ _0916_ _0797_ _0783_ net42 vssd1 vssd1 vccd1 vccd1 _0824_ sky130_fd_sc_hd__o211a_1
X_2610_ dut.ball_pos_x\[2\] _0944_ _0863_ _0905_ vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__a22o_1
XFILLER_9_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2541_ dut.ir_sensor_array.final_sensor_data\[6\] dut.ir_sensor_array.final_sensor_data\[7\]
+ _0943_ vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__mux2_1
X_1423_ dut.lcd1602.cnt_500hz\[6\] _0934_ vssd1 vssd1 vccd1 vccd1 _1021_ sky130_fd_sc_hd__and2_1
XFILLER_48_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1354_ _0968_ _0970_ _0971_ _0972_ vssd1 vssd1 vccd1 vccd1 _0973_ sky130_fd_sc_hd__or4_1
X_1285_ net156 vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__inv_2
XFILLER_63_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2808_ clknet_leaf_27_clk net15 net58 vssd1 vssd1 vccd1 vccd1 dut.microstep_x.clk_en
+ sky130_fd_sc_hd__dfrtp_4
Xclkload7 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 clkload7/Y sky130_fd_sc_hd__inv_6
XFILLER_59_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2739_ clknet_leaf_6_clk _0081_ net63 vssd1 vssd1 vccd1 vccd1 dut.microstep_y.ctr\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__1356__X dut.clkdiv_inst.reset_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1972_ dut.microstep_x.ctr\[9\] dut.microstep_x.ctr\[10\] _0434_ _0435_ vssd1 vssd1
+ vccd1 vccd1 _0436_ sky130_fd_sc_hd__or4b_1
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2524_ dut.ir_sensor_array.final_sensor_data\[37\] dut.ir_sensor_array.final_sensor_data\[36\]
+ vssd1 vssd1 vccd1 vccd1 _0864_ sky130_fd_sc_hd__nor2_1
X_2455_ _0805_ _0806_ vssd1 vssd1 vccd1 vccd1 _0807_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1406_ dut.lcd1602.cnt_200ms\[14\] dut.lcd1602.cnt_200ms\[17\] dut.lcd1602.cnt_200ms\[16\]
+ dut.lcd1602.cnt_200ms\[15\] vssd1 vssd1 vccd1 vccd1 _1010_ sky130_fd_sc_hd__or4b_1
X_2386_ dut.lcd1602.cnt_200ms\[12\] _0752_ vssd1 vssd1 vccd1 vccd1 _0754_ sky130_fd_sc_hd__and2_1
Xhold19 dut.microstep_y.ctr\[2\] vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__dlygate4sd3_1
X_1337_ dut.microstep_x.ctr\[3\] _0956_ vssd1 vssd1 vccd1 vccd1 _0957_ sky130_fd_sc_hd__and2_1
XFILLER_3_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2240_ dut.data_in\[2\] _0938_ _0631_ _0640_ vssd1 vssd1 vccd1 vccd1 _0641_ sky130_fd_sc_hd__a22o_1
X_2171_ dut.lcd1602.currentState\[3\] dut.lcd1602.currentState\[5\] _0550_ dut.lcd1602.currentState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0574_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_48_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1955_ dut.microstep_y.ctr\[28\] _0425_ vssd1 vssd1 vccd1 vccd1 _0427_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_31_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1886_ net191 net157 vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__xor2_1
X_2438_ dut.actual_duty_y\[0\] _1121_ _0789_ vssd1 vssd1 vccd1 vccd1 _0790_ sky130_fd_sc_hd__a21o_1
X_2507_ dut.ir_sensor_array.final_sensor_data\[29\] dut.ir_sensor_array.final_sensor_data\[28\]
+ vssd1 vssd1 vccd1 vccd1 _0847_ sky130_fd_sc_hd__nor2_1
X_2369_ dut.lcd1602.cnt_200ms\[4\] _1002_ net227 vssd1 vssd1 vccd1 vccd1 _0744_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_39_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1671_ net22 _1241_ _1242_ vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_y.count_d\[16\]
+ sky130_fd_sc_hd__and3_1
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1740_ _0253_ _0257_ vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__or2_1
XFILLER_30_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2154_ net43 _0549_ vssd1 vssd1 vccd1 vccd1 _0557_ sky130_fd_sc_hd__or2_1
X_2223_ _0577_ _0611_ _0625_ _0600_ vssd1 vssd1 vccd1 vccd1 _0626_ sky130_fd_sc_hd__a22o_1
XFILLER_38_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2085_ dut.ball_pos_y\[0\] dut.ball_pos_y\[1\] dut.ball_pos_y\[2\] vssd1 vssd1 vccd1
+ vccd1 _0508_ sky130_fd_sc_hd__a21oi_2
XFILLER_61_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1938_ dut.microstep_y.ctr\[21\] dut.microstep_y.ctr\[20\] _0415_ vssd1 vssd1 vccd1
+ vccd1 _0417_ sky130_fd_sc_hd__and3_1
X_1869_ dut.pwm_a_inst_x.count_q\[10\] dut.pwm_a_inst_x.count_q\[9\] _0371_ dut.pwm_a_inst_x.count_q\[11\]
+ vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__a31o_1
Xteam_02_146 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] team_02_146/LO sky130_fd_sc_hd__conb_1
Xteam_02_113 vssd1 vssd1 vccd1 vccd1 team_02_113/HI gpio_out[25] sky130_fd_sc_hd__conb_1
XFILLER_29_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xteam_02_135 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] team_02_135/LO sky130_fd_sc_hd__conb_1
Xteam_02_102 vssd1 vssd1 vccd1 vccd1 team_02_102/HI gpio_out[14] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_50_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload0_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2841_ clknet_leaf_28_clk _0194_ net57 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold138 dut.spi.clk_counter_d\[5\] vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 dut.microstep_y.ctr\[25\] vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__dlygate4sd3_1
X_1654_ dut.pwm_a_inst_y.count_q\[10\] _1230_ net22 vssd1 vssd1 vccd1 vccd1 _1232_
+ sky130_fd_sc_hd__a21boi_1
Xhold116 dut.microstep_y.ctr\[19\] vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold105 dut.microstep_y.ctr\[18\] vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 dut.ir_sensor_array.final_sensor_data\[34\] vssd1 vssd1 vccd1 vccd1 net301
+ sky130_fd_sc_hd__dlygate4sd3_1
X_2772_ clknet_leaf_28_clk _0043_ net51 vssd1 vssd1 vccd1 vccd1 dut.microstep_x.ctr\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_1723_ net48 net49 vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__nand2_1
X_1585_ _1138_ _1173_ vssd1 vssd1 vccd1 vccd1 _1174_ sky130_fd_sc_hd__and2_1
X_2206_ _0577_ _0591_ _0572_ vssd1 vssd1 vccd1 vccd1 _0609_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_64_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2068_ dut.spi.state_q\[1\] dut.spi.state_q\[0\] vssd1 vssd1 vccd1 vccd1 _0493_ sky130_fd_sc_hd__nor2_1
X_2137_ net294 _0538_ _0540_ _0514_ vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_64_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_9 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1370_ _0983_ vssd1 vssd1 vccd1 vccd1 _0984_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_18_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2824_ clknet_leaf_25_clk _0177_ net73 vssd1 vssd1 vccd1 vccd1 dut.pid_y.y_pid.last_error\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_2686_ clknet_leaf_17_clk dut.pwm_a_inst_y.count_d\[9\] net86 vssd1 vssd1 vccd1 vccd1
+ dut.pwm_a_inst_y.count_q\[9\] sky130_fd_sc_hd__dfrtp_1
X_1637_ dut.pwm_a_inst_y.count_q\[4\] _1219_ vssd1 vssd1 vccd1 vccd1 _1221_ sky130_fd_sc_hd__and2_1
X_2755_ clknet_leaf_12_clk _0066_ net79 vssd1 vssd1 vccd1 vccd1 dut.microstep_y.clk_en
+ sky130_fd_sc_hd__dfrtp_1
X_1706_ net48 _1262_ vssd1 vssd1 vccd1 vccd1 _1276_ sky130_fd_sc_hd__or2_1
X_1568_ _1144_ _1156_ vssd1 vssd1 vccd1 vccd1 _1157_ sky130_fd_sc_hd__nor2_1
X_1499_ _1075_ _1082_ _1086_ vssd1 vssd1 vccd1 vccd1 _1088_ sky130_fd_sc_hd__and3_1
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout22 _1215_ vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout44 dut.microstep_y.clk_en vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__buf_2
Xfanout33 net34 vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_4
Xfanout55 net56 vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_1_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout11 _0673_ vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__buf_2
Xfanout66 net67 vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__buf_2
XFILLER_6_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout77 net78 vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__clkbuf_4
XFILLER_49_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_41_Left_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload25 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 clkload25/Y sky130_fd_sc_hd__inv_8
X_1422_ dut.lcd1602.cnt_500hz\[6\] _0934_ vssd1 vssd1 vccd1 vccd1 _1020_ sky130_fd_sc_hd__or2_1
Xclkload14 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 clkload14/Y sky130_fd_sc_hd__inv_6
X_2471_ _0814_ _0822_ vssd1 vssd1 vccd1 vccd1 _0823_ sky130_fd_sc_hd__or2_1
X_2540_ dut.ir_sensor_array.final_sensor_data\[6\] dut.ir_sensor_array.final_sensor_data\[5\]
+ net32 vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_50_Left_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1284_ net305 vssd1 vssd1 vccd1 vccd1 _0910_ sky130_fd_sc_hd__inv_2
X_1353_ dut.clkdiv_inst.counter\[3\] dut.clkdiv_inst.counter\[5\] dut.clkdiv_inst.counter\[4\]
+ dut.clkdiv_inst.counter\[7\] vssd1 vssd1 vccd1 vccd1 _0972_ sky130_fd_sc_hd__or4b_1
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2807_ clknet_leaf_9_clk _0161_ net66 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_200ms\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_2738_ clknet_leaf_6_clk _0080_ net62 vssd1 vssd1 vccd1 vccd1 dut.microstep_y.ctr\[21\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload8 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 clkload8/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__2670__RESET_B net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2669_ clknet_leaf_14_clk _0032_ net69 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_500hz\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_42_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1971_ dut.microstep_x.ctr\[7\] dut.microstep_x.ctr\[6\] dut.microstep_x.ctr\[15\]
+ dut.microstep_x.ctr\[16\] vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__and4b_1
X_1405_ dut.lcd1602.cnt_200ms\[19\] dut.lcd1602.cnt_200ms\[20\] dut.lcd1602.cnt_200ms\[21\]
+ dut.lcd1602.cnt_200ms\[18\] vssd1 vssd1 vccd1 vccd1 _1009_ sky130_fd_sc_hd__or4bb_1
X_2385_ _0752_ _0753_ vssd1 vssd1 vccd1 vccd1 _0151_ sky130_fd_sc_hd__and2b_1
X_2523_ dut.ir_sensor_array.final_sensor_data\[35\] dut.ir_sensor_array.final_sensor_data\[34\]
+ _0926_ _0862_ vssd1 vssd1 vccd1 vccd1 _0863_ sky130_fd_sc_hd__and4bb_1
X_2454_ net39 _0794_ net38 vssd1 vssd1 vccd1 vccd1 _0806_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_26_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput1 en vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_1
X_1336_ dut.microstep_x.ctr\[1\] dut.microstep_x.ctr\[0\] dut.microstep_x.ctr\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0956_ sky130_fd_sc_hd__and3_1
XFILLER_61_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2170_ _0554_ _0565_ _0570_ vssd1 vssd1 vccd1 vccd1 _0573_ sky130_fd_sc_hd__or3_1
X_1954_ dut.microstep_y.ctr\[28\] _0425_ vssd1 vssd1 vccd1 vccd1 _0426_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_31_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1885_ _0918_ _0384_ net27 vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_x.count_d\[17\]
+ sky130_fd_sc_hd__a21boi_1
X_2506_ _0976_ _0516_ _0846_ vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__and3_1
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2368_ net13 _0743_ vssd1 vssd1 vccd1 vccd1 _0144_ sky130_fd_sc_hd__nand2_1
X_2437_ net41 _1133_ vssd1 vssd1 vccd1 vccd1 _0789_ sky130_fd_sc_hd__nor2_1
XFILLER_29_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1319_ net35 net298 _0941_ dut.ir_sensor_array.state\[1\] vssd1 vssd1 vccd1 vccd1
+ _0001_ sky130_fd_sc_hd__a22o_1
X_2299_ dut.actual_duty_x\[0\] _0672_ vssd1 vssd1 vccd1 vccd1 _0687_ sky130_fd_sc_hd__nor2_1
XFILLER_21_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1670_ dut.pwm_a_inst_y.count_q\[16\] dut.pwm_a_inst_y.count_q\[15\] _1238_ vssd1
+ vssd1 vccd1 vccd1 _1242_ sky130_fd_sc_hd__nand3_1
XFILLER_7_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2222_ _0624_ vssd1 vssd1 vccd1 vccd1 _0625_ sky130_fd_sc_hd__inv_2
X_2153_ _0549_ _0555_ dut.lcd1602.currentState\[3\] vssd1 vssd1 vccd1 vccd1 _0556_
+ sky130_fd_sc_hd__a21o_1
XFILLER_38_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2084_ dut.ball_pos_y\[0\] _0923_ _0501_ vssd1 vssd1 vccd1 vccd1 _0507_ sky130_fd_sc_hd__or3_2
X_1937_ dut.microstep_y.ctr\[20\] _0415_ net266 vssd1 vssd1 vccd1 vccd1 _0416_ sky130_fd_sc_hd__a21oi_1
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1799_ _0314_ _0316_ vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__nor2_1
X_1868_ dut.pwm_a_inst_x.count_q\[10\] _0372_ _0374_ vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_x.count_d\[10\]
+ sky130_fd_sc_hd__o21a_1
Xteam_02_114 vssd1 vssd1 vccd1 vccd1 team_02_114/HI gpio_out[26] sky130_fd_sc_hd__conb_1
Xteam_02_147 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] team_02_147/LO sky130_fd_sc_hd__conb_1
Xteam_02_136 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] team_02_136/LO sky130_fd_sc_hd__conb_1
XFILLER_29_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xteam_02_103 vssd1 vssd1 vccd1 vccd1 team_02_103/HI gpio_out[15] sky130_fd_sc_hd__conb_1
XFILLER_52_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_19_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2771_ clknet_leaf_28_clk _0042_ net51 vssd1 vssd1 vccd1 vccd1 dut.microstep_x.ctr\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_2840_ clknet_leaf_0_clk _0193_ net59 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold139 dut.lcd1602.cnt_500hz\[2\] vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__dlygate4sd3_1
X_1653_ _1230_ _1231_ vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_y.count_d\[9\] sky130_fd_sc_hd__nor2_1
Xhold128 dut.microstep_y.ctr\[22\] vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__dlygate4sd3_1
Xhold117 dut.microstep_y.ctr\[12\] vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__dlygate4sd3_1
X_1584_ _1117_ _1126_ _1137_ vssd1 vssd1 vccd1 vccd1 _1173_ sky130_fd_sc_hd__nand3_1
Xhold106 dut.microstep_x.ctr\[13\] vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__dlygate4sd3_1
X_1722_ net49 _0228_ vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2205_ _0599_ _0602_ _0603_ _0607_ _0594_ vssd1 vssd1 vccd1 vccd1 _0608_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_64_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2136_ dut.spi.bit_counter_q\[3\] _0538_ vssd1 vssd1 vccd1 vccd1 _0540_ sky130_fd_sc_hd__nand2_1
X_2067_ net176 _0491_ vssd1 vssd1 vccd1 vccd1 _0009_ sky130_fd_sc_hd__xnor2_1
XFILLER_1_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout78_A net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2823_ clknet_leaf_19_clk _0176_ net74 vssd1 vssd1 vccd1 vccd1 dut.pid_y.y_pid.last_error\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2754_ clknet_leaf_23_clk _0139_ net75 vssd1 vssd1 vccd1 vccd1 dut.actual_duty_x\[7\]
+ sky130_fd_sc_hd__dfstp_1
X_1705_ _1267_ _1274_ vssd1 vssd1 vccd1 vccd1 _1275_ sky130_fd_sc_hd__or2_1
X_2685_ clknet_leaf_15_clk dut.pwm_a_inst_y.count_d\[8\] net84 vssd1 vssd1 vccd1 vccd1
+ dut.pwm_a_inst_y.count_q\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_48_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1567_ _1072_ _1141_ _1143_ vssd1 vssd1 vccd1 vccd1 _1156_ sky130_fd_sc_hd__and3_1
X_1636_ _1219_ _1220_ net21 vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_y.count_d\[3\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_64_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2119_ _0990_ _0993_ _0494_ vssd1 vssd1 vccd1 vccd1 _0529_ sky130_fd_sc_hd__o21ai_1
XFILLER_58_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1498_ _1082_ _1086_ _1075_ vssd1 vssd1 vccd1 vccd1 _1087_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_1_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout12 _0565_ vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_2
Xfanout67 net72 vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__clkbuf_2
Xfanout34 _0942_ vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__buf_2
XFILLER_22_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout45 dut.actual_duty_x\[7\] vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__buf_2
Xfanout56 net72 vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout78 net87 vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_9_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload15 clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 clkload15/Y sky130_fd_sc_hd__clkinv_4
Xclkload26 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 clkload26/Y sky130_fd_sc_hd__inv_8
XFILLER_9_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1421_ net18 net14 vssd1 vssd1 vccd1 vccd1 _1019_ sky130_fd_sc_hd__or2_1
X_2470_ _0915_ _1183_ vssd1 vssd1 vccd1 vccd1 _0822_ sky130_fd_sc_hd__and2_1
XFILLER_36_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1283_ net157 vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__inv_2
X_1352_ dut.clkdiv_inst.counter\[6\] dut.clkdiv_inst.counter\[11\] dut.clkdiv_inst.counter\[10\]
+ dut.clkdiv_inst.counter\[12\] vssd1 vssd1 vccd1 vccd1 _0971_ sky130_fd_sc_hd__or4b_1
XFILLER_51_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2806_ clknet_leaf_8_clk _0160_ net66 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_200ms\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_2668_ clknet_leaf_14_clk _0031_ net69 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_500hz\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_2737_ clknet_leaf_6_clk _0079_ net62 vssd1 vssd1 vccd1 vccd1 dut.microstep_y.ctr\[20\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload9 clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 clkload9/Y sky130_fd_sc_hd__clkinvlp_4
X_1619_ _1042_ _1146_ _1153_ _1154_ _1207_ vssd1 vssd1 vccd1 vccd1 _1208_ sky130_fd_sc_hd__a221o_1
X_2599_ dut.ir_sensor_array.final_sensor_data\[19\] dut.ir_sensor_array.final_sensor_data\[18\]
+ _0895_ _0859_ vssd1 vssd1 vccd1 vccd1 _0896_ sky130_fd_sc_hd__o31a_1
XANTENNA_input2_A gpio_in[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_23_Left_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1970_ dut.microstep_x.ctr\[8\] dut.microstep_x.ctr\[11\] vssd1 vssd1 vccd1 vccd1
+ _0434_ sky130_fd_sc_hd__nand2_1
XFILLER_53_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2522_ dut.ir_sensor_array.final_sensor_data\[32\] net28 vssd1 vssd1 vccd1 vccd1
+ _0862_ sky130_fd_sc_hd__nor2_1
X_1404_ dut.lcd1602.cnt_200ms\[8\] dut.lcd1602.cnt_200ms\[9\] _1007_ vssd1 vssd1 vccd1
+ vccd1 _1008_ sky130_fd_sc_hd__nand3b_1
X_2384_ dut.lcd1602.cnt_200ms\[9\] dut.lcd1602.cnt_200ms\[10\] _0748_ dut.lcd1602.cnt_200ms\[11\]
+ vssd1 vssd1 vccd1 vccd1 _0753_ sky130_fd_sc_hd__a31o_1
X_1335_ _0948_ _0949_ _0950_ _0955_ vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__nor4_2
X_2453_ _1078_ _0794_ vssd1 vssd1 vccd1 vccd1 _0805_ sky130_fd_sc_hd__or2_2
XFILLER_5_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput2 gpio_in[6] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_34_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout60_A net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1953_ _0424_ _0425_ vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__nor2_1
XFILLER_33_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1884_ net26 _0383_ _0384_ vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_x.count_d\[16\]
+ sky130_fd_sc_hd__and3_1
XFILLER_21_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2505_ dut.spi.spi_clk_q _0982_ vssd1 vssd1 vccd1 vccd1 _0846_ sky130_fd_sc_hd__or2_1
X_2367_ net296 _1002_ vssd1 vssd1 vccd1 vccd1 _0743_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_39_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2436_ _0766_ _0777_ _0787_ vssd1 vssd1 vccd1 vccd1 _0788_ sky130_fd_sc_hd__o21ai_2
X_1318_ net35 _0940_ vssd1 vssd1 vccd1 vccd1 _0941_ sky130_fd_sc_hd__nand2_1
X_2298_ _0673_ _0685_ vssd1 vssd1 vccd1 vccd1 _0686_ sky130_fd_sc_hd__nand2_1
XFILLER_12_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2221_ _0582_ _0587_ vssd1 vssd1 vccd1 vccd1 _0624_ sky130_fd_sc_hd__or2_1
X_2152_ dut.lcd1602.currentState\[0\] net43 vssd1 vssd1 vccd1 vccd1 _0555_ sky130_fd_sc_hd__nand2_1
X_2083_ dut.ball_pos_x\[2\] _0502_ _0503_ _0505_ vssd1 vssd1 vccd1 vccd1 _0506_ sky130_fd_sc_hd__o211a_1
X_1936_ net194 _0415_ vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_26_Left_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1867_ dut.pwm_a_inst_x.count_q\[10\] _0372_ net26 vssd1 vssd1 vccd1 vccd1 _0374_
+ sky130_fd_sc_hd__a21boi_1
XPHY_EDGE_ROW_10_Left_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1798_ dut.pwm_a_inst_x.count_q\[4\] _0315_ _0295_ vssd1 vssd1 vccd1 vccd1 _0316_
+ sky130_fd_sc_hd__o21ba_1
Xteam_02_115 vssd1 vssd1 vccd1 vccd1 team_02_115/HI gpio_out[27] sky130_fd_sc_hd__conb_1
Xteam_02_137 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] team_02_137/LO sky130_fd_sc_hd__conb_1
Xteam_02_104 vssd1 vssd1 vccd1 vccd1 team_02_104/HI gpio_out[16] sky130_fd_sc_hd__conb_1
XFILLER_44_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2419_ _0503_ _0508_ dut.ball_pos_x\[2\] _0499_ vssd1 vssd1 vccd1 vccd1 _0771_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_29_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xteam_02_126 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] team_02_126/LO sky130_fd_sc_hd__conb_1
Xteam_02_148 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] team_02_148/LO sky130_fd_sc_hd__conb_1
XFILLER_52_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2770_ clknet_leaf_29_clk _0041_ net51 vssd1 vssd1 vccd1 vccd1 dut.microstep_x.ctr\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_1721_ _0231_ _0238_ vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__or2_1
Xhold107 dut.lcd1602.cnt_200ms\[1\] vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__dlygate4sd3_1
X_1652_ dut.pwm_a_inst_y.count_q\[9\] _1229_ net22 vssd1 vssd1 vccd1 vccd1 _1231_
+ sky130_fd_sc_hd__o21ai_1
X_1583_ _1139_ _1171_ vssd1 vssd1 vccd1 vccd1 _1172_ sky130_fd_sc_hd__and2_1
Xhold118 dut.microstep_x.ctr\[10\] vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 dut.clkdiv_inst.counter\[5\] vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2135_ net282 _0537_ _0539_ _0514_ vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__o211a_1
X_2204_ _0598_ _0606_ vssd1 vssd1 vccd1 vccd1 _0607_ sky130_fd_sc_hd__nor2_1
XFILLER_26_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2066_ _0491_ _0492_ vssd1 vssd1 vccd1 vccd1 _0008_ sky130_fd_sc_hd__and2_1
X_1919_ dut.microstep_y.ctr\[13\] dut.microstep_y.ctr\[14\] _0402_ vssd1 vssd1 vccd1
+ vccd1 _0405_ sky130_fd_sc_hd__and3_1
XFILLER_1_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2684_ clknet_leaf_13_clk dut.pwm_a_inst_y.count_d\[7\] net84 vssd1 vssd1 vccd1 vccd1
+ dut.pwm_a_inst_y.count_q\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_31_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2822_ clknet_leaf_20_clk _0175_ net77 vssd1 vssd1 vccd1 vccd1 dut.actual_duty_y\[7\]
+ sky130_fd_sc_hd__dfstp_1
X_2753_ clknet_leaf_23_clk _0138_ net75 vssd1 vssd1 vccd1 vccd1 dut.actual_duty_x\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_1704_ _0920_ _1266_ vssd1 vssd1 vccd1 vccd1 _1274_ sky130_fd_sc_hd__and2_1
X_1566_ _1148_ _1150_ vssd1 vssd1 vccd1 vccd1 _1155_ sky130_fd_sc_hd__nor2_1
X_1635_ dut.pwm_a_inst_y.count_q\[2\] dut.pwm_a_inst_y.count_q\[1\] dut.pwm_a_inst_y.count_q\[0\]
+ dut.pwm_a_inst_y.count_q\[3\] vssd1 vssd1 vccd1 vccd1 _1220_ sky130_fd_sc_hd__a31o_1
X_1497_ _1083_ _1085_ vssd1 vssd1 vccd1 vccd1 _1086_ sky130_fd_sc_hd__nand2_1
X_2118_ net177 _0517_ _0519_ net192 _0528_ vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__a221o_1
X_2049_ net292 _0480_ _0482_ _0019_ vssd1 vssd1 vccd1 vccd1 _0017_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_1_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout13 _1012_ vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_52_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_18_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout68 net71 vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__clkbuf_4
Xfanout79 net87 vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__clkbuf_4
Xfanout35 dut.clk_en vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__buf_2
Xfanout46 dut.actual_duty_x\[6\] vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_2
Xfanout57 net58 vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_9_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload16 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 clkload16/Y sky130_fd_sc_hd__inv_6
Xclkload27 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 clkload27/Y sky130_fd_sc_hd__inv_6
X_1420_ net18 net14 vssd1 vssd1 vccd1 vccd1 _1018_ sky130_fd_sc_hd__nor2_1
X_1351_ _0969_ vssd1 vssd1 vccd1 vccd1 _0970_ sky130_fd_sc_hd__inv_2
XFILLER_48_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1282_ net154 vssd1 vssd1 vccd1 vccd1 _0909_ sky130_fd_sc_hd__inv_2
X_2805_ clknet_leaf_8_clk _0159_ net65 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_200ms\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_51_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2667_ clknet_leaf_10_clk _0030_ net69 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_500hz\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_1618_ dut.pwm_a_inst_y.count_q\[13\] _1041_ dut.pwm_a_inst_y.count_q\[14\] vssd1
+ vssd1 vccd1 vccd1 _1207_ sky130_fd_sc_hd__a21oi_1
X_2736_ clknet_leaf_5_clk _0077_ net62 vssd1 vssd1 vccd1 vccd1 dut.microstep_y.ctr\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_1549_ _1126_ _1137_ _1117_ vssd1 vssd1 vccd1 vccd1 _1138_ sky130_fd_sc_hd__a21o_1
X_2598_ dut.ir_sensor_array.final_sensor_data\[23\] dut.ir_sensor_array.final_sensor_data\[22\]
+ _0894_ _0857_ vssd1 vssd1 vccd1 vccd1 _0895_ sky130_fd_sc_hd__o31a_1
XFILLER_54_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2521_ _0856_ _0858_ _0860_ _0851_ vssd1 vssd1 vccd1 vccd1 _0861_ sky130_fd_sc_hd__o31ai_1
X_1403_ dut.lcd1602.cnt_200ms\[13\] dut.lcd1602.cnt_200ms\[12\] dut.lcd1602.cnt_200ms\[11\]
+ dut.lcd1602.cnt_200ms\[10\] vssd1 vssd1 vccd1 vccd1 _1007_ sky130_fd_sc_hd__and4b_1
X_2383_ dut.lcd1602.cnt_200ms\[9\] dut.lcd1602.cnt_200ms\[11\] dut.lcd1602.cnt_200ms\[10\]
+ _0748_ vssd1 vssd1 vccd1 vccd1 _0752_ sky130_fd_sc_hd__and4_1
X_1334_ _0951_ _0952_ _0953_ _0954_ vssd1 vssd1 vccd1 vccd1 _0955_ sky130_fd_sc_hd__or4_1
X_2452_ _0792_ _0796_ _0801_ _0803_ _0800_ vssd1 vssd1 vccd1 vccd1 _0804_ sky130_fd_sc_hd__o221a_1
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput3 nrst vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_34_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2719_ clknet_leaf_2_clk _0089_ net55 vssd1 vssd1 vccd1 vccd1 dut.microstep_y.ctr\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_38_Left_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1952_ dut.microstep_y.ctr\[27\] dut.microstep_y.ctr\[26\] _0423_ vssd1 vssd1 vccd1
+ vccd1 _0425_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_31_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1883_ dut.pwm_a_inst_x.count_q\[16\] dut.pwm_a_inst_x.count_q\[15\] _0380_ vssd1
+ vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__nand3_1
XPHY_EDGE_ROW_47_Left_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2435_ _0767_ _0785_ vssd1 vssd1 vccd1 vccd1 _0787_ sky130_fd_sc_hd__or2_2
X_2504_ dut.pid_y.y_pid.last_error\[2\] _0766_ net35 vssd1 vssd1 vccd1 vccd1 _0178_
+ sky130_fd_sc_hd__mux2_1
X_2366_ _1002_ _0742_ net13 vssd1 vssd1 vccd1 vccd1 _0143_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_39_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1317_ dut.ir_sensor_array.bit_count\[4\] dut.ir_sensor_array.bit_count\[3\] _0939_
+ dut.ir_sensor_array.bit_count\[5\] vssd1 vssd1 vccd1 vccd1 _0940_ sky130_fd_sc_hd__o31a_1
X_2297_ _0269_ _0275_ vssd1 vssd1 vccd1 vccd1 _0685_ sky130_fd_sc_hd__or2_1
XFILLER_64_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_56_Left_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2151_ _0547_ _0553_ vssd1 vssd1 vccd1 vccd1 _0554_ sky130_fd_sc_hd__nand2b_1
X_2220_ _0602_ _0604_ vssd1 vssd1 vccd1 vccd1 _0623_ sky130_fd_sc_hd__nor2_1
X_2082_ _0499_ _0504_ dut.ball_pos_x\[2\] vssd1 vssd1 vccd1 vccd1 _0505_ sky130_fd_sc_hd__o21ai_1
X_1935_ _0414_ _0415_ vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__nor2_1
X_1866_ _0372_ _0373_ vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_x.count_d\[9\] sky130_fd_sc_hd__nor2_1
X_1797_ dut.pwm_a_inst_x.count_q\[8\] dut.pwm_a_inst_x.count_q\[7\] dut.pwm_a_inst_x.count_q\[6\]
+ dut.pwm_a_inst_x.count_q\[5\] vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__or4_1
Xteam_02_116 vssd1 vssd1 vccd1 vccd1 team_02_116/HI gpio_out[28] sky130_fd_sc_hd__conb_1
Xteam_02_105 vssd1 vssd1 vccd1 vccd1 team_02_105/HI gpio_out[17] sky130_fd_sc_hd__conb_1
X_2418_ dut.ball_pos_x\[1\] dut.ball_pos_x\[0\] dut.ball_pos_x\[2\] _0504_ vssd1 vssd1
+ vccd1 vccd1 _0770_ sky130_fd_sc_hd__or4_1
Xteam_02_127 vssd1 vssd1 vccd1 vccd1 gpio_oeb[1] team_02_127/LO sky130_fd_sc_hd__conb_1
Xteam_02_138 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] team_02_138/LO sky130_fd_sc_hd__conb_1
XFILLER_44_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xteam_02_149 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] team_02_149/LO sky130_fd_sc_hd__conb_1
X_2349_ net284 dut.microstep_x.clk_en _0733_ vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__o21ba_1
XFILLER_16_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold108 _0740_ vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__dlygate4sd3_1
X_1651_ dut.pwm_a_inst_y.count_q\[9\] _1229_ vssd1 vssd1 vccd1 vccd1 _1230_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_41_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1720_ _0921_ _0230_ vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__and2_1
Xhold119 dut.microstep_y.ctr\[13\] vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__dlygate4sd3_1
X_1582_ _1105_ _1115_ _1138_ vssd1 vssd1 vccd1 vccd1 _1171_ sky130_fd_sc_hd__nand3_1
X_2134_ _0538_ vssd1 vssd1 vccd1 vccd1 _0539_ sky130_fd_sc_hd__inv_2
X_2203_ _0585_ _0591_ _0605_ vssd1 vssd1 vccd1 vccd1 _0606_ sky130_fd_sc_hd__and3b_1
X_2065_ dut.clkdiv_inst.counter\[15\] _0489_ vssd1 vssd1 vccd1 vccd1 _0492_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_64_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1918_ net271 _0402_ _0404_ net17 vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__a211oi_1
X_1849_ _0361_ _0362_ net27 vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_x.count_d\[3\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_27_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_20_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_4_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2821_ clknet_leaf_20_clk _0174_ net76 vssd1 vssd1 vccd1 vccd1 dut.actual_duty_y\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_11_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2683_ clknet_leaf_13_clk dut.pwm_a_inst_y.count_d\[6\] net84 vssd1 vssd1 vccd1 vccd1
+ dut.pwm_a_inst_y.count_q\[6\] sky130_fd_sc_hd__dfrtp_1
X_1634_ dut.pwm_a_inst_y.count_q\[2\] dut.pwm_a_inst_y.count_q\[3\] dut.pwm_a_inst_y.count_q\[1\]
+ dut.pwm_a_inst_y.count_q\[0\] vssd1 vssd1 vccd1 vccd1 _1219_ sky130_fd_sc_hd__and4_1
XFILLER_31_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2752_ clknet_leaf_23_clk _0137_ net75 vssd1 vssd1 vccd1 vccd1 dut.actual_duty_x\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_1703_ _1271_ _1272_ vssd1 vssd1 vccd1 vccd1 _1273_ sky130_fd_sc_hd__nand2_1
X_1565_ net36 _1145_ _1042_ vssd1 vssd1 vccd1 vccd1 _1154_ sky130_fd_sc_hd__o21a_1
XFILLER_39_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1496_ _1082_ _1084_ vssd1 vssd1 vccd1 vccd1 _1085_ sky130_fd_sc_hd__and2_1
X_2117_ dut.data_in\[9\] dut.lcd1602.out_valid _0513_ vssd1 vssd1 vccd1 vccd1 _0528_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_52_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2048_ dut.clkdiv_inst.counter\[8\] _0480_ vssd1 vssd1 vccd1 vccd1 _0482_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_1_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout14 _1012_ vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_2
Xfanout69 net71 vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__clkbuf_4
XANTENNA__2814__RESET_B net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout36 dut.actual_duty_y\[7\] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_2
Xfanout47 dut.actual_duty_x\[5\] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__buf_2
XFILLER_13_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout58 net72 vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_9_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout83_A net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload17 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 clkload17/Y sky130_fd_sc_hd__inv_8
X_1281_ net289 vssd1 vssd1 vccd1 vccd1 _0908_ sky130_fd_sc_hd__inv_2
X_1350_ dut.clkdiv_inst.counter\[1\] dut.clkdiv_inst.counter\[0\] dut.clkdiv_inst.counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0969_ sky130_fd_sc_hd__and3_1
XFILLER_63_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_0_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2804_ clknet_leaf_8_clk _0158_ net64 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_200ms\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_2666_ clknet_leaf_9_clk _0029_ net69 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_500hz\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1617_ _1153_ _1154_ _1205_ _1151_ vssd1 vssd1 vccd1 vccd1 _1206_ sky130_fd_sc_hd__o211a_1
X_2735_ clknet_leaf_5_clk _0076_ net62 vssd1 vssd1 vccd1 vccd1 dut.microstep_y.ctr\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_2597_ dut.ir_sensor_array.final_sensor_data\[11\] dut.ir_sensor_array.final_sensor_data\[10\]
+ _0893_ _0854_ vssd1 vssd1 vccd1 vccd1 _0894_ sky130_fd_sc_hd__o31a_1
X_1548_ _1128_ _1136_ vssd1 vssd1 vccd1 vccd1 _1137_ sky130_fd_sc_hd__or2_1
XFILLER_39_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1479_ _1066_ _1067_ net41 vssd1 vssd1 vccd1 vccd1 _1068_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_37_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_45 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1402_ dut.lcd1602.cnt_200ms\[7\] _1004_ vssd1 vssd1 vccd1 vccd1 _1006_ sky130_fd_sc_hd__nand2_1
X_2451_ net39 _0794_ vssd1 vssd1 vccd1 vccd1 _0803_ sky130_fd_sc_hd__xnor2_1
X_2520_ dut.ir_sensor_array.final_sensor_data\[16\] dut.ir_sensor_array.final_sensor_data\[19\]
+ dut.ir_sensor_array.final_sensor_data\[18\] dut.ir_sensor_array.final_sensor_data\[17\]
+ vssd1 vssd1 vccd1 vccd1 _0860_ sky130_fd_sc_hd__or4_1
X_2382_ net203 _0750_ vssd1 vssd1 vccd1 vccd1 _0150_ sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_leaf_17_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1333_ dut.microstep_y.ctr\[23\] dut.microstep_y.ctr\[22\] dut.microstep_y.ctr\[25\]
+ dut.microstep_y.ctr\[24\] vssd1 vssd1 vccd1 vccd1 _0954_ sky130_fd_sc_hd__or4_1
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_2_1__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_34_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2718_ clknet_leaf_2_clk _0078_ net55 vssd1 vssd1 vccd1 vccd1 dut.microstep_y.ctr\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2649_ clknet_leaf_13_clk _0120_ vssd1 vssd1 vccd1 vccd1 dut.data_in\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1951_ dut.microstep_y.ctr\[26\] _0423_ net224 vssd1 vssd1 vccd1 vccd1 _0424_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_31_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1882_ dut.pwm_a_inst_x.count_q\[15\] dut.pwm_a_inst_x.count_q\[14\] _0379_ dut.pwm_a_inst_x.count_q\[16\]
+ vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__a31o_1
X_2365_ net253 _1001_ vssd1 vssd1 vccd1 vccd1 _0742_ sky130_fd_sc_hd__nor2_1
X_2434_ _0767_ _0785_ vssd1 vssd1 vccd1 vccd1 _0786_ sky130_fd_sc_hd__nor2_1
X_2503_ net277 _0772_ net35 vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1316_ dut.ir_sensor_array.bit_count\[2\] dut.ir_sensor_array.bit_count\[1\] vssd1
+ vssd1 vccd1 vccd1 _0939_ sky130_fd_sc_hd__and2_1
XFILLER_24_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2296_ net49 _0269_ vssd1 vssd1 vccd1 vccd1 _0684_ sky130_fd_sc_hd__xnor2_1
XFILLER_64_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2150_ _0551_ _0552_ dut.lcd1602.currentState\[5\] vssd1 vssd1 vccd1 vccd1 _0553_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_38_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2081_ dut.ball_pos_y\[0\] dut.ball_pos_y\[2\] dut.ball_pos_y\[1\] vssd1 vssd1 vccd1
+ vccd1 _0504_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_44_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1934_ dut.microstep_y.ctr\[19\] _0413_ vssd1 vssd1 vccd1 vccd1 _0415_ sky130_fd_sc_hd__and2_1
XFILLER_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1796_ _0237_ _0284_ vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__xnor2_1
X_1865_ dut.pwm_a_inst_x.count_q\[9\] _0371_ net26 vssd1 vssd1 vccd1 vccd1 _0373_
+ sky130_fd_sc_hd__o21ai_1
Xteam_02_139 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] team_02_139/LO sky130_fd_sc_hd__conb_1
Xteam_02_117 vssd1 vssd1 vccd1 vccd1 team_02_117/HI gpio_out[29] sky130_fd_sc_hd__conb_1
X_2417_ dut.pid_y.y_pid.last_error\[2\] _0767_ vssd1 vssd1 vccd1 vccd1 _0769_ sky130_fd_sc_hd__and2_1
Xteam_02_106 vssd1 vssd1 vccd1 vccd1 team_02_106/HI gpio_out[18] sky130_fd_sc_hd__conb_1
Xteam_02_128 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] team_02_128/LO sky130_fd_sc_hd__conb_1
X_2348_ _0711_ _0720_ _0732_ dut.microstep_x.clk_en vssd1 vssd1 vccd1 vccd1 _0733_
+ sky130_fd_sc_hd__o211a_1
XFILLER_37_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2279_ _0506_ _0510_ dut.pid_x.x_pid.last_error\[3\] vssd1 vssd1 vccd1 vccd1 _0667_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_20_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1650_ _1229_ net21 _1228_ vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_y.count_d\[8\]
+ sky130_fd_sc_hd__and3b_1
X_1581_ _1036_ _1037_ _1169_ vssd1 vssd1 vccd1 vccd1 _1170_ sky130_fd_sc_hd__o21a_1
Xhold109 dut.microstep_y.ctr\[10\] vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__dlygate4sd3_1
X_2202_ _0604_ vssd1 vssd1 vccd1 vccd1 _0605_ sky130_fd_sc_hd__inv_2
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2133_ dut.spi.bit_counter_q\[0\] dut.spi.bit_counter_q\[1\] dut.spi.bit_counter_q\[2\]
+ _0517_ vssd1 vssd1 vccd1 vccd1 _0538_ sky130_fd_sc_hd__and4_1
X_2064_ dut.clkdiv_inst.counter\[15\] _0489_ vssd1 vssd1 vccd1 vccd1 _0491_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_64_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1917_ dut.microstep_y.ctr\[13\] _0402_ vssd1 vssd1 vccd1 vccd1 _0404_ sky130_fd_sc_hd__nor2_1
X_1779_ dut.pwm_a_inst_x.count_q\[10\] dut.pwm_a_inst_x.count_q\[9\] _0295_ dut.pwm_a_inst_x.count_q\[11\]
+ vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__a31o_1
X_1848_ dut.pwm_a_inst_x.count_q\[2\] dut.pwm_a_inst_x.count_q\[1\] dut.pwm_a_inst_x.count_q\[0\]
+ dut.pwm_a_inst_x.count_q\[3\] vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__a31o_1
XFILLER_57_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2820_ clknet_leaf_20_clk _0173_ net77 vssd1 vssd1 vccd1 vccd1 dut.actual_duty_y\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2751_ clknet_leaf_27_clk _0136_ net75 vssd1 vssd1 vccd1 vccd1 dut.actual_duty_x\[4\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_16_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1564_ _1041_ _1152_ vssd1 vssd1 vccd1 vccd1 _1153_ sky130_fd_sc_hd__and2_1
X_2682_ clknet_leaf_18_clk dut.pwm_a_inst_y.count_d\[5\] net86 vssd1 vssd1 vccd1 vccd1
+ dut.pwm_a_inst_y.count_q\[5\] sky130_fd_sc_hd__dfrtp_1
X_1633_ net21 _1217_ _1218_ vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_y.count_d\[2\]
+ sky130_fd_sc_hd__and3_1
X_1702_ _1259_ _1268_ _1270_ vssd1 vssd1 vccd1 vccd1 _1272_ sky130_fd_sc_hd__o21ai_1
XFILLER_58_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1495_ _1077_ _1081_ vssd1 vssd1 vccd1 vccd1 _1084_ sky130_fd_sc_hd__nand2_1
X_2116_ dut.spi.shift_reg_q\[7\] _0517_ _0519_ net177 vssd1 vssd1 vccd1 vccd1 _0108_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout37 dut.actual_duty_y\[6\] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__buf_2
X_2047_ net264 _0478_ _0481_ vssd1 vssd1 vccd1 vccd1 _0016_ sky130_fd_sc_hd__o21a_1
Xfanout26 net27 vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_1_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout48 dut.actual_duty_x\[4\] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__buf_2
Xfanout59 net61 vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_4
XANTENNA__2854__RESET_B net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload18 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 clkload18/Y sky130_fd_sc_hd__inv_6
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1280_ dut.ir_sensor_array.state\[2\] vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.latch
+ sky130_fd_sc_hd__inv_2
XFILLER_36_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2803_ clknet_leaf_8_clk _0157_ net64 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_200ms\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_2734_ clknet_leaf_5_clk _0075_ net62 vssd1 vssd1 vccd1 vccd1 dut.microstep_y.ctr\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_2665_ clknet_leaf_9_clk _0028_ net70 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_500hz\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1616_ _1157_ _1158_ _1204_ _1155_ vssd1 vssd1 vccd1 vccd1 _1205_ sky130_fd_sc_hd__a211o_1
X_1547_ _1130_ _1131_ _1135_ vssd1 vssd1 vccd1 vccd1 _1136_ sky130_fd_sc_hd__a21oi_1
XFILLER_8_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2596_ dut.ir_sensor_array.final_sensor_data\[14\] dut.ir_sensor_array.final_sensor_data\[15\]
+ _0892_ _0852_ vssd1 vssd1 vccd1 vccd1 _0893_ sky130_fd_sc_hd__o31a_1
XFILLER_39_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1478_ net36 _1045_ _1065_ vssd1 vssd1 vccd1 vccd1 _1067_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_37_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1401_ dut.lcd1602.cnt_200ms\[7\] dut.lcd1602.cnt_200ms\[6\] _1003_ vssd1 vssd1 vccd1
+ vccd1 _1005_ sky130_fd_sc_hd__and3_1
X_2381_ _0750_ _0751_ vssd1 vssd1 vccd1 vccd1 _0149_ sky130_fd_sc_hd__and2_1
X_2450_ _0801_ vssd1 vssd1 vccd1 vccd1 _0802_ sky130_fd_sc_hd__inv_2
XFILLER_5_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1332_ dut.microstep_y.ctr\[27\] dut.microstep_y.ctr\[26\] dut.microstep_y.ctr\[29\]
+ dut.microstep_y.ctr\[28\] vssd1 vssd1 vccd1 vccd1 _0953_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_34_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2717_ clknet_leaf_1_clk _0067_ net55 vssd1 vssd1 vccd1 vccd1 dut.microstep_y.ctr\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2648_ clknet_leaf_10_clk _0119_ vssd1 vssd1 vccd1 vccd1 dut.data_in\[2\] sky130_fd_sc_hd__dfxtp_1
X_2579_ dut.ir_sensor_array.final_sensor_data\[12\] _0876_ dut.ir_sensor_array.final_sensor_data\[11\]
+ vssd1 vssd1 vccd1 vccd1 _0877_ sky130_fd_sc_hd__o21ba_1
XFILLER_35_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1950_ net212 _0423_ vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__xor2_1
XFILLER_21_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2502_ net173 _0775_ dut.clk_en vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__mux2_1
X_1881_ net283 _0380_ _0382_ vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_x.count_d\[15\]
+ sky130_fd_sc_hd__a21oi_1
X_1315_ _0938_ vssd1 vssd1 vccd1 vccd1 dut.lcd1602.lcd_ctrl sky130_fd_sc_hd__inv_2
X_2364_ _1001_ _0741_ net13 vssd1 vssd1 vccd1 vccd1 _0142_ sky130_fd_sc_hd__o21ai_1
X_2433_ _0768_ _0777_ vssd1 vssd1 vccd1 vccd1 _0785_ sky130_fd_sc_hd__nor2_1
XFILLER_52_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2295_ _0512_ _0666_ _0509_ vssd1 vssd1 vccd1 vccd1 _0683_ sky130_fd_sc_hd__a21o_1
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_2_0__f_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_16_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2080_ dut.ball_pos_y\[1\] dut.ball_pos_y\[2\] _0500_ vssd1 vssd1 vccd1 vccd1 _0503_
+ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_44_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1933_ net268 _0413_ vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__nor2_1
X_1795_ _0296_ _0312_ vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__nand2_1
X_1864_ dut.pwm_a_inst_x.count_q\[9\] _0371_ vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__and2_1
Xteam_02_107 vssd1 vssd1 vccd1 vccd1 team_02_107/HI gpio_out[19] sky130_fd_sc_hd__conb_1
XFILLER_29_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2416_ dut.pid_y.y_pid.last_error\[2\] _0767_ vssd1 vssd1 vccd1 vccd1 _0768_ sky130_fd_sc_hd__nor2_1
Xteam_02_118 vssd1 vssd1 vccd1 vccd1 team_02_118/HI gpio_out[30] sky130_fd_sc_hd__conb_1
Xteam_02_129 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] team_02_129/LO sky130_fd_sc_hd__conb_1
X_2347_ _0684_ _0722_ _0731_ _0719_ vssd1 vssd1 vccd1 vccd1 _0732_ sky130_fd_sc_hd__a211o_1
X_2278_ _0509_ _0665_ _0664_ vssd1 vssd1 vccd1 vccd1 _0666_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_50_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout61_X net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1580_ dut.pwm_a_inst_y.count_q\[6\] _1036_ dut.pwm_a_inst_y.count_q\[7\] vssd1 vssd1
+ vccd1 vccd1 _1169_ sky130_fd_sc_hd__o21ai_1
XFILLER_7_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2132_ _0514_ net20 _0536_ vssd1 vssd1 vccd1 vccd1 _0537_ sky130_fd_sc_hd__a21oi_1
X_2201_ _0553_ _0586_ vssd1 vssd1 vccd1 vccd1 _0604_ sky130_fd_sc_hd__or2_1
XFILLER_3_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2063_ _0489_ _0490_ vssd1 vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_14_Left_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1916_ _0402_ _0403_ vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__nor2_1
X_1847_ dut.pwm_a_inst_x.count_q\[3\] dut.pwm_a_inst_x.count_q\[2\] dut.pwm_a_inst_x.count_q\[1\]
+ dut.pwm_a_inst_x.count_q\[0\] vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__and4_1
X_1778_ dut.pwm_a_inst_x.count_q\[9\] _0295_ vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__nand2_1
XFILLER_57_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2681_ clknet_leaf_18_clk dut.pwm_a_inst_y.count_d\[4\] net86 vssd1 vssd1 vccd1 vccd1
+ dut.pwm_a_inst_y.count_q\[4\] sky130_fd_sc_hd__dfrtp_2
X_1701_ _1259_ _1268_ _1270_ vssd1 vssd1 vccd1 vccd1 _1271_ sky130_fd_sc_hd__or3_1
X_2750_ clknet_leaf_27_clk _0135_ net75 vssd1 vssd1 vccd1 vccd1 dut.actual_duty_x\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1563_ dut.pwm_a_inst_y.count_q\[12\] _1040_ vssd1 vssd1 vccd1 vccd1 _1152_ sky130_fd_sc_hd__nand2_1
X_1632_ dut.pwm_a_inst_y.count_q\[1\] dut.pwm_a_inst_y.count_q\[0\] dut.pwm_a_inst_y.count_q\[2\]
+ vssd1 vssd1 vccd1 vccd1 _1218_ sky130_fd_sc_hd__a21o_1
X_1494_ net37 _1078_ _1048_ vssd1 vssd1 vccd1 vccd1 _1083_ sky130_fd_sc_hd__a21o_1
X_2115_ dut.spi.shift_reg_q\[6\] net20 _0520_ net228 _0527_ vssd1 vssd1 vccd1 vccd1
+ _0107_ sky130_fd_sc_hd__o221a_1
XFILLER_39_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout38 dut.actual_duty_y\[5\] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__buf_2
Xfanout27 _0355_ vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_2
X_2046_ _0019_ _0480_ vssd1 vssd1 vccd1 vccd1 _0481_ sky130_fd_sc_hd__nor2_1
Xfanout49 dut.actual_duty_x\[3\] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__buf_2
XFILLER_13_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2879_ clknet_leaf_1_clk _0016_ net53 vssd1 vssd1 vccd1 vccd1 dut.clkdiv_inst.counter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_9_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout69_A net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload19 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 clkload19/Y sky130_fd_sc_hd__clkinv_4
XFILLER_48_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2664_ clknet_leaf_9_clk _0027_ net70 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_500hz\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2802_ clknet_leaf_8_clk _0156_ net64 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_200ms\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_2733_ clknet_leaf_5_clk _0074_ net63 vssd1 vssd1 vccd1 vccd1 dut.microstep_y.ctr\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2092__S dut.clk_en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1615_ _1157_ _1158_ _1162_ _1203_ vssd1 vssd1 vccd1 vccd1 _1204_ sky130_fd_sc_hd__o211a_1
X_1546_ _0915_ net42 _1121_ _1132_ vssd1 vssd1 vccd1 vccd1 _1135_ sky130_fd_sc_hd__and4_1
X_1477_ _1045_ _1065_ net36 vssd1 vssd1 vccd1 vccd1 _1066_ sky130_fd_sc_hd__a21oi_1
XFILLER_5_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2595_ dut.ir_sensor_array.final_sensor_data\[3\] dut.ir_sensor_array.final_sensor_data\[2\]
+ _0891_ net2 _0928_ vssd1 vssd1 vccd1 vccd1 _0892_ sky130_fd_sc_hd__o311a_1
XFILLER_42_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2029_ _0470_ _0471_ vssd1 vssd1 vccd1 vccd1 _0056_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_17_Left_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1400_ dut.lcd1602.cnt_200ms\[6\] _1003_ vssd1 vssd1 vccd1 vccd1 _1004_ sky130_fd_sc_hd__and2_1
X_2380_ dut.lcd1602.cnt_200ms\[9\] _0748_ vssd1 vssd1 vccd1 vccd1 _0751_ sky130_fd_sc_hd__or2_1
X_1331_ dut.microstep_y.ctr\[14\] dut.microstep_y.ctr\[15\] dut.microstep_y.ctr\[17\]
+ dut.microstep_y.ctr\[16\] vssd1 vssd1 vccd1 vccd1 _0952_ sky130_fd_sc_hd__nand4b_1
XFILLER_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2647_ clknet_leaf_13_clk _0118_ vssd1 vssd1 vccd1 vccd1 dut.data_in\[1\] sky130_fd_sc_hd__dfxtp_1
X_2716_ clknet_leaf_20_clk net122 net76 vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_x.count_q\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1529_ _1111_ _1113_ vssd1 vssd1 vccd1 vccd1 _1118_ sky130_fd_sc_hd__and2_1
X_2578_ dut.ir_sensor_array.final_sensor_data\[14\] _0875_ dut.ir_sensor_array.final_sensor_data\[13\]
+ vssd1 vssd1 vccd1 vccd1 _0876_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_25_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_2_Left_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1880_ dut.pwm_a_inst_x.count_q\[15\] _0380_ net26 vssd1 vssd1 vccd1 vccd1 _0382_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_14_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2501_ dut.microstep_y.clk_en _0816_ net36 vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__a21o_1
X_1314_ _0934_ _0937_ vssd1 vssd1 vccd1 vccd1 _0938_ sky130_fd_sc_hd__nand2_2
X_2363_ dut.lcd1602.cnt_200ms\[0\] dut.lcd1602.cnt_200ms\[1\] net251 vssd1 vssd1 vccd1
+ vccd1 _0741_ sky130_fd_sc_hd__a21oi_1
XFILLER_44_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2432_ _0780_ _0782_ _0779_ vssd1 vssd1 vccd1 vccd1 _0784_ sky130_fd_sc_hd__a21boi_1
X_2294_ _0681_ vssd1 vssd1 vccd1 vccd1 _0682_ sky130_fd_sc_hd__inv_2
XFILLER_64_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1932_ _0412_ _0413_ vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__nor2_1
X_1863_ _0371_ net26 _0370_ vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_x.count_d\[8\]
+ sky130_fd_sc_hd__and3b_1
X_2415_ dut.ball_pos_x\[2\] _0502_ _0508_ vssd1 vssd1 vccd1 vccd1 _0767_ sky130_fd_sc_hd__nand3_1
X_1794_ dut.pwm_a_inst_x.count_q\[9\] _0295_ vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__or2_1
Xteam_02_119 vssd1 vssd1 vccd1 vccd1 team_02_119/HI gpio_out[31] sky130_fd_sc_hd__conb_1
Xteam_02_108 vssd1 vssd1 vccd1 vccd1 team_02_108/HI gpio_out[20] sky130_fd_sc_hd__conb_1
XFILLER_29_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2277_ dut.pid_x.x_pid.last_error\[1\] _0506_ dut.pid_x.x_pid.last_error\[3\] vssd1
+ vssd1 vccd1 vccd1 _0665_ sky130_fd_sc_hd__a21oi_1
X_2346_ _0683_ _0722_ vssd1 vssd1 vccd1 vccd1 _0731_ sky130_fd_sc_hd__nor2_1
XFILLER_37_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_50_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_23_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_5_Left_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2131_ net20 _0536_ _0535_ _0514_ vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__o211a_1
X_2200_ _0573_ _0585_ vssd1 vssd1 vccd1 vccd1 _0603_ sky130_fd_sc_hd__or2_1
X_2062_ dut.clkdiv_inst.counter\[13\] _0487_ net287 vssd1 vssd1 vccd1 vccd1 _0490_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_34_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_14_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1915_ net269 _0400_ vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__nor2_1
X_1777_ dut.pwm_a_inst_x.count_q\[7\] _0294_ dut.pwm_a_inst_x.count_q\[8\] vssd1 vssd1
+ vccd1 vccd1 _0295_ sky130_fd_sc_hd__o21a_1
X_1846_ net27 _0359_ _0360_ vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_x.count_d\[2\]
+ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_15_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2329_ net46 _0701_ vssd1 vssd1 vccd1 vccd1 _0717_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_63_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_31_Left_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2680_ clknet_leaf_18_clk dut.pwm_a_inst_y.count_d\[3\] net79 vssd1 vssd1 vccd1 vccd1
+ dut.pwm_a_inst_y.count_q\[3\] sky130_fd_sc_hd__dfrtp_1
X_1631_ dut.pwm_a_inst_y.count_q\[2\] dut.pwm_a_inst_y.count_q\[1\] dut.pwm_a_inst_y.count_q\[0\]
+ vssd1 vssd1 vccd1 vccd1 _1217_ sky130_fd_sc_hd__nand3_1
XFILLER_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1700_ _1253_ _1269_ vssd1 vssd1 vccd1 vccd1 _1270_ sky130_fd_sc_hd__nand2_1
X_1562_ _1148_ _1150_ _1042_ _1146_ vssd1 vssd1 vccd1 vccd1 _1151_ sky130_fd_sc_hd__o2bb2a_1
X_1493_ _1077_ _1081_ vssd1 vssd1 vccd1 vccd1 _1082_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_3_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_54_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2114_ dut.data_in\[7\] _0515_ vssd1 vssd1 vccd1 vccd1 _0527_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_2_2__f_clk_X clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2045_ dut.clkdiv_inst.counter\[7\] _0478_ vssd1 vssd1 vccd1 vccd1 _0480_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_60_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout39 dut.actual_duty_y\[4\] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__buf_2
XFILLER_13_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout28 _0944_ vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__buf_2
X_1829_ _0292_ _0300_ _0305_ _0346_ _0306_ vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_9_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2878_ clknet_leaf_1_clk _0015_ net53 vssd1 vssd1 vccd1 vccd1 dut.clkdiv_inst.counter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2863__RESET_B net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2801_ clknet_leaf_8_clk _0155_ net66 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_200ms\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2663_ clknet_leaf_9_clk _0026_ net70 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_500hz\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1614_ _1141_ _1159_ _1161_ _1167_ _1202_ vssd1 vssd1 vccd1 vccd1 _1203_ sky130_fd_sc_hd__a311o_1
X_2732_ clknet_leaf_5_clk _0073_ net67 vssd1 vssd1 vccd1 vccd1 dut.microstep_y.ctr\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2594_ dut.ir_sensor_array.final_sensor_data\[6\] dut.ir_sensor_array.final_sensor_data\[7\]
+ _0868_ vssd1 vssd1 vccd1 vccd1 _0891_ sky130_fd_sc_hd__o21a_1
X_1545_ dut.actual_duty_y\[1\] net42 vssd1 vssd1 vccd1 vccd1 _1134_ sky130_fd_sc_hd__nand2_1
X_1476_ dut.actual_duty_y\[5\] dut.actual_duty_y\[6\] vssd1 vssd1 vccd1 vccd1 _1065_
+ sky130_fd_sc_hd__or2_1
XFILLER_5_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2028_ dut.microstep_x.ctr\[28\] _0469_ vssd1 vssd1 vccd1 vccd1 _0471_ sky130_fd_sc_hd__nand2_1
XFILLER_50_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1330_ dut.microstep_y.ctr\[19\] dut.microstep_y.ctr\[18\] dut.microstep_y.ctr\[21\]
+ dut.microstep_y.ctr\[20\] vssd1 vssd1 vccd1 vccd1 _0951_ sky130_fd_sc_hd__or4_1
XFILLER_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2646_ clknet_leaf_14_clk _0117_ vssd1 vssd1 vccd1 vccd1 dut.data_in\[0\] sky130_fd_sc_hd__dfxtp_1
X_2715_ clknet_leaf_20_clk net123 net76 vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_x.count_q\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_2577_ net2 _0874_ dut.ir_sensor_array.final_sensor_data\[15\] vssd1 vssd1 vccd1
+ vccd1 _0875_ sky130_fd_sc_hd__a21oi_1
X_1528_ _1115_ _1116_ vssd1 vssd1 vccd1 vccd1 _1117_ sky130_fd_sc_hd__nand2_1
X_1459_ net38 net39 vssd1 vssd1 vccd1 vccd1 _1048_ sky130_fd_sc_hd__and2_1
XFILLER_42_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2431_ _0781_ _0782_ vssd1 vssd1 vccd1 vccd1 _0783_ sky130_fd_sc_hd__xnor2_1
X_2500_ net37 dut.microstep_y.clk_en _0812_ _0845_ vssd1 vssd1 vccd1 vccd1 _0174_
+ sky130_fd_sc_hd__o22a_1
X_1313_ dut.lcd1602.cnt_500hz\[13\] _0936_ dut.lcd1602.cnt_500hz\[10\] dut.lcd1602.cnt_500hz\[14\]
+ vssd1 vssd1 vccd1 vccd1 _0937_ sky130_fd_sc_hd__and4b_1
X_2362_ net13 net260 vssd1 vssd1 vccd1 vccd1 _0141_ sky130_fd_sc_hd__nand2_1
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2293_ _0679_ _0680_ vssd1 vssd1 vccd1 vccd1 _0681_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_47_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2629_ clknet_leaf_14_clk net162 net81 vssd1 vssd1 vccd1 vccd1 dut.spi.shift_reg_q\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1931_ dut.microstep_y.ctr\[17\] dut.microstep_y.ctr\[18\] _0409_ vssd1 vssd1 vccd1
+ vccd1 _0413_ sky130_fd_sc_hd__and3_1
X_1793_ _0286_ _0310_ vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__and2_1
X_1862_ dut.pwm_a_inst_x.count_q\[8\] dut.pwm_a_inst_x.count_q\[7\] _0367_ vssd1 vssd1
+ vccd1 vccd1 _0371_ sky130_fd_sc_hd__and3_1
X_2414_ dut.ball_pos_x\[2\] _0502_ _0508_ vssd1 vssd1 vccd1 vccd1 _0766_ sky130_fd_sc_hd__and3_1
Xteam_02_109 vssd1 vssd1 vccd1 vccd1 team_02_109/HI gpio_out[21] sky130_fd_sc_hd__conb_1
X_2345_ dut.actual_duty_x\[2\] _0930_ _0729_ _0730_ vssd1 vssd1 vccd1 vccd1 _0134_
+ sky130_fd_sc_hd__a22o_1
X_2276_ dut.pid_x.x_pid.last_error\[2\] _0512_ vssd1 vssd1 vccd1 vccd1 _0664_ sky130_fd_sc_hd__xnor2_1
XFILLER_52_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_50_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_44_Left_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2130_ dut.spi.bit_counter_q\[0\] dut.spi.bit_counter_q\[1\] vssd1 vssd1 vccd1 vccd1
+ _0536_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_53_Left_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2061_ dut.clkdiv_inst.counter\[13\] dut.clkdiv_inst.counter\[14\] _0487_ vssd1 vssd1
+ vccd1 vccd1 _0489_ sky130_fd_sc_hd__and3_1
XFILLER_19_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1914_ dut.microstep_y.ctr\[11\] dut.microstep_y.ctr\[12\] _0398_ vssd1 vssd1 vccd1
+ vccd1 _0402_ sky130_fd_sc_hd__and3_1
XFILLER_34_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_62_Left_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1776_ dut.pwm_a_inst_x.count_q\[6\] dut.pwm_a_inst_x.count_q\[5\] dut.pwm_a_inst_x.count_q\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__or3_1
X_1845_ dut.pwm_a_inst_x.count_q\[1\] dut.pwm_a_inst_x.count_q\[0\] dut.pwm_a_inst_x.count_q\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0360_ sky130_fd_sc_hd__a21o_1
X_2328_ net11 _0705_ _0713_ _0677_ _0715_ vssd1 vssd1 vccd1 vccd1 _0716_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_55_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2259_ dut.ir_sensor_array.bit_count\[0\] net35 dut.ir_sensor_array.state\[1\] vssd1
+ vssd1 vccd1 vccd1 _0653_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_63_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1630_ net318 dut.pwm_a_inst_y.count_q\[0\] _1216_ vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_y.count_d\[1\]
+ sky130_fd_sc_hd__a21oi_1
X_1561_ _1038_ _1149_ _1040_ vssd1 vssd1 vccd1 vccd1 _1150_ sky130_fd_sc_hd__a21bo_1
X_1492_ _0916_ _1080_ vssd1 vssd1 vccd1 vccd1 _1081_ sky130_fd_sc_hd__or2_1
XFILLER_3_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2113_ net219 net20 _0520_ net242 _0526_ vssd1 vssd1 vccd1 vccd1 _0106_ sky130_fd_sc_hd__o221a_1
X_2044_ _0478_ _0479_ vssd1 vssd1 vccd1 vccd1 _0015_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_60_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout18 dut.lcd1602.lcd_ctrl vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_4
XFILLER_30_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2877_ clknet_leaf_0_clk _0014_ net53 vssd1 vssd1 vccd1 vccd1 dut.clkdiv_inst.counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_1828_ _0307_ _0309_ _0345_ vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__o21a_1
X_1759_ _0274_ _0276_ vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__nand2_1
XFILLER_38_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_14_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2800_ clknet_leaf_8_clk _0154_ net64 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_200ms\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2731_ clknet_leaf_5_clk _0072_ net63 vssd1 vssd1 vccd1 vccd1 dut.microstep_y.ctr\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_2662_ clknet_leaf_9_clk _0020_ net70 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_500hz\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1613_ _1170_ _1172_ _1200_ _1201_ _1168_ vssd1 vssd1 vccd1 vccd1 _1202_ sky130_fd_sc_hd__o221a_1
X_1544_ _0916_ _0917_ vssd1 vssd1 vccd1 vccd1 _1133_ sky130_fd_sc_hd__nor2_1
X_2593_ dut.ball_pos_x\[0\] _0944_ _0862_ _0890_ vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__a22o_1
XFILLER_5_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_29_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1475_ _1057_ _1063_ vssd1 vssd1 vccd1 vccd1 _1064_ sky130_fd_sc_hd__nand2_1
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2027_ dut.microstep_x.ctr\[28\] _0469_ vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__or2_1
XFILLER_40_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2714_ clknet_leaf_20_clk dut.pwm_a_inst_x.count_d\[17\] net76 vssd1 vssd1 vccd1
+ vccd1 dut.pwm_a_inst_x.count_q\[17\] sky130_fd_sc_hd__dfrtp_1
X_2645_ clknet_leaf_15_clk _0116_ net82 vssd1 vssd1 vccd1 vccd1 dut.spi.bit_counter_q\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1527_ _1107_ _1114_ vssd1 vssd1 vccd1 vccd1 _1116_ sky130_fd_sc_hd__or2_1
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2576_ dut.ir_sensor_array.final_sensor_data\[2\] _0873_ _0928_ vssd1 vssd1 vccd1
+ vccd1 _0874_ sky130_fd_sc_hd__o21ai_1
X_1389_ dut.spi.cs_low_counter_q\[1\] dut.spi.cs_low_counter_q\[0\] dut.spi.cs_low_counter_q\[3\]
+ dut.spi.cs_low_counter_q\[2\] vssd1 vssd1 vccd1 vccd1 _0996_ sky130_fd_sc_hd__and4_1
X_1458_ _1043_ _1045_ vssd1 vssd1 vccd1 vccd1 _1047_ sky130_fd_sc_hd__or2_1
XFILLER_35_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2361_ dut.lcd1602.cnt_200ms\[0\] net259 vssd1 vssd1 vccd1 vccd1 _0740_ sky130_fd_sc_hd__xnor2_1
X_2430_ dut.pid_y.y_pid.last_error\[2\] _0924_ _0772_ vssd1 vssd1 vccd1 vccd1 _0782_
+ sky130_fd_sc_hd__o21a_1
X_1312_ dut.lcd1602.cnt_500hz\[11\] dut.lcd1602.cnt_500hz\[12\] _0935_ vssd1 vssd1
+ vccd1 vccd1 _0936_ sky130_fd_sc_hd__and3_1
XFILLER_1_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2292_ dut.actual_duty_x\[4\] _0678_ vssd1 vssd1 vccd1 vccd1 _0680_ sky130_fd_sc_hd__nand2_1
XFILLER_64_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2559_ dut.ir_sensor_array.final_sensor_data\[24\] net323 _0943_ vssd1 vssd1 vccd1
+ vccd1 _0207_ sky130_fd_sc_hd__mux2_1
X_2628_ clknet_leaf_24_clk _0099_ net73 vssd1 vssd1 vccd1 vccd1 dut.pid_x.x_pid.last_error\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xmax_cap15 net16 vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__buf_1
XFILLER_62_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1930_ dut.microstep_y.ctr\[17\] _0409_ net257 vssd1 vssd1 vccd1 vccd1 _0412_ sky130_fd_sc_hd__a21oi_1
X_1792_ _1273_ _0235_ _0285_ vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__nand3_1
XFILLER_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1861_ dut.pwm_a_inst_x.count_q\[7\] dut.pwm_a_inst_x.count_q\[6\] _0366_ dut.pwm_a_inst_x.count_q\[8\]
+ vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__a31o_1
X_2413_ dut.lcd1602.currentState\[5\] _0577_ net18 vssd1 vssd1 vccd1 vccd1 _0167_
+ sky130_fd_sc_hd__mux2_1
X_2344_ _0331_ _0719_ _0930_ vssd1 vssd1 vccd1 vccd1 _0730_ sky130_fd_sc_hd__a21oi_1
X_2275_ net193 _0662_ net28 vssd1 vssd1 vccd1 vccd1 _0131_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_58_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2695__125 vssd1 vssd1 vccd1 vccd1 _2695__125/HI net125 sky130_fd_sc_hd__conb_1
XFILLER_47_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2060_ net244 _0487_ vssd1 vssd1 vccd1 vccd1 _0006_ sky130_fd_sc_hd__xor2_1
XFILLER_19_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2962_ dut.sclk_lcd vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
X_1913_ net304 _0398_ _0401_ vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__o21a_1
XFILLER_8_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1775_ dut.pwm_a_inst_x.count_q\[5\] dut.pwm_a_inst_x.count_q\[4\] vssd1 vssd1 vccd1
+ vccd1 _0293_ sky130_fd_sc_hd__nor2_1
X_1844_ dut.pwm_a_inst_x.count_q\[2\] dut.pwm_a_inst_x.count_q\[1\] dut.pwm_a_inst_x.count_q\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__nand3_1
XFILLER_57_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2258_ net168 net19 net81 _0652_ vssd1 vssd1 vccd1 vccd1 _0125_ sky130_fd_sc_hd__o211a_1
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2327_ _0683_ _0711_ _0713_ _0677_ _0712_ vssd1 vssd1 vccd1 vccd1 _0715_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_63_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2189_ net12 _0570_ vssd1 vssd1 vccd1 vccd1 _0592_ sky130_fd_sc_hd__nand2_1
XFILLER_43_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1560_ dut.pwm_a_inst_y.count_q\[10\] dut.pwm_a_inst_y.count_q\[11\] dut.pwm_a_inst_y.count_q\[9\]
+ vssd1 vssd1 vccd1 vccd1 _1149_ sky130_fd_sc_hd__and3_1
X_2112_ dut.data_in\[6\] _0515_ vssd1 vssd1 vccd1 vccd1 _0526_ sky130_fd_sc_hd__or2_1
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1491_ net37 _1079_ vssd1 vssd1 vccd1 vccd1 _1080_ sky130_fd_sc_hd__xor2_1
XFILLER_3_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout19 dut.lcd1602.lcd_ctrl vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_2
X_2043_ dut.clkdiv_inst.counter\[5\] _0476_ net295 vssd1 vssd1 vccd1 vccd1 _0479_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_17_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1827_ _0307_ _0309_ _0311_ _0313_ _0344_ vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__a221o_1
X_2876_ clknet_leaf_0_clk _0013_ net53 vssd1 vssd1 vccd1 vccd1 dut.clkdiv_inst.counter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1689_ net49 _1251_ vssd1 vssd1 vccd1 vccd1 _1259_ sky130_fd_sc_hd__xnor2_1
X_1758_ net49 _0275_ vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__and2b_1
XFILLER_57_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2661_ clknet_leaf_14_clk net19 net81 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.out_valid
+ sky130_fd_sc_hd__dfrtp_1
X_2730_ clknet_leaf_6_clk _0071_ net63 vssd1 vssd1 vccd1 vccd1 dut.microstep_y.ctr\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_1612_ _1170_ _1172_ _1174_ _1175_ vssd1 vssd1 vccd1 vccd1 _1201_ sky130_fd_sc_hd__a22o_1
X_1543_ _1130_ _1131_ vssd1 vssd1 vccd1 vccd1 _1132_ sky130_fd_sc_hd__xor2_1
X_2592_ dut.ir_sensor_array.final_sensor_data\[34\] _0889_ _0926_ vssd1 vssd1 vccd1
+ vccd1 _0890_ sky130_fd_sc_hd__o21ai_1
X_1474_ _1046_ _1056_ dut.actual_duty_y\[3\] vssd1 vssd1 vccd1 vccd1 _1063_ sky130_fd_sc_hd__a21o_1
XFILLER_54_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2026_ _0468_ _0469_ vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__nor2_1
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2859_ clknet_leaf_2_clk _0212_ net59 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_20_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout67_A net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_2_3__f_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2644_ clknet_leaf_15_clk _0115_ net84 vssd1 vssd1 vccd1 vccd1 dut.spi.bit_counter_q\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2713_ clknet_leaf_21_clk dut.pwm_a_inst_x.count_d\[16\] net76 vssd1 vssd1 vccd1
+ vccd1 dut.pwm_a_inst_x.count_q\[16\] sky130_fd_sc_hd__dfrtp_1
X_1526_ _1107_ _1114_ vssd1 vssd1 vccd1 vccd1 _1115_ sky130_fd_sc_hd__nand2_1
X_1457_ net36 net37 vssd1 vssd1 vccd1 vccd1 _1046_ sky130_fd_sc_hd__nand2_1
X_2575_ dut.ir_sensor_array.final_sensor_data\[4\] _0872_ dut.ir_sensor_array.final_sensor_data\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0873_ sky130_fd_sc_hd__o21ba_1
X_1388_ dut.spi.cs_low_counter_q\[1\] dut.spi.cs_low_counter_q\[0\] dut.spi.cs_low_counter_q\[2\]
+ dut.spi.cs_low_counter_q\[3\] vssd1 vssd1 vccd1 vccd1 _0995_ sky130_fd_sc_hd__a31o_1
XFILLER_35_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2009_ net206 _0459_ vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__xor2_1
XANTENNA_clkbuf_leaf_13_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_28_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1311_ dut.lcd1602.cnt_500hz\[6\] dut.lcd1602.cnt_500hz\[9\] dut.lcd1602.cnt_500hz\[8\]
+ dut.lcd1602.cnt_500hz\[7\] vssd1 vssd1 vccd1 vccd1 _0935_ sky130_fd_sc_hd__and4bb_1
X_2360_ net183 net13 vssd1 vssd1 vccd1 vccd1 _0140_ sky130_fd_sc_hd__nand2_1
X_2291_ dut.actual_duty_x\[4\] _0678_ vssd1 vssd1 vccd1 vccd1 _0679_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2627_ clknet_leaf_19_clk _0098_ net73 vssd1 vssd1 vccd1 vccd1 dut.pid_x.x_pid.last_error\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1509_ _0917_ _1097_ vssd1 vssd1 vccd1 vccd1 _1098_ sky130_fd_sc_hd__or2_1
X_2489_ _0790_ _0813_ _0833_ _1186_ net44 vssd1 vssd1 vccd1 vccd1 _0839_ sky130_fd_sc_hd__o221a_1
X_2558_ dut.ir_sensor_array.final_sensor_data\[24\] net317 net31 vssd1 vssd1 vccd1
+ vccd1 _0206_ sky130_fd_sc_hd__mux2_1
XFILLER_46_48 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xmax_cap16 _0035_ vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__buf_1
XFILLER_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1860_ net303 _0367_ _0369_ vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_x.count_d\[7\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_14_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_26_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1791_ _0287_ _0308_ vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__nor2_1
X_2412_ dut.lcd1602.currentState\[4\] _0582_ net18 vssd1 vssd1 vccd1 vccd1 _0166_
+ sky130_fd_sc_hd__mux2_1
X_2343_ _0685_ _0722_ _0728_ vssd1 vssd1 vccd1 vccd1 _0729_ sky130_fd_sc_hd__a21o_1
X_2274_ _0662_ _0663_ vssd1 vssd1 vccd1 vccd1 _0130_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_17_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_37_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1989_ _0446_ _0447_ vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__nor2_1
XFILLER_20_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2961_ dut.sdo_lcd vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
X_1912_ net17 _0400_ vssd1 vssd1 vccd1 vccd1 _0401_ sky130_fd_sc_hd__nor2_1
X_1843_ net240 dut.pwm_a_inst_x.count_q\[0\] _0358_ vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_x.count_d\[1\]
+ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_6_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1774_ net45 _0290_ _0291_ vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__o21ba_1
X_2257_ _0603_ _0627_ _0642_ _0938_ vssd1 vssd1 vccd1 vccd1 _0652_ sky130_fd_sc_hd__a31o_1
X_2326_ _0713_ vssd1 vssd1 vccd1 vccd1 _0714_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_63_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2188_ net12 _0570_ vssd1 vssd1 vccd1 vccd1 _0591_ sky130_fd_sc_hd__and2_1
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1490_ _1048_ _1078_ vssd1 vssd1 vccd1 vccd1 _1079_ sky130_fd_sc_hd__nand2b_1
XFILLER_3_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1 dut.lcd1602.cnt_200ms\[21\] vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__dlygate4sd3_1
X_2111_ net216 net20 _0520_ net219 _0525_ vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__o221a_1
XFILLER_39_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2042_ dut.clkdiv_inst.counter\[5\] dut.clkdiv_inst.counter\[6\] _0476_ vssd1 vssd1
+ vccd1 vccd1 _0478_ sky130_fd_sc_hd__and3_1
XFILLER_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2875_ clknet_leaf_0_clk _0012_ net54 vssd1 vssd1 vccd1 vccd1 dut.clkdiv_inst.counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1826_ _0311_ _0313_ _0317_ _0343_ _0318_ vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1688_ _1253_ _1256_ vssd1 vssd1 vccd1 vccd1 _1258_ sky130_fd_sc_hd__xor2_1
X_1757_ _0920_ _0268_ vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__nor2_1
XFILLER_57_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2309_ _0677_ _0681_ _0696_ net11 _0693_ vssd1 vssd1 vccd1 vccd1 _0697_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1611_ _1174_ _1175_ _1198_ _1199_ _1179_ vssd1 vssd1 vccd1 vccd1 _1200_ sky130_fd_sc_hd__o221a_1
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2660_ clknet_leaf_25_clk _0131_ net60 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.bit_count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_1473_ _1053_ _1061_ vssd1 vssd1 vccd1 vccd1 _1062_ sky130_fd_sc_hd__nor2_1
X_1542_ _0915_ net42 _1123_ _1108_ dut.actual_duty_y\[1\] vssd1 vssd1 vccd1 vccd1
+ _1131_ sky130_fd_sc_hd__a32o_1
X_2591_ dut.ir_sensor_array.final_sensor_data\[36\] _0888_ dut.ir_sensor_array.final_sensor_data\[35\]
+ vssd1 vssd1 vccd1 vccd1 _0889_ sky130_fd_sc_hd__o21ba_1
XFILLER_54_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2025_ dut.microstep_x.ctr\[27\] dut.microstep_x.ctr\[26\] _0467_ vssd1 vssd1 vccd1
+ vccd1 _0469_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_59_Left_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2789_ clknet_leaf_9_clk _0143_ net65 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_200ms\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_2858_ clknet_leaf_2_clk _0211_ net55 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_1809_ dut.pwm_a_inst_x.count_q\[5\] dut.pwm_a_inst_x.count_q\[4\] vssd1 vssd1 vccd1
+ vccd1 _0327_ sky130_fd_sc_hd__and2_1
XFILLER_41_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2643_ clknet_leaf_15_clk _0114_ net82 vssd1 vssd1 vccd1 vccd1 dut.spi.bit_counter_q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2712_ clknet_leaf_20_clk dut.pwm_a_inst_x.count_d\[15\] net76 vssd1 vssd1 vccd1
+ vccd1 dut.pwm_a_inst_x.count_q\[15\] sky130_fd_sc_hd__dfrtp_1
X_2574_ _0927_ dut.ir_sensor_array.final_sensor_data\[7\] dut.ir_sensor_array.final_sensor_data\[5\]
+ vssd1 vssd1 vccd1 vccd1 _0872_ sky130_fd_sc_hd__a21oi_1
X_1387_ _0991_ _0993_ _0994_ vssd1 vssd1 vccd1 vccd1 dut.spi.cs_low_counter_d\[2\]
+ sky130_fd_sc_hd__and3_1
X_1525_ _1111_ _1113_ vssd1 vssd1 vccd1 vccd1 _1114_ sky130_fd_sc_hd__nor2_1
X_1456_ net38 net37 vssd1 vssd1 vccd1 vccd1 _1045_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_25_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2008_ _0458_ _0459_ vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__nor2_1
XFILLER_51_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1310_ dut.lcd1602.cnt_500hz\[5\] dut.lcd1602.cnt_500hz\[4\] _0933_ vssd1 vssd1 vccd1
+ vccd1 _0934_ sky130_fd_sc_hd__and3_1
XFILLER_49_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_22_Left_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2290_ _0255_ _0268_ vssd1 vssd1 vccd1 vccd1 _0678_ sky130_fd_sc_hd__nand2_1
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2626_ clknet_leaf_24_clk _0097_ net73 vssd1 vssd1 vccd1 vccd1 dut.pid_x.x_pid.last_error\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2557_ net317 dut.ir_sensor_array.final_sensor_data\[22\] net31 vssd1 vssd1 vccd1
+ vccd1 _0205_ sky130_fd_sc_hd__mux2_1
XFILLER_55_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1439_ dut.lcd1602.cnt_500hz\[11\] _1028_ dut.lcd1602.cnt_500hz\[12\] vssd1 vssd1
+ vccd1 vccd1 _1031_ sky130_fd_sc_hd__a21o_1
Xmax_cap17 _0066_ vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_2
X_1508_ net38 _1096_ vssd1 vssd1 vccd1 vccd1 _1097_ sky130_fd_sc_hd__xor2_1
X_2488_ _0787_ _0834_ vssd1 vssd1 vccd1 vccd1 _0838_ sky130_fd_sc_hd__or2_1
XFILLER_62_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1790_ _1258_ _1271_ _0286_ vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__and3_1
X_2411_ dut.lcd1602.currentState\[3\] _0553_ net18 vssd1 vssd1 vccd1 vccd1 _0165_
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2342_ net11 _0722_ _0719_ vssd1 vssd1 vccd1 vccd1 _0728_ sky130_fd_sc_hd__o21bai_1
X_2273_ net297 _0660_ net28 vssd1 vssd1 vccd1 vccd1 _0663_ sky130_fd_sc_hd__o21ai_1
XFILLER_60_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_12_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1988_ net278 _0444_ vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__nor2_1
XFILLER_20_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2609_ _0850_ _0904_ net30 vssd1 vssd1 vccd1 vccd1 _0905_ sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_leaf_27_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_2__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_41_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2960_ dut.cs_n_lcd vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
X_1911_ dut.microstep_y.ctr\[11\] _0398_ vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__and2_1
X_1842_ dut.pwm_a_inst_x.count_q\[1\] dut.pwm_a_inst_x.count_q\[0\] net27 vssd1 vssd1
+ vccd1 vccd1 _0358_ sky130_fd_sc_hd__o21ai_1
X_1773_ net45 _0290_ _0288_ vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__a21bo_1
X_2256_ net81 _0651_ vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__and2_1
X_2187_ _0554_ _0583_ vssd1 vssd1 vccd1 vccd1 _0590_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_40_Left_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_25_Left_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2325_ net48 _0700_ vssd1 vssd1 vccd1 vccd1 _0713_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_63_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2110_ dut.data_in\[5\] _0515_ vssd1 vssd1 vccd1 vccd1 _0525_ sky130_fd_sc_hd__or2_1
Xhold2 dut.ir_sensor_array.state\[0\] vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__dlygate4sd3_1
X_2041_ net281 _0476_ vssd1 vssd1 vccd1 vccd1 _0014_ sky130_fd_sc_hd__xor2_1
X_1825_ _0320_ _0321_ _0342_ vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__a21o_1
X_1756_ _0272_ _0273_ vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__and2_1
X_2874_ clknet_leaf_0_clk _0011_ net53 vssd1 vssd1 vccd1 vccd1 dut.clkdiv_inst.counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_57_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1687_ _1253_ _1256_ vssd1 vssd1 vccd1 vccd1 _1257_ sky130_fd_sc_hd__and2b_1
X_2308_ _0694_ _0695_ vssd1 vssd1 vccd1 vccd1 _0696_ sky130_fd_sc_hd__nor2_1
XFILLER_57_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2239_ net12 _0625_ _0639_ _0598_ _0616_ vssd1 vssd1 vccd1 vccd1 _0640_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_0_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1610_ _1036_ _1177_ _1178_ _1181_ dut.pwm_a_inst_y.count_q\[4\] vssd1 vssd1 vccd1
+ vccd1 _1199_ sky130_fd_sc_hd__a32o_1
X_2590_ dut.ir_sensor_array.final_sensor_data\[38\] _0887_ dut.ir_sensor_array.final_sensor_data\[37\]
+ vssd1 vssd1 vccd1 vccd1 _0888_ sky130_fd_sc_hd__o21ba_1
X_1541_ _1125_ _1129_ vssd1 vssd1 vccd1 vccd1 _1130_ sky130_fd_sc_hd__nor2_1
X_1472_ _1058_ _1060_ _1046_ vssd1 vssd1 vccd1 vccd1 _1061_ sky130_fd_sc_hd__o21a_1
XFILLER_35_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2024_ dut.microstep_x.ctr\[26\] _0467_ net233 vssd1 vssd1 vccd1 vccd1 _0468_ sky130_fd_sc_hd__a21oi_1
X_2857_ clknet_leaf_2_clk _0210_ net55 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2788_ clknet_leaf_11_clk _0142_ net70 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_200ms\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1739_ dut.actual_duty_x\[1\] _0256_ _0254_ vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__a21oi_1
X_1808_ _0280_ _0325_ vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__nor2_1
XFILLER_58_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2711_ clknet_leaf_20_clk dut.pwm_a_inst_x.count_d\[14\] net76 vssd1 vssd1 vccd1
+ vccd1 dut.pwm_a_inst_x.count_q\[14\] sky130_fd_sc_hd__dfrtp_1
X_2642_ clknet_leaf_14_clk _0113_ net83 vssd1 vssd1 vccd1 vccd1 dut.spi.bit_counter_q\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1524_ _1098_ _1112_ vssd1 vssd1 vccd1 vccd1 _1113_ sky130_fd_sc_hd__nand2_1
X_2573_ net286 dut.ir_sensor_array.final_sensor_data\[38\] net33 vssd1 vssd1 vccd1
+ vccd1 _0221_ sky130_fd_sc_hd__mux2_1
X_1386_ dut.spi.cs_low_counter_q\[1\] dut.spi.cs_low_counter_q\[0\] dut.spi.cs_low_counter_q\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0994_ sky130_fd_sc_hd__a21o_1
X_1455_ net38 net37 vssd1 vssd1 vccd1 vccd1 _1044_ sky130_fd_sc_hd__and2_1
X_2716__122 vssd1 vssd1 vccd1 vccd1 _2716__122/HI net122 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_25_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2007_ dut.microstep_x.ctr\[19\] _0457_ vssd1 vssd1 vccd1 vccd1 _0459_ sky130_fd_sc_hd__and2_1
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout72_A dut.clkdiv_inst.reset_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2625_ clknet_leaf_15_clk net290 net85 vssd1 vssd1 vccd1 vccd1 dut.spi.clk_counter_q\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_1507_ _1094_ _1095_ vssd1 vssd1 vccd1 vccd1 _1096_ sky130_fd_sc_hd__nand2_1
X_2487_ dut.actual_duty_y\[1\] _0931_ _0836_ _0837_ vssd1 vssd1 vccd1 vccd1 _0169_
+ sky130_fd_sc_hd__a22o_1
X_2556_ dut.ir_sensor_array.final_sensor_data\[22\] net321 net31 vssd1 vssd1 vccd1
+ vccd1 _0204_ sky130_fd_sc_hd__mux2_1
X_1369_ _0977_ _0982_ vssd1 vssd1 vccd1 vccd1 _0983_ sky130_fd_sc_hd__nor2_1
XFILLER_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1438_ net312 _1028_ _1030_ vssd1 vssd1 vccd1 vccd1 _0022_ sky130_fd_sc_hd__o21a_1
Xmax_cap29 net30 vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_55_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2410_ net43 _0586_ net18 vssd1 vssd1 vccd1 vccd1 _0164_ sky130_fd_sc_hd__mux2_1
X_2341_ dut.actual_duty_x\[1\] _0727_ dut.microstep_x.clk_en vssd1 vssd1 vccd1 vccd1
+ _0133_ sky130_fd_sc_hd__mux2_1
XFILLER_37_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2272_ dut.ir_sensor_array.bit_count\[4\] _0660_ vssd1 vssd1 vccd1 vccd1 _0662_ sky130_fd_sc_hd__and2_1
X_1987_ dut.microstep_x.ctr\[11\] dut.microstep_x.ctr\[12\] _0442_ vssd1 vssd1 vccd1
+ vccd1 _0446_ sky130_fd_sc_hd__and3_1
XFILLER_20_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2608_ _0848_ _0903_ vssd1 vssd1 vccd1 vccd1 _0904_ sky130_fd_sc_hd__nor2_1
X_2539_ dut.ir_sensor_array.final_sensor_data\[5\] dut.ir_sensor_array.final_sensor_data\[4\]
+ net32 vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout35_A dut.clk_en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1910_ _0398_ _0399_ vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__nor2_1
X_2890_ clknet_leaf_26_clk _0225_ net60 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1841_ dut.pwm_a_inst_x.count_q\[0\] net27 vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_x.count_d\[0\]
+ sky130_fd_sc_hd__and2b_1
X_1772_ _1257_ _0287_ _0289_ vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__o21a_1
XFILLER_6_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2324_ _0331_ _0674_ _0683_ _0711_ _0709_ vssd1 vssd1 vccd1 vccd1 _0712_ sky130_fd_sc_hd__a221o_1
X_2255_ dut.data_in\[7\] _0938_ _0631_ _0650_ vssd1 vssd1 vccd1 vccd1 _0651_ sky130_fd_sc_hd__a22o_1
X_2186_ _0573_ _0582_ _0584_ _0588_ vssd1 vssd1 vccd1 vccd1 _0589_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_25_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2889__Q dut.clk_en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_11_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold3 dut.clkdiv_inst.counter\[0\] vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__dlygate4sd3_1
X_2040_ _0476_ _0477_ vssd1 vssd1 vccd1 vccd1 _0013_ sky130_fd_sc_hd__nor2_1
XFILLER_62_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2873_ clknet_leaf_0_clk _0010_ net50 vssd1 vssd1 vccd1 vccd1 dut.clkdiv_inst.counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_26_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1686_ _1254_ _1255_ vssd1 vssd1 vccd1 vccd1 _1256_ sky130_fd_sc_hd__nor2_1
X_1755_ _0265_ _0271_ vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__nand2_1
X_1824_ _0320_ _0321_ _0340_ _0341_ _0324_ vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__o221a_1
XFILLER_57_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2238_ dut.ball_pos_x\[2\] _0610_ _0632_ dut.ball_pos_y\[2\] _0593_ vssd1 vssd1 vccd1
+ vccd1 _0639_ sky130_fd_sc_hd__a221o_1
X_2307_ net47 _0679_ vssd1 vssd1 vccd1 vccd1 _0695_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_51_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2169_ net12 _0570_ vssd1 vssd1 vccd1 vccd1 _0572_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1540_ _1120_ _1124_ vssd1 vssd1 vccd1 vccd1 _1129_ sky130_fd_sc_hd__nor2_1
XFILLER_5_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_222 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1471_ _1055_ _1057_ vssd1 vssd1 vccd1 vccd1 _1060_ sky130_fd_sc_hd__and2_1
XFILLER_10_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2023_ net215 _0467_ vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__xor2_1
XFILLER_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2856_ clknet_leaf_2_clk _0209_ net63 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_1807_ _0277_ _0279_ vssd1 vssd1 vccd1 vccd1 _0325_ sky130_fd_sc_hd__and2_1
X_1669_ dut.pwm_a_inst_y.count_q\[14\] dut.pwm_a_inst_y.count_q\[15\] _1237_ dut.pwm_a_inst_y.count_q\[16\]
+ vssd1 vssd1 vccd1 vccd1 _1241_ sky130_fd_sc_hd__a31o_1
X_2787_ clknet_leaf_7_clk _0141_ net65 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_200ms\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1738_ _0254_ _0255_ vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_28_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2710_ clknet_leaf_21_clk dut.pwm_a_inst_x.count_d\[13\] net76 vssd1 vssd1 vccd1
+ vccd1 dut.pwm_a_inst_x.count_q\[13\] sky130_fd_sc_hd__dfrtp_2
X_2641_ clknet_leaf_14_clk _0112_ net83 vssd1 vssd1 vccd1 vccd1 dut.spi.state_q\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1454_ net40 dut.actual_duty_y\[7\] vssd1 vssd1 vccd1 vccd1 _1043_ sky130_fd_sc_hd__nand2_1
X_1523_ _0917_ _1097_ vssd1 vssd1 vccd1 vccd1 _1112_ sky130_fd_sc_hd__nand2_1
X_2572_ dut.ir_sensor_array.final_sensor_data\[38\] net319 net34 vssd1 vssd1 vccd1
+ vccd1 _0220_ sky130_fd_sc_hd__mux2_1
XFILLER_4_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1385_ dut.spi.cs_low_counter_q\[1\] dut.spi.cs_low_counter_q\[0\] dut.spi.cs_low_counter_q\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0993_ sky130_fd_sc_hd__nand3_1
XFILLER_55_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2006_ net255 _0457_ vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_33_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2839_ clknet_leaf_26_clk _0192_ net59 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_29_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_17_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2624_ clknet_leaf_16_clk dut.spi.clk_counter_d\[4\] net85 vssd1 vssd1 vccd1 vccd1
+ dut.spi.clk_counter_q\[4\] sky130_fd_sc_hd__dfrtp_1
X_1437_ dut.lcd1602.cnt_500hz\[11\] _1028_ _1019_ vssd1 vssd1 vccd1 vccd1 _1030_ sky130_fd_sc_hd__a21oi_1
X_1506_ net39 dut.actual_duty_y\[3\] vssd1 vssd1 vccd1 vccd1 _1095_ sky130_fd_sc_hd__nand2_1
X_2486_ _1188_ _0833_ _0834_ _0825_ net44 vssd1 vssd1 vccd1 vccd1 _0837_ sky130_fd_sc_hd__o221a_1
X_2555_ net321 dut.ir_sensor_array.final_sensor_data\[20\] net31 vssd1 vssd1 vccd1
+ vccd1 _0203_ sky130_fd_sc_hd__mux2_1
X_1368_ _0979_ _0981_ vssd1 vssd1 vccd1 vccd1 _0982_ sky130_fd_sc_hd__nor2_1
X_1299_ dut.ball_pos_y\[2\] vssd1 vssd1 vccd1 vccd1 _0923_ sky130_fd_sc_hd__inv_2
XFILLER_23_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2271_ net28 _0659_ _0661_ vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__and3_1
X_2340_ _0332_ _0720_ _0725_ _0726_ vssd1 vssd1 vccd1 vccd1 _0727_ sky130_fd_sc_hd__o22a_1
XFILLER_52_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1986_ net314 _0442_ _0445_ vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_9_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2607_ _0858_ _0902_ _0860_ vssd1 vssd1 vccd1 vccd1 _0903_ sky130_fd_sc_hd__o21ba_1
X_2469_ _0815_ _0820_ vssd1 vssd1 vccd1 vccd1 _0821_ sky130_fd_sc_hd__or2_1
X_2538_ dut.ir_sensor_array.final_sensor_data\[4\] dut.ir_sensor_array.final_sensor_data\[3\]
+ net32 vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_41_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1840_ _0350_ _0351_ net26 net25 vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_x.pwm_out
+ sky130_fd_sc_hd__o211a_1
X_1771_ net46 _1254_ _0288_ vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__o21a_1
XFILLER_6_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2254_ _0583_ _0624_ _0603_ vssd1 vssd1 vccd1 vccd1 _0650_ sky130_fd_sc_hd__o21ai_1
XFILLER_40_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2323_ _0700_ _0710_ vssd1 vssd1 vccd1 vccd1 _0711_ sky130_fd_sc_hd__or2_1
X_2185_ _0585_ _0587_ vssd1 vssd1 vccd1 vccd1 _0588_ sky130_fd_sc_hd__nor2_1
XFILLER_40_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1969_ dut.microstep_x.ctr\[7\] dut.microstep_x.ctr\[6\] _0958_ vssd1 vssd1 vccd1
+ vccd1 _0433_ sky130_fd_sc_hd__nand3_1
XFILLER_0_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4 dut.microstep_x.ctr\[0\] vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_62_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1823_ _0282_ _0322_ _0323_ _0326_ _0328_ vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__a32o_1
X_2872_ clknet_leaf_0_clk _0002_ net50 vssd1 vssd1 vccd1 vccd1 dut.clkdiv_inst.counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1685_ dut.actual_duty_x\[5\] _1244_ _1245_ vssd1 vssd1 vccd1 vccd1 _1255_ sky130_fd_sc_hd__nor3_1
X_1754_ _0265_ _0271_ vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__or2_1
XFILLER_57_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2237_ net81 _0638_ vssd1 vssd1 vccd1 vccd1 _0118_ sky130_fd_sc_hd__and2_1
XFILLER_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2306_ _0227_ _0678_ vssd1 vssd1 vccd1 vccd1 _0694_ sky130_fd_sc_hd__nor2_1
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2099_ _0515_ _0518_ vssd1 vssd1 vccd1 vccd1 _0519_ sky130_fd_sc_hd__and2_1
X_2168_ _0570_ vssd1 vssd1 vccd1 vccd1 _0571_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1470_ _1053_ _1058_ _1050_ _1052_ vssd1 vssd1 vccd1 vccd1 _1059_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_22_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2022_ _0466_ _0467_ vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__nor2_1
X_2786_ clknet_leaf_7_clk _0140_ net65 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_200ms\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_2855_ clknet_leaf_3_clk _0208_ net59 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_1806_ _0282_ _0322_ _0323_ vssd1 vssd1 vccd1 vccd1 _0324_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1668_ net236 _1238_ _1240_ vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_y.count_d\[15\]
+ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_37_Left_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1599_ _1134_ _1182_ vssd1 vssd1 vccd1 vccd1 _1188_ sky130_fd_sc_hd__nand2_1
X_1737_ net49 dut.actual_duty_x\[2\] vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_28_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_46_Left_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_10_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_55_Left_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_25_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2640_ clknet_leaf_14_clk _0111_ net83 vssd1 vssd1 vccd1 vccd1 dut.spi.state_q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1453_ dut.pwm_a_inst_y.count_q\[13\] _1041_ vssd1 vssd1 vccd1 vccd1 _1042_ sky130_fd_sc_hd__xnor2_1
X_1522_ net39 _1109_ _1108_ vssd1 vssd1 vccd1 vccd1 _1111_ sky130_fd_sc_hd__a21oi_1
X_2571_ net319 dut.ir_sensor_array.final_sensor_data\[36\] net34 vssd1 vssd1 vccd1
+ vccd1 _0219_ sky130_fd_sc_hd__mux2_1
X_1384_ dut.spi.cs_low_counter_q\[1\] net231 _0992_ vssd1 vssd1 vccd1 vccd1 dut.spi.cs_low_counter_d\[1\]
+ sky130_fd_sc_hd__a21oi_1
X_2005_ _0456_ _0457_ vssd1 vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__nor2_1
XFILLER_23_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2769_ clknet_leaf_28_clk _0040_ net51 vssd1 vssd1 vccd1 vccd1 dut.microstep_x.ctr\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_2838_ clknet_leaf_26_clk _0191_ net59 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout58_A net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2623_ clknet_leaf_15_clk dut.spi.clk_counter_d\[3\] net84 vssd1 vssd1 vccd1 vccd1
+ dut.spi.clk_counter_q\[3\] sky130_fd_sc_hd__dfrtp_1
X_2554_ dut.ir_sensor_array.final_sensor_data\[20\] dut.ir_sensor_array.final_sensor_data\[19\]
+ net33 vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__mux2_1
X_1367_ dut.spi.clk_counter_q\[3\] dut.spi.clk_counter_q\[2\] dut.spi.clk_counter_q\[5\]
+ dut.spi.clk_counter_q\[4\] vssd1 vssd1 vccd1 vccd1 _0981_ sky130_fd_sc_hd__or4b_1
X_1436_ net200 _1026_ _1029_ vssd1 vssd1 vccd1 vccd1 _0021_ sky130_fd_sc_hd__o21a_1
X_1505_ net39 dut.actual_duty_y\[3\] vssd1 vssd1 vccd1 vccd1 _1094_ sky130_fd_sc_hd__or2_1
X_2485_ _1189_ _0813_ vssd1 vssd1 vccd1 vccd1 _0836_ sky130_fd_sc_hd__or2_1
XFILLER_28_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1298_ dut.actual_duty_x\[0\] vssd1 vssd1 vccd1 vccd1 _0922_ sky130_fd_sc_hd__inv_2
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2270_ _0660_ vssd1 vssd1 vccd1 vccd1 _0661_ sky130_fd_sc_hd__inv_2
X_1985_ net16 _0444_ vssd1 vssd1 vccd1 vccd1 _0445_ sky130_fd_sc_hd__nor2_1
X_2606_ _0853_ _0901_ _0855_ vssd1 vssd1 vccd1 vccd1 _0902_ sky130_fd_sc_hd__o21ba_1
X_2537_ dut.ir_sensor_array.final_sensor_data\[3\] dut.ir_sensor_array.final_sensor_data\[2\]
+ net32 vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__mux2_1
X_1419_ _0934_ net14 _1017_ vssd1 vssd1 vccd1 vccd1 _0030_ sky130_fd_sc_hd__nor3_1
X_2399_ _0760_ net209 vssd1 vssd1 vccd1 vccd1 _0157_ sky130_fd_sc_hd__nor2_1
X_2468_ net39 _0814_ vssd1 vssd1 vccd1 vccd1 _0820_ sky130_fd_sc_hd__nor2_1
XFILLER_43_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_6_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1770_ net47 _1245_ vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__nand2_1
XFILLER_6_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2253_ net159 net19 net79 _0649_ vssd1 vssd1 vccd1 vccd1 _0123_ sky130_fd_sc_hd__o211a_1
X_2184_ _0553_ _0586_ vssd1 vssd1 vccd1 vccd1 _0587_ sky130_fd_sc_hd__nand2b_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2322_ dut.actual_duty_x\[2\] _0267_ dut.actual_duty_x\[3\] vssd1 vssd1 vccd1 vccd1
+ _0710_ sky130_fd_sc_hd__a21oi_1
X_1899_ dut.microstep_y.ctr\[9\] dut.microstep_y.ctr\[10\] _0390_ _0391_ vssd1 vssd1
+ vccd1 vccd1 _0392_ sky130_fd_sc_hd__or4b_1
XFILLER_33_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1968_ dut.microstep_x.ctr\[6\] _0958_ dut.microstep_x.ctr\[7\] vssd1 vssd1 vccd1
+ vccd1 _0432_ sky130_fd_sc_hd__a21o_1
XFILLER_0_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5 dut.microstep_y.ctr\[0\] vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_62_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_364 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2871_ clknet_leaf_3_clk _0224_ net61 vssd1 vssd1 vccd1 vccd1 dut.ball_pos_x\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_29_Left_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1753_ _0266_ _0270_ vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__or2_1
X_1822_ _0326_ _0328_ _0330_ _0338_ _0339_ vssd1 vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__o221a_1
XANTENNA__2502__S dut.clk_en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1684_ _1244_ _1245_ net47 vssd1 vssd1 vccd1 vccd1 _1254_ sky130_fd_sc_hd__o21a_1
X_2236_ dut.data_in\[1\] _0938_ _0631_ _0637_ vssd1 vssd1 vccd1 vccd1 _0638_ sky130_fd_sc_hd__a22o_1
X_2167_ _0560_ _0566_ _0569_ _0907_ vssd1 vssd1 vccd1 vccd1 _0570_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_0_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2305_ _0677_ _0681_ _0683_ _0684_ _0692_ vssd1 vssd1 vccd1 vccd1 _0693_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_13_Left_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2098_ _0977_ _0516_ vssd1 vssd1 vccd1 vccd1 _0518_ sky130_fd_sc_hd__or2_1
XFILLER_53_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2021_ dut.microstep_x.ctr\[25\] _0465_ vssd1 vssd1 vccd1 vccd1 _0467_ sky130_fd_sc_hd__and2_1
XFILLER_62_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2854_ clknet_leaf_3_clk _0207_ net61 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_1736_ net49 dut.actual_duty_x\[2\] vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__and2_1
X_2785_ clknet_leaf_0_clk _0057_ net51 vssd1 vssd1 vccd1 vccd1 dut.microstep_x.ctr\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_1805_ dut.pwm_a_inst_x.count_q\[6\] _0293_ vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__xnor2_1
X_1667_ dut.pwm_a_inst_y.count_q\[15\] _1238_ net22 vssd1 vssd1 vccd1 vccd1 _1240_
+ sky130_fd_sc_hd__o21ai_1
X_1598_ dut.pwm_a_inst_y.count_q\[2\] _1185_ vssd1 vssd1 vccd1 vccd1 _1187_ sky130_fd_sc_hd__nand2_1
XFILLER_53_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2219_ _0621_ vssd1 vssd1 vccd1 vccd1 _0622_ sky130_fd_sc_hd__inv_2
XFILLER_26_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2570_ dut.ir_sensor_array.final_sensor_data\[36\] net274 net34 vssd1 vssd1 vccd1
+ vccd1 _0218_ sky130_fd_sc_hd__mux2_1
X_1383_ dut.spi.cs_low_counter_q\[1\] dut.spi.cs_low_counter_q\[0\] _0991_ vssd1 vssd1
+ vccd1 vccd1 _0992_ sky130_fd_sc_hd__o21ai_1
X_1452_ dut.pwm_a_inst_y.count_q\[12\] _1040_ vssd1 vssd1 vccd1 vccd1 _1041_ sky130_fd_sc_hd__or2_1
X_1521_ _1108_ _1109_ vssd1 vssd1 vccd1 vccd1 _1110_ sky130_fd_sc_hd__nand2b_1
X_2004_ dut.microstep_x.ctr\[17\] dut.microstep_x.ctr\[18\] _0453_ vssd1 vssd1 vccd1
+ vccd1 _0457_ sky130_fd_sc_hd__and3_1
XFILLER_50_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2768_ clknet_leaf_28_clk _0039_ net51 vssd1 vssd1 vccd1 vccd1 dut.microstep_x.ctr\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_1719_ _0235_ _0236_ vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__nand2_1
X_2837_ clknet_leaf_25_clk _0190_ net60 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_2699_ clknet_leaf_24_clk dut.pwm_a_inst_x.count_d\[2\] net74 vssd1 vssd1 vccd1 vccd1
+ dut.pwm_a_inst_x.count_q\[2\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_16_Left_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2622_ clknet_leaf_16_clk dut.spi.clk_counter_d\[2\] net84 vssd1 vssd1 vccd1 vccd1
+ dut.spi.clk_counter_q\[2\] sky130_fd_sc_hd__dfrtp_1
X_1504_ _1081_ _1092_ vssd1 vssd1 vccd1 vccd1 _1093_ sky130_fd_sc_hd__nand2_1
X_2553_ dut.ir_sensor_array.final_sensor_data\[19\] dut.ir_sensor_array.final_sensor_data\[18\]
+ net33 vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__mux2_1
X_1366_ _0976_ _0979_ _0980_ vssd1 vssd1 vccd1 vccd1 dut.spi.clk_counter_d\[1\] sky130_fd_sc_hd__and3_1
X_1435_ _1019_ _1028_ vssd1 vssd1 vccd1 vccd1 _1029_ sky130_fd_sc_hd__nor2_1
X_2484_ net42 _0835_ net44 vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__mux2_1
X_1297_ dut.actual_duty_x\[1\] vssd1 vssd1 vccd1 vccd1 _0921_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_24_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout70_A net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_1_Left_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1984_ dut.microstep_x.ctr\[11\] _0442_ vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__and2_1
X_2467_ _1048_ _0814_ _0818_ vssd1 vssd1 vccd1 vccd1 _0819_ sky130_fd_sc_hd__a21o_1
X_2605_ _0870_ _0869_ vssd1 vssd1 vccd1 vccd1 _0901_ sky130_fd_sc_hd__and2b_1
X_2536_ dut.ir_sensor_array.final_sensor_data\[2\] net307 net32 vssd1 vssd1 vccd1
+ vccd1 _0184_ sky130_fd_sc_hd__mux2_1
X_2398_ dut.lcd1602.cnt_200ms\[16\] _0758_ net208 vssd1 vssd1 vccd1 vccd1 _0761_ sky130_fd_sc_hd__a21oi_1
X_1418_ dut.lcd1602.cnt_500hz\[4\] _0933_ net288 vssd1 vssd1 vccd1 vccd1 _1017_ sky130_fd_sc_hd__a21oi_1
X_1349_ dut.clkdiv_inst.counter\[16\] dut.clkdiv_inst.counter\[13\] _0967_ vssd1 vssd1
+ vccd1 vccd1 _0968_ sky130_fd_sc_hd__or3_1
XFILLER_28_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire30 _0865_ vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_1
XFILLER_11_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2321_ dut.actual_duty_x\[2\] _0674_ _0708_ _0267_ vssd1 vssd1 vccd1 vccd1 _0709_
+ sky130_fd_sc_hd__o211a_1
X_2252_ net19 _0608_ vssd1 vssd1 vccd1 vccd1 _0649_ sky130_fd_sc_hd__nand2_1
X_2183_ _0907_ _0558_ _0547_ vssd1 vssd1 vccd1 vccd1 _0586_ sky130_fd_sc_hd__o21ba_1
X_1898_ dut.microstep_y.ctr\[7\] dut.microstep_y.ctr\[6\] dut.microstep_y.ctr\[15\]
+ dut.microstep_y.ctr\[16\] vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__and4b_1
X_1967_ net272 _0958_ vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__xor2_1
X_2519_ dut.ir_sensor_array.final_sensor_data\[16\] dut.ir_sensor_array.final_sensor_data\[17\]
+ vssd1 vssd1 vccd1 vccd1 _0859_ sky130_fd_sc_hd__nor2_1
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6 dut.data_in\[3\] vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_47_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2870_ clknet_leaf_12_clk _0223_ net71 vssd1 vssd1 vccd1 vccd1 dut.ball_pos_x\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_10_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_30_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1683_ _1243_ _1244_ _1252_ vssd1 vssd1 vccd1 vccd1 _1253_ sky130_fd_sc_hd__or3_1
X_1752_ _0921_ _0922_ _0269_ vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__a21o_1
X_1821_ _0277_ _0329_ _0338_ dut.pwm_a_inst_x.count_q\[4\] vssd1 vssd1 vccd1 vccd1
+ _0339_ sky130_fd_sc_hd__a31o_1
X_2304_ _0683_ _0684_ _0690_ _0691_ _0686_ vssd1 vssd1 vccd1 vccd1 _0692_ sky130_fd_sc_hd__o221a_1
X_2097_ _0977_ _0516_ vssd1 vssd1 vccd1 vccd1 _0517_ sky130_fd_sc_hd__nor2_1
X_2235_ _0616_ _0626_ _0636_ vssd1 vssd1 vccd1 vccd1 _0637_ sky130_fd_sc_hd__or3_1
X_2166_ dut.lcd1602.currentState\[4\] _0567_ _0568_ vssd1 vssd1 vccd1 vccd1 _0569_
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Left_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2020_ net285 _0465_ vssd1 vssd1 vccd1 vccd1 _0466_ sky130_fd_sc_hd__nor2_1
XFILLER_62_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2853_ clknet_leaf_2_clk _0206_ net59 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_1666_ _1238_ _1239_ vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_y.count_d\[14\] sky130_fd_sc_hd__nor2_1
X_2784_ clknet_leaf_28_clk _0056_ net51 vssd1 vssd1 vccd1 vccd1 dut.microstep_x.ctr\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_1735_ _0920_ _0243_ vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__xnor2_1
X_1804_ _0263_ _0280_ _0281_ vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__or3_1
X_1597_ _1185_ vssd1 vssd1 vccd1 vccd1 _1186_ sky130_fd_sc_hd__inv_2
X_2149_ dut.lcd1602.currentState\[4\] dut.lcd1602.currentState\[0\] net43 vssd1 vssd1
+ vccd1 vccd1 _0552_ sky130_fd_sc_hd__or3b_1
X_2218_ _0613_ _0616_ _0619_ _0620_ vssd1 vssd1 vccd1 vccd1 _0621_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_11_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2657__RESET_B net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1520_ dut.actual_duty_y\[3\] net41 vssd1 vssd1 vccd1 vccd1 _1109_ sky130_fd_sc_hd__or2_1
X_1382_ dut.spi.cs_low_counter_q\[0\] _0991_ vssd1 vssd1 vccd1 vccd1 dut.spi.cs_low_counter_d\[0\]
+ sky130_fd_sc_hd__and2b_1
X_1451_ dut.pwm_a_inst_y.count_q\[10\] dut.pwm_a_inst_y.count_q\[9\] _1038_ dut.pwm_a_inst_y.count_q\[11\]
+ vssd1 vssd1 vccd1 vccd1 _1040_ sky130_fd_sc_hd__a31o_1
XFILLER_4_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2003_ dut.microstep_x.ctr\[17\] _0453_ net263 vssd1 vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__a21oi_1
XFILLER_31_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2836_ clknet_leaf_26_clk _0189_ net60 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_1649_ dut.pwm_a_inst_y.count_q\[8\] dut.pwm_a_inst_y.count_q\[7\] _1225_ vssd1 vssd1
+ vccd1 vccd1 _1229_ sky130_fd_sc_hd__and3_1
X_2698_ clknet_leaf_19_clk net241 net74 vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_x.count_q\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2767_ clknet_leaf_28_clk _0038_ net57 vssd1 vssd1 vccd1 vccd1 dut.microstep_x.ctr\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_1718_ _0233_ _0234_ vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__nand2_1
XFILLER_58_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2621_ clknet_leaf_16_clk dut.spi.clk_counter_d\[1\] net84 vssd1 vssd1 vccd1 vccd1
+ dut.spi.clk_counter_q\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_56_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1503_ _0916_ _1080_ vssd1 vssd1 vccd1 vccd1 _1092_ sky130_fd_sc_hd__nand2_1
X_2483_ _0783_ _0917_ _0834_ vssd1 vssd1 vccd1 vccd1 _0835_ sky130_fd_sc_hd__mux2_1
X_2552_ dut.ir_sensor_array.final_sensor_data\[18\] dut.ir_sensor_array.final_sensor_data\[17\]
+ net33 vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__mux2_1
X_1365_ dut.spi.clk_counter_q\[1\] dut.spi.clk_counter_q\[0\] vssd1 vssd1 vccd1 vccd1
+ _0980_ sky130_fd_sc_hd__or2_1
X_1434_ dut.lcd1602.cnt_500hz\[9\] dut.lcd1602.cnt_500hz\[10\] _1025_ vssd1 vssd1
+ vccd1 vccd1 _1028_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_38_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1296_ dut.actual_duty_x\[2\] vssd1 vssd1 vccd1 vccd1 _0920_ sky130_fd_sc_hd__inv_2
X_2819_ clknet_leaf_20_clk _0172_ net77 vssd1 vssd1 vccd1 vccd1 dut.actual_duty_y\[4\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2604_ _0926_ _0862_ _0900_ _0944_ dut.ball_pos_x\[1\] vssd1 vssd1 vccd1 vccd1 _0223_
+ sky130_fd_sc_hd__a32o_1
X_1983_ _0442_ _0443_ vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__nor2_1
X_1417_ net14 _1016_ vssd1 vssd1 vccd1 vccd1 _0029_ sky130_fd_sc_hd__nor2_1
X_2466_ net38 _0815_ vssd1 vssd1 vccd1 vccd1 _0818_ sky130_fd_sc_hd__nor2_1
X_2535_ net307 _0929_ net32 vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__mux2_1
X_2397_ dut.lcd1602.cnt_200ms\[17\] dut.lcd1602.cnt_200ms\[16\] _0758_ vssd1 vssd1
+ vccd1 vccd1 _0760_ sky130_fd_sc_hd__and3_1
X_1279_ dut.lcd1602.currentState\[5\] vssd1 vssd1 vccd1 vccd1 _0907_ sky130_fd_sc_hd__inv_2
X_1348_ dut.clkdiv_inst.counter\[15\] dut.clkdiv_inst.counter\[14\] dut.clkdiv_inst.counter\[9\]
+ dut.clkdiv_inst.counter\[8\] vssd1 vssd1 vccd1 vccd1 _0967_ sky130_fd_sc_hd__or4bb_1
XFILLER_28_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_57_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2251_ net187 net19 _0621_ _0630_ net79 vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__o221a_1
XFILLER_6_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2320_ _0688_ _0707_ _0676_ vssd1 vssd1 vccd1 vccd1 _0708_ sky130_fd_sc_hd__a21o_1
X_2182_ _0576_ _0580_ vssd1 vssd1 vccd1 vccd1 _0585_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_23_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1966_ _0958_ net164 vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__nor2_1
XFILLER_18_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1897_ dut.microstep_y.ctr\[8\] dut.microstep_y.ctr\[11\] vssd1 vssd1 vccd1 vccd1
+ _0390_ sky130_fd_sc_hd__nand2_1
X_2449_ _0775_ _0777_ _0788_ vssd1 vssd1 vccd1 vccd1 _0801_ sky130_fd_sc_hd__o21a_1
XFILLER_0_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2518_ dut.ir_sensor_array.final_sensor_data\[23\] dut.ir_sensor_array.final_sensor_data\[22\]
+ dut.ir_sensor_array.final_sensor_data\[21\] dut.ir_sensor_array.final_sensor_data\[20\]
+ vssd1 vssd1 vccd1 vccd1 _0858_ sky130_fd_sc_hd__or4_1
XFILLER_56_388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7 dut.data_in\[6\] vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_47_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1820_ dut.pwm_a_inst_x.count_q\[3\] _0335_ _0337_ _0276_ vssd1 vssd1 vccd1 vccd1
+ _0338_ sky130_fd_sc_hd__o22ai_1
XTAP_TAPCELL_ROW_17_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1682_ net49 _1248_ _1250_ vssd1 vssd1 vccd1 vccd1 _1252_ sky130_fd_sc_hd__a21oi_1
X_1751_ _0920_ _0268_ vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__and2_1
X_2234_ dut.ball_pos_y\[1\] _0923_ _0632_ _0610_ dut.ball_pos_x\[1\] vssd1 vssd1 vccd1
+ vccd1 _0636_ sky130_fd_sc_hd__a32o_1
X_2303_ net11 _0685_ _0688_ _0332_ vssd1 vssd1 vccd1 vccd1 _0691_ sky130_fd_sc_hd__a2bb2o_1
X_2096_ dut.spi.spi_clk_q _0982_ vssd1 vssd1 vccd1 vccd1 _0516_ sky130_fd_sc_hd__nand2_1
XFILLER_53_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2165_ dut.lcd1602.currentState\[1\] _0563_ vssd1 vssd1 vccd1 vccd1 _0568_ sky130_fd_sc_hd__xnor2_1
XFILLER_38_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1949_ _0422_ _0423_ vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__nor2_1
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2783_ clknet_leaf_0_clk _0055_ net52 vssd1 vssd1 vccd1 vccd1 dut.microstep_x.ctr\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_1803_ dut.pwm_a_inst_x.count_q\[7\] _0294_ vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__xor2_1
X_2852_ clknet_leaf_2_clk _0205_ net54 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_1665_ dut.pwm_a_inst_y.count_q\[14\] _1237_ net22 vssd1 vssd1 vccd1 vccd1 _1239_
+ sky130_fd_sc_hd__o21ai_1
X_1596_ _1183_ _1184_ vssd1 vssd1 vccd1 vccd1 _1185_ sky130_fd_sc_hd__nand2_1
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1734_ _0239_ _0247_ vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__xnor2_1
X_2217_ _0592_ _0599_ _0601_ _0554_ _0617_ vssd1 vssd1 vccd1 vccd1 _0620_ sky130_fd_sc_hd__o221a_1
XFILLER_38_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2148_ dut.lcd1602.currentState\[3\] _0550_ vssd1 vssd1 vccd1 vccd1 _0551_ sky130_fd_sc_hd__nand2_1
X_2079_ dut.ball_pos_y\[0\] dut.ball_pos_y\[2\] _0501_ vssd1 vssd1 vccd1 vccd1 _0502_
+ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1450_ dut.pwm_a_inst_y.count_q\[9\] _1038_ vssd1 vssd1 vccd1 vccd1 _1039_ sky130_fd_sc_hd__nand2_1
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1381_ dut.spi.cs_low_counter_q\[5\] _0990_ _0975_ vssd1 vssd1 vccd1 vccd1 _0991_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_4_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2002_ dut.microstep_x.ctr\[17\] _0453_ _0455_ vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__o21ba_1
XANTENNA_clkbuf_0_clk_X clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2766_ clknet_leaf_27_clk _0037_ net57 vssd1 vssd1 vccd1 vccd1 dut.microstep_x.ctr\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_2835_ clknet_leaf_26_clk _0188_ net58 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_1648_ dut.pwm_a_inst_y.count_q\[7\] dut.pwm_a_inst_y.count_q\[6\] _1224_ dut.pwm_a_inst_y.count_q\[8\]
+ vssd1 vssd1 vccd1 vccd1 _1228_ sky130_fd_sc_hd__a31o_1
X_1579_ _1164_ _1166_ vssd1 vssd1 vccd1 vccd1 _1168_ sky130_fd_sc_hd__nand2_1
X_2697_ clknet_leaf_19_clk dut.pwm_a_inst_x.count_d\[0\] net74 vssd1 vssd1 vccd1 vccd1
+ dut.pwm_a_inst_x.count_q\[0\] sky130_fd_sc_hd__dfrtp_2
X_1717_ _0233_ _0234_ vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__or2_1
XFILLER_41_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2620_ clknet_leaf_15_clk dut.spi.clk_counter_d\[0\] net82 vssd1 vssd1 vccd1 vccd1
+ dut.spi.clk_counter_q\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1433_ net250 _1025_ _1027_ vssd1 vssd1 vccd1 vccd1 _0034_ sky130_fd_sc_hd__o21a_1
X_1502_ _1086_ _1090_ vssd1 vssd1 vccd1 vccd1 _1091_ sky130_fd_sc_hd__nand2_1
X_2482_ _1056_ _0805_ _0813_ _0833_ vssd1 vssd1 vccd1 vccd1 _0834_ sky130_fd_sc_hd__o211ai_4
X_2551_ net310 dut.ir_sensor_array.final_sensor_data\[17\] _0943_ vssd1 vssd1 vccd1
+ vccd1 _0199_ sky130_fd_sc_hd__mux2_1
X_1364_ dut.spi.clk_counter_q\[1\] dut.spi.clk_counter_q\[0\] vssd1 vssd1 vccd1 vccd1
+ _0979_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_38_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1295_ dut.actual_duty_x\[6\] vssd1 vssd1 vccd1 vccd1 _0919_ sky130_fd_sc_hd__inv_2
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2818_ clknet_leaf_19_clk _0171_ net74 vssd1 vssd1 vccd1 vccd1 dut.actual_duty_y\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_2749_ clknet_leaf_27_clk _0134_ net75 vssd1 vssd1 vccd1 vccd1 dut.actual_duty_x\[2\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_54_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout56_A net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1982_ dut.microstep_x.ctr\[9\] _0440_ net270 vssd1 vssd1 vccd1 vccd1 _0443_ sky130_fd_sc_hd__a21oi_1
X_2603_ dut.ir_sensor_array.final_sensor_data\[35\] dut.ir_sensor_array.final_sensor_data\[34\]
+ _0899_ vssd1 vssd1 vccd1 vccd1 _0900_ sky130_fd_sc_hd__or3_1
X_2534_ dut.ball_pos_y\[2\] _0944_ _0867_ _0871_ vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__a22o_1
X_1416_ dut.lcd1602.cnt_500hz\[4\] _0933_ vssd1 vssd1 vccd1 vccd1 _1016_ sky130_fd_sc_hd__xnor2_1
X_2396_ net201 _0758_ vssd1 vssd1 vccd1 vccd1 _0156_ sky130_fd_sc_hd__xor2_1
X_2465_ net36 _0816_ vssd1 vssd1 vccd1 vccd1 _0817_ sky130_fd_sc_hd__or2_1
X_1347_ _0959_ _0960_ _0961_ _0966_ vssd1 vssd1 vccd1 vccd1 _0035_ sky130_fd_sc_hd__nor4_1
X_1278_ dut.lcd1602.currentState\[4\] vssd1 vssd1 vccd1 vccd1 _0906_ sky130_fd_sc_hd__inv_2
XFILLER_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_86 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2250_ net160 net18 net79 _0648_ vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__o211a_1
X_2181_ _0583_ vssd1 vssd1 vccd1 vccd1 _0584_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_63_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1965_ dut.microstep_x.ctr\[4\] _0957_ net163 vssd1 vssd1 vccd1 vccd1 _0431_ sky130_fd_sc_hd__a21oi_1
X_1896_ dut.microstep_y.ctr\[7\] dut.microstep_y.ctr\[6\] _0947_ vssd1 vssd1 vccd1
+ vccd1 _0389_ sky130_fd_sc_hd__nand3_1
X_2517_ dut.ir_sensor_array.final_sensor_data\[21\] dut.ir_sensor_array.final_sensor_data\[20\]
+ vssd1 vssd1 vccd1 vccd1 _0857_ sky130_fd_sc_hd__nor2_1
X_2379_ dut.lcd1602.cnt_200ms\[9\] _0748_ vssd1 vssd1 vccd1 vccd1 _0750_ sky130_fd_sc_hd__nand2_1
X_2448_ _0792_ _0796_ _0799_ _0791_ vssd1 vssd1 vccd1 vccd1 _0800_ sky130_fd_sc_hd__a22o_1
XFILLER_24_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold8 dut.data_in\[4\] vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__dlygate4sd3_1
X_1750_ dut.actual_duty_x\[1\] dut.actual_duty_x\[0\] vssd1 vssd1 vccd1 vccd1 _0268_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_17_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1681_ _1247_ _1250_ vssd1 vssd1 vccd1 vccd1 _1251_ sky130_fd_sc_hd__nor2_1
X_2233_ net81 _0635_ vssd1 vssd1 vccd1 vccd1 _0117_ sky130_fd_sc_hd__and2_1
X_2164_ net43 _0544_ dut.lcd1602.currentState\[4\] vssd1 vssd1 vccd1 vccd1 _0567_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_38_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2302_ _0267_ _0268_ _0689_ _0687_ vssd1 vssd1 vccd1 vccd1 _0690_ sky130_fd_sc_hd__a31oi_1
X_2095_ dut.lcd1602.out_valid _0513_ vssd1 vssd1 vccd1 vccd1 _0515_ sky130_fd_sc_hd__nand2_2
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1948_ dut.microstep_y.ctr\[25\] _0421_ vssd1 vssd1 vccd1 vccd1 _0423_ sky130_fd_sc_hd__and2_1
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_80 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1879_ _0380_ _0381_ vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_x.count_d\[14\] sky130_fd_sc_hd__nor2_1
XFILLER_0_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_3__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_35_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkload1_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1733_ _0248_ _0250_ vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__xnor2_1
X_1802_ _0283_ _0319_ vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__nor2_1
X_2782_ clknet_leaf_0_clk _0054_ net50 vssd1 vssd1 vccd1 vccd1 dut.microstep_x.ctr\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_2851_ clknet_leaf_2_clk _0204_ net54 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_1664_ dut.pwm_a_inst_y.count_q\[14\] _1237_ vssd1 vssd1 vccd1 vccd1 _1238_ sky130_fd_sc_hd__and2_1
X_1595_ net41 _1182_ vssd1 vssd1 vccd1 vccd1 _1184_ sky130_fd_sc_hd__or2_1
X_2147_ net43 _0548_ vssd1 vssd1 vccd1 vccd1 _0550_ sky130_fd_sc_hd__nand2_1
X_2216_ _0585_ _0618_ vssd1 vssd1 vccd1 vccd1 _0619_ sky130_fd_sc_hd__nor2_1
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2078_ dut.ball_pos_y\[1\] _0498_ _0500_ vssd1 vssd1 vccd1 vccd1 _0501_ sky130_fd_sc_hd__or3b_1
XANTENNA_fanout86_A net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1380_ dut.spi.cs_low_counter_q\[3\] dut.spi.cs_low_counter_q\[4\] dut.spi.cs_low_counter_q\[5\]
+ vssd1 vssd1 vccd1 vccd1 _0990_ sky130_fd_sc_hd__or3b_1
X_2001_ dut.microstep_x.ctr\[17\] dut.microstep_x.ctr\[16\] _0451_ _0035_ vssd1 vssd1
+ vccd1 vccd1 _0455_ sky130_fd_sc_hd__a31o_1
XFILLER_50_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2696_ clknet_leaf_15_clk net124 net84 vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_y.count_q\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1716_ _1259_ _1268_ vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__xnor2_1
X_2765_ clknet_leaf_27_clk _0065_ net57 vssd1 vssd1 vccd1 vccd1 dut.microstep_x.ctr\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_2834_ clknet_leaf_26_clk _0187_ net58 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_1647_ net237 _1225_ _1227_ vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_y.count_d\[7\]
+ sky130_fd_sc_hd__a21oi_1
X_1578_ _1164_ _1166_ vssd1 vssd1 vccd1 vccd1 _1167_ sky130_fd_sc_hd__nor2_1
XFILLER_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2550_ dut.ir_sensor_array.final_sensor_data\[16\] dut.ir_sensor_array.final_sensor_data\[15\]
+ net31 vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__mux2_1
X_1363_ dut.spi.clk_counter_q\[1\] dut.spi.clk_counter_q\[0\] vssd1 vssd1 vccd1 vccd1
+ _0978_ sky130_fd_sc_hd__and2_1
X_1432_ net14 _1026_ vssd1 vssd1 vccd1 vccd1 _1027_ sky130_fd_sc_hd__nor2_1
X_1501_ _1083_ _1085_ vssd1 vssd1 vccd1 vccd1 _1090_ sky130_fd_sc_hd__or2_1
X_2481_ _0831_ _0832_ _0817_ vssd1 vssd1 vccd1 vccd1 _0833_ sky130_fd_sc_hd__a21boi_4
XFILLER_48_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Left_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1294_ net313 vssd1 vssd1 vccd1 vccd1 _0918_ sky130_fd_sc_hd__inv_2
XFILLER_63_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_52_Left_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2679_ clknet_leaf_13_clk dut.pwm_a_inst_y.count_d\[2\] net80 vssd1 vssd1 vccd1 vccd1
+ dut.pwm_a_inst_y.count_q\[2\] sky130_fd_sc_hd__dfrtp_1
X_2817_ clknet_leaf_18_clk _0170_ net77 vssd1 vssd1 vccd1 vccd1 dut.actual_duty_y\[2\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_11_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2748_ clknet_leaf_26_clk _0133_ net75 vssd1 vssd1 vccd1 vccd1 dut.actual_duty_x\[1\]
+ sky130_fd_sc_hd__dfstp_2
XPHY_EDGE_ROW_61_Left_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1981_ dut.microstep_x.ctr\[9\] dut.microstep_x.ctr\[10\] _0440_ vssd1 vssd1 vccd1
+ vccd1 _0442_ sky130_fd_sc_hd__and3_1
X_2602_ dut.ir_sensor_array.final_sensor_data\[39\] dut.ir_sensor_array.final_sensor_data\[38\]
+ _0898_ _0864_ vssd1 vssd1 vccd1 vccd1 _0899_ sky130_fd_sc_hd__o31a_1
X_2533_ _0869_ _0870_ _0866_ vssd1 vssd1 vccd1 vccd1 _0871_ sky130_fd_sc_hd__o21ba_1
XANTENNA__2090__S dut.clk_en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1415_ _0933_ net14 _1015_ vssd1 vssd1 vccd1 vccd1 _0028_ sky130_fd_sc_hd__nor3_1
X_2395_ _0758_ _0759_ vssd1 vssd1 vccd1 vccd1 _0155_ sky130_fd_sc_hd__nor2_1
X_2464_ net40 _1044_ _0814_ vssd1 vssd1 vccd1 vccd1 _0816_ sky130_fd_sc_hd__and3_1
X_1346_ _0962_ _0963_ _0964_ _0965_ vssd1 vssd1 vccd1 vccd1 _0966_ sky130_fd_sc_hd__or4_1
XFILLER_51_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_1__f_clk_X clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2180_ net12 _0571_ vssd1 vssd1 vccd1 vccd1 _0583_ sky130_fd_sc_hd__or2_1
XFILLER_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_13_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1895_ dut.microstep_y.ctr\[6\] _0947_ dut.microstep_y.ctr\[7\] vssd1 vssd1 vccd1
+ vccd1 _0388_ sky130_fd_sc_hd__a21o_1
XFILLER_33_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1964_ net167 _0957_ vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__xor2_1
X_2447_ _1134_ _0788_ _0798_ _0790_ _0786_ vssd1 vssd1 vccd1 vccd1 _0799_ sky130_fd_sc_hd__a32o_1
X_2516_ _0853_ _0855_ vssd1 vssd1 vccd1 vccd1 _0856_ sky130_fd_sc_hd__nor2_1
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2378_ _1011_ _0747_ _0749_ vssd1 vssd1 vccd1 vccd1 _0148_ sky130_fd_sc_hd__and3_1
X_1329_ dut.microstep_y.ctr\[7\] dut.microstep_y.ctr\[9\] _0910_ dut.microstep_y.ctr\[6\]
+ vssd1 vssd1 vccd1 vccd1 _0950_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_3_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold9 dut.spi.shift_reg_q\[0\] vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout71_X net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1680_ net47 _1246_ _1248_ vssd1 vssd1 vccd1 vccd1 _1250_ sky130_fd_sc_hd__and3_1
X_2301_ _0512_ _0668_ _0670_ net11 _0675_ vssd1 vssd1 vccd1 vccd1 _0689_ sky130_fd_sc_hd__o32a_1
XFILLER_53_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2232_ dut.data_in\[0\] _0938_ _0631_ _0634_ vssd1 vssd1 vccd1 vccd1 _0635_ sky130_fd_sc_hd__a22o_1
X_2163_ _0555_ dut.lcd1602.currentState\[2\] dut.lcd1602.currentState\[1\] vssd1 vssd1
+ vccd1 vccd1 _0566_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_2_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_24_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2094_ dut.spi.state_q\[2\] dut.spi.state_q\[1\] dut.spi.state_q\[0\] vssd1 vssd1
+ vccd1 vccd1 _0514_ sky130_fd_sc_hd__or3_2
XFILLER_53_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1947_ net279 _0421_ vssd1 vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__nor2_1
XFILLER_9_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1878_ dut.pwm_a_inst_x.count_q\[14\] _0379_ net26 vssd1 vssd1 vccd1 vccd1 _0381_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_37_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Left_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2850_ clknet_leaf_2_clk _0203_ net54 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_1663_ _1237_ net22 _1236_ vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_y.count_d\[13\]
+ sky130_fd_sc_hd__and3b_1
X_1732_ _0233_ _0249_ vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__nand2_1
X_2781_ clknet_leaf_29_clk _0053_ net52 vssd1 vssd1 vccd1 vccd1 dut.microstep_x.ctr\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_1801_ _0251_ _0261_ _0282_ vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_13_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1594_ net41 _1182_ vssd1 vssd1 vccd1 vccd1 _1183_ sky130_fd_sc_hd__nand2_1
XFILLER_7_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2215_ _0586_ _0601_ _0614_ _0595_ vssd1 vssd1 vccd1 vccd1 _0618_ sky130_fd_sc_hd__o211a_1
X_2146_ dut.lcd1602.currentState\[1\] dut.lcd1602.currentState\[0\] vssd1 vssd1 vccd1
+ vccd1 _0549_ sky130_fd_sc_hd__or2_1
XFILLER_38_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2077_ dut.ball_pos_x\[1\] dut.ball_pos_x\[0\] dut.ball_pos_x\[2\] vssd1 vssd1 vccd1
+ vccd1 _0500_ sky130_fd_sc_hd__a21o_1
XFILLER_34_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout79_A net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_34_Left_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2000_ dut.microstep_x.ctr\[16\] _0451_ _0454_ _0439_ vssd1 vssd1 vccd1 vccd1 _0043_
+ sky130_fd_sc_hd__o211a_1
XFILLER_50_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2833_ clknet_leaf_27_clk _0186_ net58 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_2695_ clknet_leaf_15_clk net125 net84 vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_y.count_q\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_1646_ dut.pwm_a_inst_y.count_q\[7\] _1225_ net21 vssd1 vssd1 vccd1 vccd1 _1227_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_6_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1715_ _1275_ _0232_ vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__or2_1
X_2764_ clknet_leaf_28_clk _0064_ net57 vssd1 vssd1 vccd1 vccd1 dut.microstep_x.ctr\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_1577_ dut.pwm_a_inst_y.count_q\[4\] _1165_ _1038_ vssd1 vssd1 vccd1 vccd1 _1166_
+ sky130_fd_sc_hd__o21ba_1
XANTENNA_clkbuf_leaf_21_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2129_ dut.spi.bit_counter_q\[0\] _0517_ dut.spi.bit_counter_q\[1\] vssd1 vssd1 vccd1
+ vccd1 _0535_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_49_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1500_ _1087_ _1088_ vssd1 vssd1 vccd1 vccd1 _1089_ sky130_fd_sc_hd__or2_1
XFILLER_31_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2480_ _0786_ _0819_ _0830_ _0816_ _1046_ vssd1 vssd1 vccd1 vccd1 _0832_ sky130_fd_sc_hd__o221a_1
XFILLER_9_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1362_ net184 _0977_ vssd1 vssd1 vccd1 vccd1 dut.spi.clk_counter_d\[0\] sky130_fd_sc_hd__nor2_1
X_1431_ dut.lcd1602.cnt_500hz\[9\] _1025_ vssd1 vssd1 vccd1 vccd1 _1026_ sky130_fd_sc_hd__and2_1
X_1293_ net42 vssd1 vssd1 vccd1 vccd1 _0917_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_46_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2816_ clknet_leaf_18_clk _0169_ net80 vssd1 vssd1 vccd1 vccd1 dut.actual_duty_y\[1\]
+ sky130_fd_sc_hd__dfstp_2
X_1629_ dut.pwm_a_inst_y.count_q\[1\] dut.pwm_a_inst_y.count_q\[0\] net21 vssd1 vssd1
+ vccd1 vccd1 _1216_ sky130_fd_sc_hd__o21ai_1
X_2678_ clknet_leaf_12_clk dut.pwm_a_inst_y.count_d\[1\] net79 vssd1 vssd1 vccd1 vccd1
+ dut.pwm_a_inst_y.count_q\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2747_ clknet_leaf_26_clk _0132_ net75 vssd1 vssd1 vccd1 vccd1 dut.actual_duty_x\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input3_A nrst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1980_ net256 _0440_ vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__xor2_1
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2463_ _1095_ _1183_ vssd1 vssd1 vccd1 vccd1 _0815_ sky130_fd_sc_hd__nor2_1
X_2601_ dut.ir_sensor_array.final_sensor_data\[27\] dut.ir_sensor_array.final_sensor_data\[26\]
+ _0897_ _0849_ vssd1 vssd1 vccd1 vccd1 _0898_ sky130_fd_sc_hd__o31a_1
X_2532_ dut.ir_sensor_array.final_sensor_data\[3\] dut.ir_sensor_array.final_sensor_data\[2\]
+ dut.ir_sensor_array.final_sensor_data\[1\] _0929_ vssd1 vssd1 vccd1 vccd1 _0870_
+ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_21_Left_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1414_ net302 _0932_ vssd1 vssd1 vccd1 vccd1 _1015_ sky130_fd_sc_hd__nor2_1
X_2394_ net211 _0756_ vssd1 vssd1 vccd1 vccd1 _0759_ sky130_fd_sc_hd__nor2_1
X_1345_ dut.microstep_x.ctr\[23\] dut.microstep_x.ctr\[22\] dut.microstep_x.ctr\[25\]
+ dut.microstep_x.ctr\[24\] vssd1 vssd1 vccd1 vccd1 _0965_ sky130_fd_sc_hd__or4_1
XFILLER_36_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire23 net24 vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
XANTENNA_fanout61_A net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1894_ net273 _0947_ vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__xor2_1
X_1963_ _0957_ _0430_ vssd1 vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__nor2_1
X_2446_ net42 _0783_ _0797_ dut.actual_duty_y\[1\] vssd1 vssd1 vccd1 vccd1 _0798_
+ sky130_fd_sc_hd__a211o_1
X_2515_ dut.ir_sensor_array.final_sensor_data\[8\] dut.ir_sensor_array.final_sensor_data\[11\]
+ dut.ir_sensor_array.final_sensor_data\[10\] dut.ir_sensor_array.final_sensor_data\[9\]
+ vssd1 vssd1 vccd1 vccd1 _0855_ sky130_fd_sc_hd__or4_1
XFILLER_56_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2377_ _0748_ vssd1 vssd1 vccd1 vccd1 _0749_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_54_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1328_ dut.microstep_y.ctr\[10\] dut.microstep_y.ctr\[12\] dut.microstep_y.ctr\[13\]
+ dut.microstep_y.ctr\[11\] vssd1 vssd1 vccd1 vccd1 _0949_ sky130_fd_sc_hd__or4bb_1
XTAP_TAPCELL_ROW_3_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2231_ dut.ball_pos_y\[0\] _0923_ _0632_ _0633_ vssd1 vssd1 vccd1 vccd1 _0634_ sky130_fd_sc_hd__a31o_1
X_2300_ _0512_ _0668_ _0671_ _0676_ vssd1 vssd1 vccd1 vccd1 _0688_ sky130_fd_sc_hd__a211oi_1
X_2093_ dut.spi.state_q\[2\] _0493_ vssd1 vssd1 vccd1 vccd1 _0513_ sky130_fd_sc_hd__and2b_1
X_2162_ _0907_ _0562_ _0564_ _0556_ _0560_ vssd1 vssd1 vccd1 vccd1 _0565_ sky130_fd_sc_hd__a32o_1
XFILLER_17_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1946_ _0420_ _0421_ vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__nor2_1
X_1877_ dut.pwm_a_inst_x.count_q\[14\] _0379_ vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__and2_1
X_2429_ _0779_ _0780_ vssd1 vssd1 vccd1 vccd1 _0781_ sky130_fd_sc_hd__nand2_1
XFILLER_29_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1800_ _0314_ _0316_ vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_13_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1662_ dut.pwm_a_inst_y.count_q\[13\] dut.pwm_a_inst_y.count_q\[12\] _1234_ vssd1
+ vssd1 vccd1 vccd1 _1237_ sky130_fd_sc_hd__and3_1
XFILLER_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1731_ _1275_ _0232_ vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__nand2_1
X_2780_ clknet_leaf_29_clk _0052_ net50 vssd1 vssd1 vccd1 vccd1 dut.microstep_x.ctr\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_2214_ _0586_ _0600_ _0577_ vssd1 vssd1 vccd1 vccd1 _0617_ sky130_fd_sc_hd__o21ai_1
X_1593_ dut.actual_duty_y\[1\] net42 vssd1 vssd1 vccd1 vccd1 _1182_ sky130_fd_sc_hd__or2_1
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2145_ dut.lcd1602.currentState\[1\] dut.lcd1602.currentState\[0\] vssd1 vssd1 vccd1
+ vccd1 _0548_ sky130_fd_sc_hd__nor2_1
XFILLER_38_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2076_ dut.ball_pos_x\[1\] dut.ball_pos_x\[0\] vssd1 vssd1 vccd1 vccd1 _0499_ sky130_fd_sc_hd__nand2_1
XFILLER_26_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1929_ dut.microstep_y.ctr\[17\] _0409_ _0411_ vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__o21ba_1
XFILLER_30_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold90 dut.spi.shift_reg_q\[6\] vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2832_ clknet_leaf_27_clk _0185_ net58 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_2763_ clknet_leaf_28_clk _0063_ net58 vssd1 vssd1 vccd1 vccd1 dut.microstep_x.ctr\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2694_ clknet_leaf_15_clk dut.pwm_a_inst_y.count_d\[17\] net84 vssd1 vssd1 vccd1
+ vccd1 dut.pwm_a_inst_y.count_q\[17\] sky130_fd_sc_hd__dfrtp_1
X_1645_ dut.pwm_a_inst_y.count_q\[6\] _1224_ _1226_ net21 vssd1 vssd1 vccd1 vccd1
+ dut.pwm_a_inst_y.count_d\[6\] sky130_fd_sc_hd__o211a_1
X_1576_ dut.pwm_a_inst_y.count_q\[8\] dut.pwm_a_inst_y.count_q\[5\] _1037_ vssd1 vssd1
+ vccd1 vccd1 _1165_ sky130_fd_sc_hd__or3_1
X_1714_ _1277_ _0229_ _0231_ vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__o21ba_1
X_2128_ _0517_ _0534_ dut.spi.bit_counter_q\[0\] vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2059_ net235 _0485_ _0488_ vssd1 vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__o21a_1
XFILLER_41_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1430_ _1025_ _1018_ _1024_ vssd1 vssd1 vccd1 vccd1 _0033_ sky130_fd_sc_hd__and3b_1
XFILLER_49_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1361_ dut.spi.spi_clk_q _0977_ vssd1 vssd1 vccd1 vccd1 dut.sclk_lcd sky130_fd_sc_hd__or2_1
XFILLER_48_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1292_ dut.actual_duty_y\[1\] vssd1 vssd1 vccd1 vccd1 _0916_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_46_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2746_ clknet_leaf_7_clk _0088_ net65 vssd1 vssd1 vccd1 vccd1 dut.microstep_y.ctr\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_2815_ clknet_leaf_19_clk _0168_ net79 vssd1 vssd1 vccd1 vccd1 dut.actual_duty_y\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1559_ _1145_ _1147_ vssd1 vssd1 vccd1 vccd1 _1148_ sky130_fd_sc_hd__or2_1
X_1628_ _0914_ net21 vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_y.count_d\[0\] sky130_fd_sc_hd__and2_1
X_2677_ clknet_leaf_18_clk dut.pwm_a_inst_y.count_d\[0\] net80 vssd1 vssd1 vccd1 vccd1
+ dut.pwm_a_inst_y.count_q\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_36_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2089__A1 dut.clk_en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2600_ dut.ir_sensor_array.final_sensor_data\[31\] dut.ir_sensor_array.final_sensor_data\[30\]
+ _0896_ _0847_ vssd1 vssd1 vccd1 vccd1 _0897_ sky130_fd_sc_hd__o31a_1
XANTENNA_clkbuf_leaf_20_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1413_ _0932_ net13 _1014_ vssd1 vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__nor3_1
X_2393_ dut.lcd1602.cnt_200ms\[15\] _0756_ vssd1 vssd1 vccd1 vccd1 _0758_ sky130_fd_sc_hd__and2_1
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2462_ _0915_ _1183_ vssd1 vssd1 vccd1 vccd1 _0814_ sky130_fd_sc_hd__nor2_1
XFILLER_5_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2531_ dut.ir_sensor_array.final_sensor_data\[6\] dut.ir_sensor_array.final_sensor_data\[7\]
+ dut.ir_sensor_array.final_sensor_data\[5\] dut.ir_sensor_array.final_sensor_data\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0869_ sky130_fd_sc_hd__or4_1
XFILLER_36_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire24 dut.clkdiv_inst.sck vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
XFILLER_3_84 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1344_ dut.microstep_x.ctr\[27\] dut.microstep_x.ctr\[26\] dut.microstep_x.ctr\[29\]
+ dut.microstep_x.ctr\[28\] vssd1 vssd1 vccd1 vccd1 _0964_ sky130_fd_sc_hd__or4_1
XFILLER_51_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2729_ clknet_leaf_6_clk _0070_ net63 vssd1 vssd1 vccd1 vccd1 dut.microstep_y.ctr\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xteam_02_90 vssd1 vssd1 vccd1 vccd1 team_02_90/HI gpio_oeb[5] sky130_fd_sc_hd__conb_1
XFILLER_6_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2871__RESET_B net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1962_ net190 _0956_ vssd1 vssd1 vccd1 vccd1 _0430_ sky130_fd_sc_hd__nor2_1
X_1893_ _0947_ net175 vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__nor2_1
X_2376_ dut.lcd1602.cnt_200ms\[8\] _1005_ vssd1 vssd1 vccd1 vccd1 _0748_ sky130_fd_sc_hd__and2_1
X_2445_ _0784_ _0788_ vssd1 vssd1 vccd1 vccd1 _0797_ sky130_fd_sc_hd__nand2_1
X_2514_ dut.ir_sensor_array.final_sensor_data\[8\] dut.ir_sensor_array.final_sensor_data\[9\]
+ vssd1 vssd1 vccd1 vccd1 _0854_ sky130_fd_sc_hd__nor2_1
XFILLER_64_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1327_ _0947_ vssd1 vssd1 vccd1 vccd1 _0948_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_49_Left_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_58_Left_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2230_ dut.ball_pos_x\[0\] _0610_ _0623_ _0589_ _0606_ vssd1 vssd1 vccd1 vccd1 _0633_
+ sky130_fd_sc_hd__a2111o_1
X_2161_ dut.lcd1602.currentState\[0\] _0563_ _0544_ _0906_ vssd1 vssd1 vccd1 vccd1
+ _0564_ sky130_fd_sc_hd__a211o_1
XANTENNA_clkbuf_2_2__f_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2092_ dut.pid_x.x_pid.last_error\[2\] _0512_ dut.clk_en vssd1 vssd1 vccd1 vccd1
+ _0099_ sky130_fd_sc_hd__mux2_1
XFILLER_61_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1945_ dut.microstep_y.ctr\[23\] dut.microstep_y.ctr\[24\] _0419_ vssd1 vssd1 vccd1
+ vccd1 _0421_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_16_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1876_ _0379_ net26 _0378_ vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_x.count_d\[13\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_29_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2428_ _0766_ _0777_ _0778_ vssd1 vssd1 vccd1 vccd1 _0780_ sky130_fd_sc_hd__or3_1
XFILLER_28_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2359_ net46 dut.microstep_x.clk_en _0701_ net45 vssd1 vssd1 vccd1 vccd1 _0139_ sky130_fd_sc_hd__a31o_1
XFILLER_56_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1661_ dut.pwm_a_inst_y.count_q\[12\] _1149_ _1229_ dut.pwm_a_inst_y.count_q\[13\]
+ vssd1 vssd1 vccd1 vccd1 _1236_ sky130_fd_sc_hd__a31o_1
X_1592_ _1135_ _1180_ vssd1 vssd1 vccd1 vccd1 _1181_ sky130_fd_sc_hd__and2b_1
X_1730_ _0239_ _0247_ vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__or2_1
XFILLER_11_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2144_ _0543_ _0545_ _0546_ vssd1 vssd1 vccd1 vccd1 _0547_ sky130_fd_sc_hd__o21ai_1
X_2213_ _0576_ _0614_ _0615_ vssd1 vssd1 vccd1 vccd1 _0616_ sky130_fd_sc_hd__o21ai_1
XFILLER_34_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2075_ dut.ball_pos_x\[1\] dut.ball_pos_x\[0\] dut.ball_pos_x\[2\] vssd1 vssd1 vccd1
+ vccd1 _0498_ sky130_fd_sc_hd__o21a_1
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1928_ dut.microstep_y.ctr\[17\] dut.microstep_y.ctr\[16\] _0407_ net17 vssd1 vssd1
+ vccd1 vccd1 _0411_ sky130_fd_sc_hd__a31o_1
X_1859_ dut.pwm_a_inst_x.count_q\[7\] _0367_ net27 vssd1 vssd1 vccd1 vccd1 _0369_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_79 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold80 dut.spi.cs_low_counter_d\[1\] vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 _0106_ vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1713_ _0921_ _0230_ vssd1 vssd1 vccd1 vccd1 _0231_ sky130_fd_sc_hd__nor2_1
X_2831_ clknet_leaf_28_clk _0184_ net57 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2762_ clknet_leaf_28_clk _0062_ net51 vssd1 vssd1 vccd1 vccd1 dut.microstep_x.ctr\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_2693_ clknet_leaf_15_clk dut.pwm_a_inst_y.count_d\[16\] net85 vssd1 vssd1 vccd1
+ vccd1 dut.pwm_a_inst_y.count_q\[16\] sky130_fd_sc_hd__dfrtp_1
X_1644_ _1225_ vssd1 vssd1 vccd1 vccd1 _1226_ sky130_fd_sc_hd__inv_2
X_1575_ _1140_ _1163_ vssd1 vssd1 vccd1 vccd1 _1164_ sky130_fd_sc_hd__or2_1
XFILLER_6_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2127_ _0513_ _0517_ vssd1 vssd1 vccd1 vccd1 _0534_ sky130_fd_sc_hd__nor2_1
XFILLER_54_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2058_ _0019_ _0487_ vssd1 vssd1 vccd1 vccd1 _0488_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_24_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1360_ dut.spi.state_q\[0\] _0975_ vssd1 vssd1 vccd1 vccd1 _0977_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_38_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1291_ dut.actual_duty_y\[3\] vssd1 vssd1 vccd1 vccd1 _0915_ sky130_fd_sc_hd__inv_2
XFILLER_63_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_9_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2676_ clknet_leaf_11_clk _0025_ net70 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_500hz\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_2745_ clknet_leaf_7_clk _0087_ net65 vssd1 vssd1 vccd1 vccd1 dut.microstep_y.ctr\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_2814_ clknet_leaf_3_clk _0167_ net71 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.currentState\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_31_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1627_ dut.pwm_a_inst_y.count_q\[18\] dut.pwm_a_inst_y.count_q\[19\] _1214_ vssd1
+ vssd1 vccd1 vccd1 _1215_ sky130_fd_sc_hd__nor3_1
X_1558_ _1051_ _1059_ _1144_ vssd1 vssd1 vccd1 vccd1 _1147_ sky130_fd_sc_hd__nor3_1
X_1489_ net38 net39 vssd1 vssd1 vccd1 vccd1 _1078_ sky130_fd_sc_hd__or2_1
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout87_X net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_61_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2707__CLK clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2530_ dut.ir_sensor_array.final_sensor_data\[5\] dut.ir_sensor_array.final_sensor_data\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0868_ sky130_fd_sc_hd__nor2_1
X_1412_ dut.lcd1602.cnt_500hz\[1\] dut.lcd1602.cnt_500hz\[0\] net291 vssd1 vssd1 vccd1
+ vccd1 _1014_ sky130_fd_sc_hd__a21oi_1
X_2392_ _0756_ _0757_ vssd1 vssd1 vccd1 vccd1 _0154_ sky130_fd_sc_hd__nor2_1
X_2461_ _0811_ _0812_ vssd1 vssd1 vccd1 vccd1 _0813_ sky130_fd_sc_hd__nor2_2
XFILLER_3_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1343_ dut.microstep_x.ctr\[14\] dut.microstep_x.ctr\[15\] dut.microstep_x.ctr\[17\]
+ dut.microstep_x.ctr\[16\] vssd1 vssd1 vccd1 vccd1 _0963_ sky130_fd_sc_hd__nand4b_1
XFILLER_51_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwire25 _0357_ vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_16_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2728_ clknet_leaf_6_clk _0069_ net63 vssd1 vssd1 vccd1 vccd1 dut.microstep_y.ctr\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_2659_ clknet_leaf_25_clk _0130_ net73 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.bit_count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xteam_02_91 vssd1 vssd1 vccd1 vccd1 team_02_91/HI gpio_oeb[7] sky130_fd_sc_hd__conb_1
XFILLER_2_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1892_ dut.microstep_y.ctr\[4\] _0946_ net174 vssd1 vssd1 vccd1 vccd1 _0387_ sky130_fd_sc_hd__a21oi_1
X_1961_ _0956_ net180 vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__nor2_1
X_2513_ dut.ir_sensor_array.final_sensor_data\[14\] dut.ir_sensor_array.final_sensor_data\[15\]
+ dut.ir_sensor_array.final_sensor_data\[13\] dut.ir_sensor_array.final_sensor_data\[12\]
+ vssd1 vssd1 vccd1 vccd1 _0853_ sky130_fd_sc_hd__or4_1
X_2375_ dut.lcd1602.cnt_200ms\[8\] _1005_ vssd1 vssd1 vccd1 vccd1 _0747_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_5_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1326_ dut.microstep_y.ctr\[5\] dut.microstep_y.ctr\[4\] _0946_ vssd1 vssd1 vccd1
+ vccd1 _0947_ sky130_fd_sc_hd__and3_2
X_2444_ _0794_ _0795_ vssd1 vssd1 vccd1 vccd1 _0796_ sky130_fd_sc_hd__nand2_1
XFILLER_64_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2160_ dut.lcd1602.currentState\[3\] net43 vssd1 vssd1 vccd1 vccd1 _0563_ sky130_fd_sc_hd__xor2_1
XFILLER_38_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2091_ _0506_ _0509_ vssd1 vssd1 vccd1 vccd1 _0512_ sky130_fd_sc_hd__nor2_2
XFILLER_61_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1944_ dut.microstep_y.ctr\[23\] _0419_ net238 vssd1 vssd1 vccd1 vccd1 _0420_ sky130_fd_sc_hd__a21oi_1
X_1875_ dut.pwm_a_inst_x.count_q\[13\] dut.pwm_a_inst_x.count_q\[12\] _0376_ vssd1
+ vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_16_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2427_ _0777_ _0778_ _0766_ vssd1 vssd1 vccd1 vccd1 _0779_ sky130_fd_sc_hd__o21ai_1
X_1309_ dut.lcd1602.cnt_500hz\[3\] _0932_ vssd1 vssd1 vccd1 vccd1 _0933_ sky130_fd_sc_hd__and2_1
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2358_ net46 _0930_ _0738_ _0739_ vssd1 vssd1 vccd1 vccd1 _0138_ sky130_fd_sc_hd__a22o_1
X_2289_ _0509_ net11 vssd1 vssd1 vccd1 vccd1 _0677_ sky130_fd_sc_hd__nor2_1
XFILLER_52_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1660_ net225 _1234_ _1235_ vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_y.count_d\[12\]
+ sky130_fd_sc_hd__a21oi_1
X_1591_ _0915_ net42 _1121_ _1132_ vssd1 vssd1 vccd1 vccd1 _1180_ sky130_fd_sc_hd__a31o_1
X_2143_ dut.lcd1602.currentState\[3\] dut.lcd1602.currentState\[5\] _0544_ net43 vssd1
+ vssd1 vccd1 vccd1 _0546_ sky130_fd_sc_hd__a211o_1
X_2212_ _0570_ _0585_ _0611_ vssd1 vssd1 vccd1 vccd1 _0615_ sky130_fd_sc_hd__or3b_1
XFILLER_38_168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2074_ dut.clkdiv_inst.counter\[11\] _0496_ _0497_ dut.clkdiv_inst.counter\[15\]
+ dut.clkdiv_inst.counter\[14\] vssd1 vssd1 vccd1 vccd1 dut.clkdiv_inst.sck sky130_fd_sc_hd__a2111oi_1
XFILLER_14_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1927_ dut.microstep_y.ctr\[16\] _0407_ _0410_ _0395_ vssd1 vssd1 vccd1 vccd1 _0074_
+ sky130_fd_sc_hd__o211a_1
X_1858_ dut.pwm_a_inst_x.count_q\[6\] _0366_ _0368_ net27 vssd1 vssd1 vccd1 vccd1
+ dut.pwm_a_inst_x.count_d\[6\] sky130_fd_sc_hd__o211a_1
X_1789_ dut.pwm_a_inst_x.count_q\[10\] _0296_ vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__xor2_1
XFILLER_44_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold70 dut.spi.shift_reg_q\[3\] vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 dut.clkdiv_inst.counter\[13\] vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 dut.microstep_x.ctr\[27\] vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_31_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2830_ clknet_leaf_26_clk _0183_ net57 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.final_sensor_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2692_ clknet_leaf_16_clk dut.pwm_a_inst_y.count_d\[15\] net85 vssd1 vssd1 vccd1
+ vccd1 dut.pwm_a_inst_y.count_q\[15\] sky130_fd_sc_hd__dfrtp_1
X_1643_ dut.pwm_a_inst_y.count_q\[6\] _1224_ vssd1 vssd1 vccd1 vccd1 _1225_ sky130_fd_sc_hd__and2_1
XFILLER_6_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1712_ _1277_ _0229_ vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__xnor2_1
X_2761_ clknet_leaf_28_clk _0061_ net51 vssd1 vssd1 vccd1 vccd1 dut.microstep_x.ctr\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_1574_ _1089_ _1103_ _1139_ vssd1 vssd1 vccd1 vccd1 _1163_ sky130_fd_sc_hd__and3_1
X_2126_ dut.spi.state_q\[2\] _0976_ _0532_ vssd1 vssd1 vccd1 vccd1 _0112_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2057_ dut.clkdiv_inst.counter\[12\] _0485_ vssd1 vssd1 vccd1 vccd1 _0487_ sky130_fd_sc_hd__and2_1
XFILLER_26_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2959_ dut.pwm_a_inst_y.pwm_out vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_32_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1290_ dut.pwm_a_inst_y.count_q\[0\] vssd1 vssd1 vccd1 vccd1 _0914_ sky130_fd_sc_hd__inv_2
XFILLER_0_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2813_ clknet_leaf_11_clk _0166_ net69 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.currentState\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_46_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1626_ _1212_ _1213_ dut.pwm_a_inst_y.count_q\[17\] dut.pwm_a_inst_y.count_q\[16\]
+ vssd1 vssd1 vccd1 vccd1 _1214_ sky130_fd_sc_hd__o211a_1
X_2675_ clknet_leaf_9_clk _0024_ net70 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_500hz\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_2744_ clknet_leaf_7_clk _0086_ net64 vssd1 vssd1 vccd1 vccd1 dut.microstep_y.ctr\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1557_ dut.actual_duty_y\[7\] _1145_ _1047_ vssd1 vssd1 vccd1 vccd1 _1146_ sky130_fd_sc_hd__a21bo_1
XFILLER_39_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1488_ _1068_ _1076_ vssd1 vssd1 vccd1 vccd1 _1077_ sky130_fd_sc_hd__nand2_1
XFILLER_52_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2109_ dut.spi.shift_reg_q\[3\] net20 _0520_ net216 _0524_ vssd1 vssd1 vccd1 vccd1
+ _0104_ sky130_fd_sc_hd__o221a_1
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2460_ net36 net37 _0805_ vssd1 vssd1 vccd1 vccd1 _0812_ sky130_fd_sc_hd__and3_1
XFILLER_5_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1411_ net13 _1013_ vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__nor2_1
X_2391_ net322 _0754_ net204 vssd1 vssd1 vccd1 vccd1 _0757_ sky130_fd_sc_hd__a21oi_1
X_1342_ dut.microstep_x.ctr\[19\] dut.microstep_x.ctr\[18\] dut.microstep_x.ctr\[21\]
+ dut.microstep_x.ctr\[20\] vssd1 vssd1 vccd1 vccd1 _0962_ sky130_fd_sc_hd__or4_1
XFILLER_3_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2727_ clknet_leaf_4_clk _0068_ net63 vssd1 vssd1 vccd1 vccd1 dut.microstep_y.ctr\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_1609_ dut.pwm_a_inst_y.count_q\[4\] _1181_ _1195_ _1197_ vssd1 vssd1 vccd1 vccd1
+ _1198_ sky130_fd_sc_hd__o211a_1
X_2589_ dut.ir_sensor_array.final_sensor_data\[24\] _0886_ dut.ir_sensor_array.final_sensor_data\[39\]
+ vssd1 vssd1 vccd1 vccd1 _0887_ sky130_fd_sc_hd__o21ba_1
X_2658_ clknet_leaf_24_clk _0129_ net73 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.bit_count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_57_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input1_A en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_02_92 vssd1 vssd1 vccd1 vccd1 team_02_92/HI gpio_oeb[8] sky130_fd_sc_hd__conb_1
XFILLER_42_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_8_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1891_ net166 _0946_ vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__xor2_1
X_1960_ dut.microstep_x.ctr\[1\] dut.microstep_x.ctr\[0\] net179 vssd1 vssd1 vccd1
+ vccd1 _0429_ sky130_fd_sc_hd__a21oi_1
XFILLER_52_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2443_ net41 _1133_ dut.actual_duty_y\[3\] vssd1 vssd1 vccd1 vccd1 _0795_ sky130_fd_sc_hd__o21ai_1
XFILLER_5_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2512_ dut.ir_sensor_array.final_sensor_data\[13\] dut.ir_sensor_array.final_sensor_data\[12\]
+ vssd1 vssd1 vccd1 vccd1 _0852_ sky130_fd_sc_hd__nor2_1
X_2374_ net226 _1004_ _0746_ vssd1 vssd1 vccd1 vccd1 _0147_ sky130_fd_sc_hd__o21a_1
X_1325_ dut.microstep_y.ctr\[3\] _0945_ vssd1 vssd1 vccd1 vccd1 _0946_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_62_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2090_ dut.pid_x.x_pid.last_error\[3\] _0509_ dut.clk_en vssd1 vssd1 vccd1 vccd1
+ _0098_ sky130_fd_sc_hd__mux2_1
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1943_ net196 _0419_ vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__xor2_1
X_1874_ dut.pwm_a_inst_x.count_q\[12\] _0301_ _0371_ dut.pwm_a_inst_x.count_q\[13\]
+ vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__a31o_1
X_2426_ _0768_ _0769_ _0774_ _0776_ vssd1 vssd1 vccd1 vccd1 _0778_ sky130_fd_sc_hd__o211a_1
X_1308_ dut.lcd1602.cnt_500hz\[1\] dut.lcd1602.cnt_500hz\[0\] dut.lcd1602.cnt_500hz\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0932_ sky130_fd_sc_hd__and3_1
XFILLER_56_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2357_ _0719_ _0721_ dut.microstep_x.clk_en vssd1 vssd1 vccd1 vccd1 _0739_ sky130_fd_sc_hd__o21a_1
X_2288_ net11 _0675_ vssd1 vssd1 vccd1 vccd1 _0676_ sky130_fd_sc_hd__nor2_1
XFILLER_60_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1590_ _1036_ _1178_ _1177_ vssd1 vssd1 vccd1 vccd1 _1179_ sky130_fd_sc_hd__a21o_1
XFILLER_53_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2211_ _0583_ _0604_ vssd1 vssd1 vccd1 vccd1 _0614_ sky130_fd_sc_hd__or2_1
X_2142_ dut.lcd1602.currentState\[0\] dut.lcd1602.currentState\[1\] vssd1 vssd1 vccd1
+ vccd1 _0545_ sky130_fd_sc_hd__nand2b_1
X_2073_ dut.clkdiv_inst.counter\[16\] dut.clkdiv_inst.counter\[13\] dut.clkdiv_inst.counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _0497_ sky130_fd_sc_hd__or3_1
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Left_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1926_ _0409_ vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__inv_2
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1857_ _0367_ vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__inv_2
X_1788_ _0302_ _0304_ vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_12_Left_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2409_ dut.lcd1602.currentState\[1\] net12 net18 vssd1 vssd1 vccd1 vccd1 _0163_ sky130_fd_sc_hd__mux2_1
XFILLER_55_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold60 dut.microstep_y.ctr\[26\] vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold71 _0103_ vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 dut.microstep_y.ctr\[9\] vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 dut.ir_sensor_array.final_sensor_data\[32\] vssd1 vssd1 vccd1 vccd1 net234
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_31_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2691_ clknet_leaf_16_clk dut.pwm_a_inst_y.count_d\[14\] net85 vssd1 vssd1 vccd1
+ vccd1 dut.pwm_a_inst_y.count_q\[14\] sky130_fd_sc_hd__dfrtp_2
X_1642_ _1224_ net21 _1223_ vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_y.count_d\[5\]
+ sky130_fd_sc_hd__and3b_1
X_1711_ net49 _0227_ _0226_ vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__a21oi_1
X_2760_ clknet_leaf_0_clk _0060_ net52 vssd1 vssd1 vccd1 vccd1 dut.microstep_x.ctr\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1573_ _1141_ _1159_ _1161_ vssd1 vssd1 vccd1 vccd1 _1162_ sky130_fd_sc_hd__a21o_1
XFILLER_39_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2125_ dut.spi.state_q\[1\] _0493_ _0532_ vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2056_ _0485_ _0486_ vssd1 vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__nor2_1
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1909_ dut.microstep_y.ctr\[9\] _0396_ net261 vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_32_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2958_ dut.pwm_a_inst_x.pwm_out vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
X_2889_ clknet_leaf_2_clk _0019_ net54 vssd1 vssd1 vccd1 vccd1 dut.clk_en sky130_fd_sc_hd__dfrtp_4
XFILLER_1_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput4 net4 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
XFILLER_63_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2743_ clknet_leaf_7_clk _0085_ net64 vssd1 vssd1 vccd1 vccd1 dut.microstep_y.ctr\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_2812_ clknet_leaf_11_clk _0165_ net71 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.currentState\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_16_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2674_ clknet_leaf_10_clk _0023_ net69 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_500hz\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_1625_ dut.pwm_a_inst_y.count_q\[10\] dut.pwm_a_inst_y.count_q\[11\] dut.pwm_a_inst_y.count_q\[8\]
+ _1037_ _1149_ vssd1 vssd1 vccd1 vccd1 _1213_ sky130_fd_sc_hd__a41o_1
X_1556_ _1059_ _1144_ _1051_ vssd1 vssd1 vccd1 vccd1 _1145_ sky130_fd_sc_hd__o21a_1
XFILLER_8_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1487_ _1066_ _1067_ dut.actual_duty_y\[2\] vssd1 vssd1 vccd1 vccd1 _1076_ sky130_fd_sc_hd__o21bai_1
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2108_ dut.data_in\[4\] _0515_ vssd1 vssd1 vccd1 vccd1 _0524_ sky130_fd_sc_hd__or2_1
XFILLER_39_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2039_ dut.clkdiv_inst.counter\[3\] _0969_ net265 vssd1 vssd1 vccd1 vccd1 _0477_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_22_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_15_Left_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1410_ dut.lcd1602.cnt_500hz\[1\] dut.lcd1602.cnt_500hz\[0\] vssd1 vssd1 vccd1 vccd1
+ _1013_ sky130_fd_sc_hd__xnor2_1
XFILLER_54_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2390_ dut.lcd1602.cnt_200ms\[13\] dut.lcd1602.cnt_200ms\[14\] _0754_ vssd1 vssd1
+ vccd1 vccd1 _0756_ sky130_fd_sc_hd__and3_1
XFILLER_3_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1341_ dut.microstep_x.ctr\[7\] dut.microstep_x.ctr\[9\] _0911_ dut.microstep_x.ctr\[6\]
+ vssd1 vssd1 vccd1 vccd1 _0961_ sky130_fd_sc_hd__or4b_1
XFILLER_36_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2726_ clknet_leaf_4_clk _0096_ net68 vssd1 vssd1 vccd1 vccd1 dut.microstep_y.ctr\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_1539_ _1126_ _1127_ vssd1 vssd1 vccd1 vccd1 _1128_ sky130_fd_sc_hd__nand2_1
X_1608_ dut.pwm_a_inst_y.count_q\[3\] _1193_ _1194_ _1196_ vssd1 vssd1 vccd1 vccd1
+ _1197_ sky130_fd_sc_hd__o2bb2a_1
X_2588_ dut.ir_sensor_array.final_sensor_data\[26\] _0885_ dut.ir_sensor_array.final_sensor_data\[25\]
+ vssd1 vssd1 vccd1 vccd1 _0886_ sky130_fd_sc_hd__o21ba_1
X_2657_ clknet_leaf_25_clk _0128_ net61 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.bit_count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_63_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xteam_02_93 vssd1 vssd1 vccd1 vccd1 team_02_93/HI gpio_oeb[9] sky130_fd_sc_hd__conb_1
XFILLER_27_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Left_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_92 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1890_ _0946_ _0386_ vssd1 vssd1 vccd1 vccd1 _0090_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2373_ _1005_ _1011_ vssd1 vssd1 vccd1 vccd1 _0746_ sky130_fd_sc_hd__nand2_1
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2442_ _1109_ _1133_ vssd1 vssd1 vccd1 vccd1 _0794_ sky130_fd_sc_hd__or2_1
X_2511_ _0848_ _0850_ vssd1 vssd1 vccd1 vccd1 _0851_ sky130_fd_sc_hd__nor2_1
XFILLER_5_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1324_ dut.microstep_y.ctr\[1\] dut.microstep_y.ctr\[0\] dut.microstep_y.ctr\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0945_ sky130_fd_sc_hd__and3_1
XFILLER_64_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2709_ clknet_leaf_21_clk dut.pwm_a_inst_x.count_d\[12\] net78 vssd1 vssd1 vccd1
+ vccd1 dut.pwm_a_inst_x.count_q\[12\] sky130_fd_sc_hd__dfrtp_2
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_36_Left_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_45_Left_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1942_ _0418_ _0419_ vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_16_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1873_ net221 _0376_ _0377_ vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_x.count_d\[12\]
+ sky130_fd_sc_hd__a21oi_1
X_2425_ _0774_ _0776_ _0768_ _0769_ vssd1 vssd1 vccd1 vccd1 _0777_ sky130_fd_sc_hd__a211oi_2
X_2356_ _0718_ _0719_ vssd1 vssd1 vccd1 vccd1 _0738_ sky130_fd_sc_hd__nand2_1
XFILLER_64_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1307_ net44 vssd1 vssd1 vccd1 vccd1 _0931_ sky130_fd_sc_hd__inv_2
X_2287_ dut.pid_x.x_pid.last_error\[2\] _0666_ _0512_ vssd1 vssd1 vccd1 vccd1 _0675_
+ sky130_fd_sc_hd__o21ba_1
XANTENNA_clkbuf_leaf_7_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_50 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2210_ _0582_ _0605_ _0609_ _0610_ _0612_ vssd1 vssd1 vccd1 vccd1 _0613_ sky130_fd_sc_hd__a311o_1
X_2141_ dut.lcd1602.currentState\[0\] dut.lcd1602.currentState\[1\] vssd1 vssd1 vccd1
+ vccd1 _0544_ sky130_fd_sc_hd__and2b_1
X_2072_ dut.clkdiv_inst.counter\[7\] dut.clkdiv_inst.counter\[9\] dut.clkdiv_inst.counter\[8\]
+ _0495_ dut.clkdiv_inst.counter\[10\] vssd1 vssd1 vccd1 vccd1 _0496_ sky130_fd_sc_hd__a41o_1
XFILLER_19_362 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1925_ dut.microstep_y.ctr\[15\] dut.microstep_y.ctr\[16\] _0405_ vssd1 vssd1 vccd1
+ vccd1 _0409_ sky130_fd_sc_hd__and3_1
XFILLER_34_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1787_ _0302_ _0304_ vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__nand2_1
X_1856_ dut.pwm_a_inst_x.count_q\[6\] _0327_ _0361_ vssd1 vssd1 vccd1 vccd1 _0367_
+ sky130_fd_sc_hd__and3_1
X_2408_ dut.lcd1602.currentState\[0\] _0570_ net18 vssd1 vssd1 vccd1 vccd1 _0162_
+ sky130_fd_sc_hd__mux2_1
XFILLER_39_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2339_ _0267_ _0268_ _0722_ _0719_ vssd1 vssd1 vccd1 vccd1 _0726_ sky130_fd_sc_hd__a31o_1
XFILLER_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold61 dut.lcd1602.cnt_200ms\[20\] vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 dut.spi.shift_reg_q\[2\] vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__dlygate4sd3_1
Xhold50 dut.lcd1602.cnt_500hz\[13\] vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 dut.microstep_y.ctr\[27\] vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 dut.clkdiv_inst.counter\[12\] vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_43_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2690_ clknet_leaf_17_clk dut.pwm_a_inst_y.count_d\[13\] net85 vssd1 vssd1 vccd1
+ vccd1 dut.pwm_a_inst_y.count_q\[13\] sky130_fd_sc_hd__dfrtp_2
X_1572_ _1039_ _1160_ vssd1 vssd1 vccd1 vccd1 _1161_ sky130_fd_sc_hd__nand2_1
X_1641_ dut.pwm_a_inst_y.count_q\[5\] dut.pwm_a_inst_y.count_q\[4\] _1219_ vssd1 vssd1
+ vccd1 vccd1 _1224_ sky130_fd_sc_hd__and3_1
X_1710_ _0226_ _0227_ vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__and2b_1
X_2124_ dut.spi.state_q\[0\] _0533_ _0532_ vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2055_ dut.clkdiv_inst.counter\[10\] _0484_ net267 vssd1 vssd1 vccd1 vccd1 _0486_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_24_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1908_ dut.microstep_y.ctr\[9\] dut.microstep_y.ctr\[10\] _0396_ vssd1 vssd1 vccd1
+ vccd1 _0398_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_32_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2888_ clknet_leaf_5_clk _0009_ net62 vssd1 vssd1 vccd1 vccd1 dut.clkdiv_inst.counter\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_1839_ dut.pwm_a_inst_x.count_q\[14\] _0356_ dut.pwm_a_inst_x.count_q\[17\] dut.pwm_a_inst_x.count_q\[16\]
+ dut.pwm_a_inst_x.count_q\[15\] vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__a2111oi_1
X_2957_ dut.ir_sensor_array.latch vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2715__123 vssd1 vssd1 vccd1 vccd1 _2715__123/HI net123 sky130_fd_sc_hd__conb_1
XFILLER_25_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput5 net5 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__buf_2
XFILLER_31_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_28_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2742_ clknet_leaf_7_clk _0084_ net64 vssd1 vssd1 vccd1 vccd1 dut.microstep_y.ctr\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_2811_ clknet_leaf_11_clk _0164_ net68 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.currentState\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1624_ dut.pwm_a_inst_y.count_q\[13\] dut.pwm_a_inst_y.count_q\[14\] dut.pwm_a_inst_y.count_q\[15\]
+ dut.pwm_a_inst_y.count_q\[12\] vssd1 vssd1 vccd1 vccd1 _1212_ sky130_fd_sc_hd__or4_1
X_2673_ clknet_leaf_11_clk _0022_ net69 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_500hz\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_1555_ _1072_ _1141_ _1143_ vssd1 vssd1 vccd1 vccd1 _1144_ sky130_fd_sc_hd__a21oi_1
X_2107_ dut.spi.shift_reg_q\[2\] net20 _0520_ net222 _0523_ vssd1 vssd1 vccd1 vccd1
+ _0103_ sky130_fd_sc_hd__o221a_1
XFILLER_39_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1486_ _1070_ _1074_ vssd1 vssd1 vccd1 vccd1 _1075_ sky130_fd_sc_hd__nand2_1
XFILLER_27_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_19_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_52_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2038_ dut.clkdiv_inst.counter\[3\] dut.clkdiv_inst.counter\[4\] _0969_ vssd1 vssd1
+ vccd1 vccd1 _0476_ sky130_fd_sc_hd__and3_1
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1340_ dut.microstep_x.ctr\[10\] dut.microstep_x.ctr\[12\] dut.microstep_x.ctr\[13\]
+ dut.microstep_x.ctr\[11\] vssd1 vssd1 vccd1 vccd1 _0960_ sky130_fd_sc_hd__or4bb_1
XFILLER_5_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_8_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2725_ clknet_leaf_4_clk _0095_ net68 vssd1 vssd1 vccd1 vccd1 dut.microstep_y.ctr\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_2656_ clknet_leaf_24_clk _0127_ net73 vssd1 vssd1 vccd1 vccd1 dut.ir_sensor_array.bit_count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1538_ _1119_ _1125_ vssd1 vssd1 vccd1 vccd1 _1127_ sky130_fd_sc_hd__or2_1
X_1607_ dut.pwm_a_inst_y.count_q\[0\] _0917_ _1191_ vssd1 vssd1 vccd1 vccd1 _1196_
+ sky130_fd_sc_hd__o21ai_1
X_1469_ _1055_ _1057_ vssd1 vssd1 vccd1 vccd1 _1058_ sky130_fd_sc_hd__nor2_1
X_2587_ dut.ir_sensor_array.final_sensor_data\[28\] _0884_ dut.ir_sensor_array.final_sensor_data\[27\]
+ vssd1 vssd1 vccd1 vccd1 _0885_ sky130_fd_sc_hd__o21ba_1
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xteam_02_94 vssd1 vssd1 vccd1 vccd1 team_02_94/HI gpio_oeb[10] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_40_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_5_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2510_ dut.ir_sensor_array.final_sensor_data\[24\] dut.ir_sensor_array.final_sensor_data\[27\]
+ dut.ir_sensor_array.final_sensor_data\[26\] dut.ir_sensor_array.final_sensor_data\[25\]
+ vssd1 vssd1 vccd1 vccd1 _0850_ sky130_fd_sc_hd__or4_1
X_2372_ _1004_ _0745_ net13 vssd1 vssd1 vccd1 vccd1 _0146_ sky130_fd_sc_hd__o21ai_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2441_ _0792_ vssd1 vssd1 vccd1 vccd1 _0793_ sky130_fd_sc_hd__inv_2
X_1323_ net35 _0909_ net28 vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__o21ai_1
XFILLER_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2639_ clknet_leaf_14_clk _0110_ net82 vssd1 vssd1 vccd1 vccd1 dut.spi.state_q\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_2708_ clknet_leaf_21_clk dut.pwm_a_inst_x.count_d\[11\] net78 vssd1 vssd1 vccd1
+ vccd1 dut.pwm_a_inst_x.count_q\[11\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1941_ dut.microstep_y.ctr\[22\] _0417_ vssd1 vssd1 vccd1 vccd1 _0419_ sky130_fd_sc_hd__and2_1
X_1872_ dut.pwm_a_inst_x.count_q\[12\] _0376_ net26 vssd1 vssd1 vccd1 vccd1 _0377_
+ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_16_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2424_ dut.pid_y.y_pid.last_error\[2\] dut.pid_y.y_pid.last_error\[1\] _0775_ vssd1
+ vssd1 vccd1 vccd1 _0776_ sky130_fd_sc_hd__o21bai_1
X_1306_ dut.microstep_x.clk_en vssd1 vssd1 vccd1 vccd1 _0930_ sky130_fd_sc_hd__inv_2
X_2355_ net47 dut.microstep_x.clk_en _0736_ _0737_ vssd1 vssd1 vccd1 vccd1 _0137_
+ sky130_fd_sc_hd__o22a_1
X_2286_ net11 vssd1 vssd1 vccd1 vccd1 _0674_ sky130_fd_sc_hd__inv_2
XFILLER_64_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2140_ dut.lcd1602.currentState\[4\] _0542_ _0541_ vssd1 vssd1 vccd1 vccd1 _0543_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_38_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2071_ dut.clkdiv_inst.counter\[3\] dut.clkdiv_inst.counter\[5\] dut.clkdiv_inst.counter\[4\]
+ dut.clkdiv_inst.counter\[6\] vssd1 vssd1 vccd1 vccd1 _0495_ sky130_fd_sc_hd__a31o_1
XFILLER_19_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1924_ dut.microstep_y.ctr\[15\] _0405_ _0408_ vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__o21a_1
X_1855_ _0366_ net27 _0365_ vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_x.count_d\[5\]
+ sky130_fd_sc_hd__and3b_1
X_1786_ _0290_ _0303_ vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__or2_1
X_2407_ net153 _0764_ vssd1 vssd1 vccd1 vccd1 _0161_ sky130_fd_sc_hd__xor2_1
XFILLER_44_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2269_ dut.ir_sensor_array.bit_count\[3\] _0939_ _0653_ vssd1 vssd1 vccd1 vccd1 _0660_
+ sky130_fd_sc_hd__and3_1
X_2338_ _0689_ _0722_ vssd1 vssd1 vccd1 vccd1 _0725_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_64_Left_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold40 dut.sdo_lcd vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 _0765_ vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 dut.pwm_a_inst_y.count_q\[15\] vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 dut.pwm_a_inst_y.count_q\[12\] vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 dut.lcd1602.cnt_200ms\[10\] vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 _0102_ vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_31_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1571_ dut.pwm_a_inst_y.count_q\[9\] _1038_ vssd1 vssd1 vccd1 vccd1 _1160_ sky130_fd_sc_hd__or2_1
X_1640_ dut.pwm_a_inst_y.count_q\[5\] _1221_ vssd1 vssd1 vccd1 vccd1 _1223_ sky130_fd_sc_hd__or2_1
X_2123_ dut.spi.state_q\[1\] _0974_ _0513_ vssd1 vssd1 vccd1 vccd1 _0533_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_6_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2054_ dut.clkdiv_inst.counter\[11\] dut.clkdiv_inst.counter\[10\] _0484_ vssd1 vssd1
+ vccd1 vccd1 _0485_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_24_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1907_ net245 _0396_ vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__xor2_1
X_2956_ net23 vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
X_2887_ clknet_leaf_5_clk _0008_ net62 vssd1 vssd1 vccd1 vccd1 dut.clkdiv_inst.counter\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_32_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1838_ _0301_ _0315_ dut.pwm_a_inst_x.count_q\[13\] dut.pwm_a_inst_x.count_q\[12\]
+ vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__a211o_1
X_1769_ _1271_ _0286_ _1258_ vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__a21oi_1
Xoutput6 net6 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__buf_2
XFILLER_36_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2672_ clknet_leaf_9_clk _0021_ net70 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.cnt_500hz\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_2810_ clknet_leaf_4_clk _0163_ net68 vssd1 vssd1 vccd1 vccd1 dut.lcd1602.currentState\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_2741_ clknet_leaf_6_clk _0083_ net62 vssd1 vssd1 vccd1 vccd1 dut.microstep_y.ctr\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1623_ _1206_ _1208_ _1211_ vssd1 vssd1 vccd1 vccd1 dut.pwm_a_inst_y.pwm_out sky130_fd_sc_hd__o21ba_1
X_1554_ _1059_ _1142_ vssd1 vssd1 vccd1 vccd1 _1143_ sky130_fd_sc_hd__or2_1
X_1485_ _1044_ _1067_ _1069_ vssd1 vssd1 vccd1 vccd1 _1074_ sky130_fd_sc_hd__or3_1
.ends

