* NGSPICE file created from team_04.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_1 abstract view
.subckt sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_2 abstract view
.subckt sky130_fd_sc_hd__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_4 abstract view
.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

.subckt team_04 ACK_I ADR_O[0] ADR_O[10] ADR_O[11] ADR_O[12] ADR_O[13] ADR_O[14] ADR_O[15]
+ ADR_O[16] ADR_O[17] ADR_O[18] ADR_O[19] ADR_O[1] ADR_O[20] ADR_O[21] ADR_O[22] ADR_O[23]
+ ADR_O[24] ADR_O[25] ADR_O[26] ADR_O[27] ADR_O[28] ADR_O[29] ADR_O[2] ADR_O[30] ADR_O[31]
+ ADR_O[3] ADR_O[4] ADR_O[5] ADR_O[6] ADR_O[7] ADR_O[8] ADR_O[9] CYC_O DAT_I[0] DAT_I[10]
+ DAT_I[11] DAT_I[12] DAT_I[13] DAT_I[14] DAT_I[15] DAT_I[16] DAT_I[17] DAT_I[18]
+ DAT_I[19] DAT_I[1] DAT_I[20] DAT_I[21] DAT_I[22] DAT_I[23] DAT_I[24] DAT_I[25] DAT_I[26]
+ DAT_I[27] DAT_I[28] DAT_I[29] DAT_I[2] DAT_I[30] DAT_I[31] DAT_I[3] DAT_I[4] DAT_I[5]
+ DAT_I[6] DAT_I[7] DAT_I[8] DAT_I[9] DAT_O[0] DAT_O[10] DAT_O[11] DAT_O[12] DAT_O[13]
+ DAT_O[14] DAT_O[15] DAT_O[16] DAT_O[17] DAT_O[18] DAT_O[19] DAT_O[1] DAT_O[20] DAT_O[21]
+ DAT_O[22] DAT_O[23] DAT_O[24] DAT_O[25] DAT_O[26] DAT_O[27] DAT_O[28] DAT_O[29]
+ DAT_O[2] DAT_O[30] DAT_O[31] DAT_O[3] DAT_O[4] DAT_O[5] DAT_O[6] DAT_O[7] DAT_O[8]
+ DAT_O[9] SEL_O[0] SEL_O[1] SEL_O[2] SEL_O[3] STB_O WE_O clk en gpio_in[0] gpio_in[10]
+ gpio_in[11] gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17]
+ gpio_in[18] gpio_in[19] gpio_in[1] gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23]
+ gpio_in[24] gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2]
+ gpio_in[30] gpio_in[31] gpio_in[32] gpio_in[33] gpio_in[3] gpio_in[4] gpio_in[5]
+ gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9] gpio_oeb[0] gpio_oeb[10] gpio_oeb[11]
+ gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15] gpio_oeb[16] gpio_oeb[17] gpio_oeb[18]
+ gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21] gpio_oeb[22] gpio_oeb[23] gpio_oeb[24]
+ gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28] gpio_oeb[29] gpio_oeb[2] gpio_oeb[30]
+ gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[3] gpio_oeb[4] gpio_oeb[5] gpio_oeb[6]
+ gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12]
+ gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19]
+ gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25]
+ gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31]
+ gpio_out[32] gpio_out[33] gpio_out[3] gpio_out[4] gpio_out[5] gpio_out[6] gpio_out[7]
+ gpio_out[8] gpio_out[9] nrst vccd1 vssd1
XFILLER_67_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09671_ net381 _03924_ _04506_ _03614_ vssd1 vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__a211o_1
X_06883_ net985 net938 vssd1 vssd1 vccd1 vccd1 _01719_ sky130_fd_sc_hd__and2_1
XANTENNA__07316__C net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08622_ _03453_ _03456_ _02387_ vssd1 vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__a21o_1
XANTENNA__08709__A _03263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09287__A1 _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08553_ datapath.rf.registers\[20\]\[0\] net964 net912 _01809_ vssd1 vssd1 vccd1
+ vccd1 _03389_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_124_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout162_A _05933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07504_ datapath.rf.registers\[16\]\[20\] _01707_ net929 vssd1 vssd1 vccd1 vccd1
+ _02340_ sky130_fd_sc_hd__and3_1
XANTENNA__07298__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08484_ datapath.rf.registers\[0\]\[1\] net869 _03309_ _03319_ vssd1 vssd1 vccd1
+ vccd1 _03320_ sky130_fd_sc_hd__o22ai_4
XFILLER_50_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07435_ datapath.rf.registers\[3\]\[22\] net770 net706 datapath.rf.registers\[10\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__a22o_1
XANTENNA__09039__A1 _02125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout427_A _05716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09099__X _03935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12043__B1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07366_ datapath.rf.registers\[3\]\[23\] net982 net927 vssd1 vssd1 vccd1 vccd1 _02202_
+ sky130_fd_sc_hd__and3_1
X_09105_ net344 _03806_ _03940_ vssd1 vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__a21oi_1
XFILLER_149_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08262__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07297_ datapath.rf.registers\[26\]\[25\] net780 net720 datapath.rf.registers\[20\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__a22o_1
XFILLER_136_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09036_ net368 _03631_ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__or2_1
XFILLER_124_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout796_A net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold340 datapath.rf.registers\[5\]\[15\] vssd1 vssd1 vccd1 vccd1 net1688 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10913__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold351 datapath.rf.registers\[7\]\[31\] vssd1 vssd1 vccd1 vccd1 net1699 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06899__A net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10357__B1 net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold362 datapath.rf.registers\[31\]\[19\] vssd1 vssd1 vccd1 vccd1 net1710 sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 datapath.rf.registers\[1\]\[8\] vssd1 vssd1 vccd1 vccd1 net1721 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold384 datapath.rf.registers\[14\]\[23\] vssd1 vssd1 vccd1 vccd1 net1732 sky130_fd_sc_hd__dlygate4sd3_1
Xhold395 datapath.rf.registers\[26\]\[20\] vssd1 vssd1 vccd1 vccd1 net1743 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout963_A net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout820 _01756_ vssd1 vssd1 vccd1 vccd1 net820 sky130_fd_sc_hd__buf_4
Xfanout831 _01748_ vssd1 vssd1 vccd1 vccd1 net831 sky130_fd_sc_hd__clkbuf_8
Xfanout842 net844 vssd1 vssd1 vccd1 vccd1 net842 sky130_fd_sc_hd__buf_2
XANTENNA__07507__B net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09938_ _04772_ _04773_ vssd1 vssd1 vccd1 vccd1 _04774_ sky130_fd_sc_hd__nand2_1
Xfanout853 net855 vssd1 vssd1 vccd1 vccd1 net853 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_144_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout864 _01726_ vssd1 vssd1 vccd1 vccd1 net864 sky130_fd_sc_hd__clkbuf_8
Xfanout875 _01723_ vssd1 vssd1 vccd1 vccd1 net875 sky130_fd_sc_hd__clkbuf_2
Xfanout886 _01716_ vssd1 vssd1 vccd1 vccd1 net886 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout751_X net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09869_ _04679_ _04694_ _04704_ _04681_ vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__o22a_1
Xfanout897 _01626_ vssd1 vssd1 vccd1 vccd1 net897 sky130_fd_sc_hd__clkbuf_4
Xhold1040 datapath.rf.registers\[11\]\[27\] vssd1 vssd1 vccd1 vccd1 net2388 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1051 datapath.rf.registers\[11\]\[18\] vssd1 vssd1 vccd1 vccd1 net2399 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout849_X net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11900_ _02680_ net657 vssd1 vssd1 vccd1 vccd1 _05964_ sky130_fd_sc_hd__nand2_1
Xhold1062 datapath.rf.registers\[18\]\[16\] vssd1 vssd1 vccd1 vccd1 net2410 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1073 datapath.rf.registers\[7\]\[29\] vssd1 vssd1 vccd1 vccd1 net2421 sky130_fd_sc_hd__dlygate4sd3_1
X_12880_ net241 net1593 net400 vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__mux2_1
Xhold1084 keypad.apps.app_c\[1\] vssd1 vssd1 vccd1 vccd1 net2432 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08619__A _02311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1095 datapath.rf.registers\[5\]\[19\] vssd1 vssd1 vccd1 vccd1 net2443 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11831_ _05302_ _05785_ _05794_ vssd1 vssd1 vccd1 vccd1 _05910_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_16_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ clknet_leaf_140_clk _01255_ net1097 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07289__B1 _02124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07828__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11762_ net1497 net145 net140 _02283_ vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__a22o_1
XFILLER_14_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13501_ clknet_leaf_145_clk _00311_ net1088 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08057__C net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10713_ datapath.multiplication_module.multiplicand_i\[1\] _03262_ net573 vssd1 vssd1
+ vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[2\] sky130_fd_sc_hd__mux2_1
XANTENNA__14038__SET_B net1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14481_ clknet_leaf_40_clk _01186_ net1140 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11693_ _04977_ net153 net148 net1427 vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__a22o_1
X_13432_ clknet_leaf_6_clk _00242_ net1068 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10644_ _05428_ _05429_ _05436_ vssd1 vssd1 vccd1 vccd1 _05464_ sky130_fd_sc_hd__or3_2
X_10575_ _03205_ _03263_ net559 net558 vssd1 vssd1 vccd1 vccd1 _05398_ sky130_fd_sc_hd__and4_1
X_13363_ clknet_leaf_36_clk _00173_ net1129 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08253__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13809__RESET_B net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12314_ _05595_ _06253_ _06290_ vssd1 vssd1 vccd1 vccd1 _06291_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07461__B1 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13294_ clknet_leaf_5_clk _00104_ net1069 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12337__A1 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09738__C1 _03614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12245_ _06238_ _06239_ vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_75_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12176_ _06195_ _06196_ vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__and2_1
XFILLER_150_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11127_ net233 net1639 net426 vssd1 vssd1 vccd1 vccd1 _00182_ sky130_fd_sc_hd__mux2_1
XFILLER_96_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08664__A_N _02284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11058_ net232 net2480 net430 vssd1 vssd1 vccd1 vccd1 _00118_ sky130_fd_sc_hd__mux2_1
XFILLER_67_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10009_ _04768_ _04793_ vssd1 vssd1 vccd1 vccd1 _04845_ sky130_fd_sc_hd__xnor2_1
XFILLER_76_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08248__B net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07819__A2 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12485__S net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14679_ clknet_leaf_126_clk _01384_ net1206 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08492__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06991__B _01816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07220_ datapath.rf.registers\[10\]\[26\] net879 net810 datapath.rf.registers\[13\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__a22o_1
XANTENNA__08229__C1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07151_ datapath.rf.registers\[28\]\[28\] net753 net663 datapath.rf.registers\[5\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__a22o_1
XANTENNA__09079__B _03914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07082_ datapath.rf.registers\[15\]\[29\] net799 net790 datapath.rf.registers\[18\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__a22o_1
XFILLER_145_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12514__A datapath.multiplication_module.multiplier_i\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08711__B _03418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07204__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout127 _06369_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__clkbuf_2
Xfanout138 net142 vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__buf_2
Xfanout149 net150 vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__clkbuf_2
XFILLER_87_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07984_ datapath.rf.registers\[22\]\[11\] net736 net670 datapath.rf.registers\[21\]\[11\]
+ _02819_ vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__a221o_2
XFILLER_86_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09723_ net609 _04557_ vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_126_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06935_ _01630_ _01639_ _01656_ net961 vssd1 vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__and4_1
XFILLER_28_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09654_ net644 _04486_ _04488_ _04489_ vssd1 vssd1 vccd1 vccd1 _04490_ sky130_fd_sc_hd__or4_1
X_06866_ net469 vssd1 vssd1 vccd1 vccd1 _01702_ sky130_fd_sc_hd__clkinv_4
XFILLER_83_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08605_ _02704_ _02726_ vssd1 vssd1 vccd1 vccd1 _03441_ sky130_fd_sc_hd__or2_1
X_09585_ net351 _04418_ _04420_ net360 vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__o211a_1
X_06797_ datapath.ru.latched_instruction\[22\] net1026 vssd1 vssd1 vccd1 vccd1 _01633_
+ sky130_fd_sc_hd__and2_1
XANTENNA_fanout165_X net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout544_A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08536_ datapath.rf.registers\[10\]\[0\] net881 net791 datapath.rf.registers\[18\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03372_ sky130_fd_sc_hd__a22o_1
XANTENNA__07630__X _02466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10275__C1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout711_A net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08467_ datapath.rf.registers\[19\]\[1\] net975 net927 vssd1 vssd1 vccd1 vccd1 _03303_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07997__B net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09680__A1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07418_ datapath.rf.registers\[10\]\[22\] net879 net810 datapath.rf.registers\[13\]\[22\]
+ _02253_ vssd1 vssd1 vccd1 vccd1 _02254_ sky130_fd_sc_hd__a221o_1
XANTENNA__07691__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08398_ datapath.rf.registers\[9\]\[2\] net988 net943 vssd1 vssd1 vccd1 vccd1 _03234_
+ sky130_fd_sc_hd__and3_1
XFILLER_137_801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_93_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12567__A1 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07349_ _02175_ _02181_ _02183_ _02184_ vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__or4_1
XANTENNA__08235__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1241_X net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07443__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10360_ _04846_ _04847_ vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__and2_1
XFILLER_137_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout799_X net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09019_ net340 _03706_ vssd1 vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__or2_1
X_10291_ _04429_ _04455_ vssd1 vssd1 vccd1 vccd1 _05127_ sky130_fd_sc_hd__xnor2_1
X_12030_ _05820_ _05852_ _05856_ _05847_ vssd1 vssd1 vccd1 vccd1 _06072_ sky130_fd_sc_hd__o211ai_1
XFILLER_3_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold170 screen.counter.currentCt\[14\] vssd1 vssd1 vccd1 vccd1 net1518 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold181 mmio.memload_or_instruction\[1\] vssd1 vssd1 vccd1 vccd1 net1529 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_151_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold192 datapath.rf.registers\[4\]\[23\] vssd1 vssd1 vccd1 vccd1 net1540 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout966_X net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08340__C net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_31_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout650 net651 vssd1 vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__clkbuf_2
Xfanout661 net663 vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__clkbuf_4
XFILLER_120_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout672 net674 vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__clkbuf_4
X_13981_ clknet_leaf_107_clk _00758_ net1221 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout683 net686 vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__buf_4
Xfanout694 net697 vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__clkbuf_8
XFILLER_74_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11474__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12932_ net304 net1972 net397 vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__mux2_1
XFILLER_74_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12863_ net207 net2097 net401 vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_46_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14602_ clknet_leaf_58_clk _01307_ net1167 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11814_ _01493_ net1015 net313 net334 datapath.ru.latched_instruction\[20\] vssd1
+ vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__a32o_1
XFILLER_73_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12794_ net174 net1905 net496 vssd1 vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__mux2_1
X_14533_ clknet_leaf_116_clk _01238_ net1187 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11745_ net1492 net143 net139 _03123_ vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__a22o_1
XANTENNA__10818__S net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08474__A2 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12007__B1 _06018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14464_ clknet_leaf_133_clk _01169_ net1111 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_11676_ _05136_ net154 net150 net1416 vssd1 vssd1 vccd1 vccd1 _00561_ sky130_fd_sc_hd__a22o_1
X_13415_ clknet_leaf_140_clk _00225_ net1093 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10627_ _05444_ _05445_ vssd1 vssd1 vccd1 vccd1 _05447_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_104_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14395_ clknet_leaf_37_clk _01100_ net1147 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_40_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13346_ clknet_leaf_152_clk _00156_ net1054 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_154_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10558_ _05315_ _05317_ _05326_ vssd1 vssd1 vccd1 vccd1 screen.register.controlFill
+ sky130_fd_sc_hd__or3_1
XANTENNA__08812__A _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13277_ clknet_leaf_149_clk _00087_ net1060 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10489_ screen.controlBus\[1\] _05314_ _05318_ screen.controlBus\[0\] vssd1 vssd1
+ vccd1 vccd1 _05319_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_90_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12228_ net2453 _06227_ net602 vssd1 vssd1 vccd1 vccd1 _06229_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_90_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_119_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12159_ net1275 _06161_ _06172_ vssd1 vssd1 vccd1 vccd1 _06186_ sky130_fd_sc_hd__and3_1
XFILLER_96_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_108_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11384__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06720_ _01441_ _01443_ _01502_ vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__or3_1
X_06651_ net1289 net1283 mmio.memload_or_instruction\[10\] vssd1 vssd1 vccd1 vccd1
+ _01490_ sky130_fd_sc_hd__or3b_2
XFILLER_25_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06582_ screen.counter.ct\[5\] vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__inv_2
XFILLER_52_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09370_ _04181_ _04182_ _04205_ vssd1 vssd1 vccd1 vccd1 _04206_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09111__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08321_ datapath.rf.registers\[12\]\[4\] net754 net679 datapath.rf.registers\[6\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03157_ sky130_fd_sc_hd__a22o_1
XFILLER_21_913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08465__A2 _01758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10728__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13104__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08252_ datapath.rf.registers\[25\]\[5\] net842 _03085_ _03087_ vssd1 vssd1 vccd1
+ vccd1 _03088_ sky130_fd_sc_hd__a211o_1
XANTENNA__07610__B net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07673__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07203_ datapath.rf.registers\[11\]\[27\] net711 net692 datapath.rf.registers\[13\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02039_ sky130_fd_sc_hd__a22o_1
XFILLER_119_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08183_ datapath.rf.registers\[24\]\[7\] net768 net728 datapath.rf.registers\[25\]\[7\]
+ _03018_ vssd1 vssd1 vccd1 vccd1 _03019_ sky130_fd_sc_hd__a221o_1
XANTENNA__08217__A2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12943__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_12_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_12_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_20_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xteam_04_1303 vssd1 vssd1 vccd1 vccd1 team_04_1303/HI gpio_oeb[12] sky130_fd_sc_hd__conb_1
XFILLER_9_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07134_ net874 _01965_ _01967_ _01969_ vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_119_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xteam_04_1314 vssd1 vssd1 vccd1 vccd1 team_04_1314/HI gpio_out[7] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_136_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xteam_04_1325 vssd1 vssd1 vccd1 vccd1 team_04_1325/HI gpio_out[29] sky130_fd_sc_hd__conb_1
Xteam_04_1336 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] team_04_1336/LO sky130_fd_sc_hd__conb_1
Xteam_04_1347 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] team_04_1347/LO sky130_fd_sc_hd__conb_1
X_07065_ datapath.rf.registers\[9\]\[30\] net704 net681 datapath.rf.registers\[6\]\[30\]
+ _01900_ vssd1 vssd1 vccd1 vccd1 _01901_ sky130_fd_sc_hd__a221o_1
XANTENNA__09178__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout494_A _06550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14232__Q datapath.multiplication_module.multiplier_i\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08925__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout661_A net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07967_ _02795_ _02800_ _02802_ vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__or3_4
XANTENNA_fanout759_A _01802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11294__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09706_ net358 _04355_ vssd1 vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__nor2_1
X_06918_ datapath.rf.registers\[6\]\[31\] net954 net933 vssd1 vssd1 vccd1 vccd1 _01754_
+ sky130_fd_sc_hd__and3_1
XFILLER_56_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07898_ datapath.rf.registers\[9\]\[12\] net886 net800 datapath.rf.registers\[15\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02734_ sky130_fd_sc_hd__a22o_1
XANTENNA__09350__B1 _02612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09637_ net578 _04471_ _04472_ _03607_ net606 vssd1 vssd1 vccd1 vccd1 _04473_ sky130_fd_sc_hd__a221oi_1
X_06849_ _01409_ _01583_ _01587_ _01410_ vssd1 vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__o22ai_1
XANTENNA__07504__C net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout926_A _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09568_ _02805_ net440 _04371_ net366 vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_26_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07801__A _02613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08519_ datapath.rf.registers\[20\]\[1\] net721 _03352_ _03353_ _03354_ vssd1 vssd1
+ vccd1 vccd1 _03355_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07113__C1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout714_X net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09499_ net648 _04332_ _04334_ vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_156_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13014__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11530_ screen.counter.ct\[3\] screen.counter.ct\[2\] vssd1 vssd1 vccd1 vccd1 _05754_
+ sky130_fd_sc_hd__nand2_1
XFILLER_8_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_137_Right_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10584__D _02980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12853__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11461_ net1681 net242 net408 vssd1 vssd1 vccd1 vccd1 _00499_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_122_Left_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13200_ clknet_leaf_57_clk _00010_ net1161 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07416__B1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10412_ net324 _04142_ vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__nor2_1
X_14180_ clknet_leaf_47_clk _00935_ net1175 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_136_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11392_ net1805 net250 net411 vssd1 vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__mux2_1
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11469__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13131_ net1609 net303 net384 vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__mux2_1
X_10343_ _05178_ net891 _04563_ vssd1 vssd1 vccd1 vccd1 _05179_ sky130_fd_sc_hd__or3b_1
XANTENNA__08351__B net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10274_ net1267 _03736_ vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__xnor2_1
X_13062_ net1569 net207 net388 vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12013_ _06039_ _06044_ _06056_ _06045_ vssd1 vssd1 vccd1 vccd1 _06057_ sky130_fd_sc_hd__o31a_1
XFILLER_78_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07195__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08392__A1 _03226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_131_Left_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout480 _06556_ vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__clkbuf_8
XFILLER_17_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout491 _06551_ vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__buf_4
X_13964_ clknet_leaf_104_clk _00742_ net1224 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12915_ net2099 net235 net484 vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10121__B _04057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13895_ clknet_leaf_43_clk net1368 net1150 vssd1 vssd1 vccd1 vccd1 keypad.decode.q2
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12846_ net244 net2401 net486 vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08807__A net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12777_ net254 net2065 net495 vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__mux2_1
XANTENNA__08447__A2 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08526__B net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14516_ clknet_leaf_20_clk _01221_ net1118 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11728_ net15 net1035 net1025 net1817 vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_140_Left_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14447_ clknet_leaf_23_clk _01152_ net1134 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_104_Right_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11659_ button\[3\] _05874_ vssd1 vssd1 vccd1 vccd1 _05879_ sky130_fd_sc_hd__and2_1
XFILLER_7_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14378_ clknet_leaf_59_clk _01083_ net1180 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold906 datapath.rf.registers\[23\]\[27\] vssd1 vssd1 vccd1 vccd1 net2254 sky130_fd_sc_hd__dlygate4sd3_1
Xhold917 datapath.rf.registers\[7\]\[30\] vssd1 vssd1 vccd1 vccd1 net2265 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11379__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13329_ clknet_leaf_40_clk _00139_ net1143 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold928 datapath.rf.registers\[17\]\[4\] vssd1 vssd1 vccd1 vccd1 net2276 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08080__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold939 datapath.rf.registers\[1\]\[30\] vssd1 vssd1 vccd1 vccd1 net2287 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_142_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08870_ _03704_ _03705_ net451 vssd1 vssd1 vccd1 vccd1 _03706_ sky130_fd_sc_hd__mux2_1
XFILLER_97_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07186__A2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07821_ datapath.rf.registers\[20\]\[14\] net839 _02638_ _02639_ _02640_ vssd1 vssd1
+ vccd1 vccd1 _02657_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09373__A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07752_ net612 _02587_ net564 vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__a21o_1
X_06703_ datapath.ru.latched_instruction\[16\] datapath.ru.latched_instruction\[17\]
+ datapath.ru.latched_instruction\[18\] datapath.ru.latched_instruction\[19\] vssd1
+ vssd1 vccd1 vccd1 _01542_ sky130_fd_sc_hd__or4_1
XFILLER_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12938__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07683_ datapath.rf.registers\[24\]\[17\] net858 _02499_ _02500_ _02506_ vssd1 vssd1
+ vccd1 vccd1 _02519_ sky130_fd_sc_hd__a2111oi_1
XFILLER_44_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09422_ net561 net442 _04195_ net364 vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__o211a_1
X_06634_ datapath.ru.latched_instruction\[2\] _01444_ _01462_ datapath.ru.latched_instruction\[3\]
+ _01472_ vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__o221a_1
XANTENNA__08717__A _03205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09353_ _04130_ _04131_ net459 vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__a21o_1
X_06565_ datapath.ru.zero_multi1 vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_23_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout242_A _05605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08436__B net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08304_ datapath.rf.registers\[11\]\[4\] net882 net794 datapath.rf.registers\[31\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03140_ sky130_fd_sc_hd__a22o_1
XANTENNA__07646__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09284_ _03448_ _04119_ vssd1 vssd1 vccd1 vccd1 _04120_ sky130_fd_sc_hd__xor2_2
XANTENNA__07110__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08235_ datapath.rf.registers\[18\]\[6\] net722 net698 datapath.rf.registers\[23\]\[6\]
+ _03068_ vssd1 vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__a221o_1
XFILLER_20_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout507_A net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1249_A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08166_ datapath.rf.registers\[20\]\[7\] net840 net816 datapath.rf.registers\[21\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03002_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_151_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11289__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07117_ _01939_ _01940_ _01947_ _01952_ vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__or4_1
XFILLER_106_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08097_ _02923_ _02930_ _02932_ vssd1 vssd1 vccd1 vccd1 _02933_ sky130_fd_sc_hd__and3_2
X_07048_ datapath.rf.registers\[3\]\[30\] net802 net797 datapath.rf.registers\[29\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__a22o_1
Xclkload90 clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 clkload90/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_54_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout876_A net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout497_X net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1204_X net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07177__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout664_X net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08999_ _01980_ _02025_ net442 vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__mux2_1
XFILLER_75_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13009__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12458__B1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09323__B1 _02567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10579__D _02364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout831_X net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10961_ datapath.mulitply_result\[0\] net598 net620 vssd1 vssd1 vccd1 vccd1 _05699_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__12848__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout929_X net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12700_ _01432_ _01434_ vssd1 vssd1 vccd1 vccd1 _06530_ sky130_fd_sc_hd__nor2_2
XANTENNA__07885__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13680_ clknet_leaf_24_clk _00490_ net1160 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10892_ net902 _05638_ vssd1 vssd1 vccd1 vccd1 _05639_ sky130_fd_sc_hd__nand2_2
XANTENNA__08627__A _02125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12631_ _06461_ _06465_ _06467_ vssd1 vssd1 vccd1 vccd1 _06473_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08346__B net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07637__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12562_ _06411_ _06412_ _06410_ vssd1 vssd1 vccd1 vccd1 _06415_ sky130_fd_sc_hd__o21ba_1
XANTENNA__07101__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14301_ clknet_leaf_145_clk _01006_ net1085 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11513_ net1280 net1275 net1271 _05335_ vssd1 vssd1 vccd1 vccd1 _05738_ sky130_fd_sc_hd__and4_1
XANTENNA__11984__A2 _05778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10892__A net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12493_ net248 net2140 net506 vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__mux2_1
XFILLER_8_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14232_ clknet_leaf_123_clk datapath.multiplication_module.multiplier_i_n\[0\] net1215
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i\[0\] sky130_fd_sc_hd__dfrtp_2
X_11444_ net1676 net209 net409 vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__mux2_1
XFILLER_137_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11199__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14163_ clknet_leaf_66_clk _00918_ net1237 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08062__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11375_ _05514_ _05724_ vssd1 vssd1 vccd1 vccd1 _05729_ sky130_fd_sc_hd__or2_1
XFILLER_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13114_ net235 net1735 net471 vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__mux2_1
X_10326_ _04207_ _04583_ vssd1 vssd1 vccd1 vccd1 _05162_ sky130_fd_sc_hd__and2_1
X_14094_ clknet_leaf_122_clk _00860_ net1201 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07409__C net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13045_ net243 net2504 net475 vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__mux2_1
X_10257_ _04855_ _05092_ vssd1 vssd1 vccd1 vccd1 _05093_ sky130_fd_sc_hd__or2_1
Xfanout1220 net1221 vssd1 vssd1 vccd1 vccd1 net1220 sky130_fd_sc_hd__clkbuf_4
Xfanout1231 net1262 vssd1 vssd1 vccd1 vccd1 net1231 sky130_fd_sc_hd__buf_2
Xfanout1242 net1243 vssd1 vssd1 vccd1 vccd1 net1242 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14023__RESET_B net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10188_ net894 _04146_ vssd1 vssd1 vccd1 vccd1 _05024_ sky130_fd_sc_hd__nor2_1
XFILLER_79_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1253 net1261 vssd1 vssd1 vccd1 vccd1 net1253 sky130_fd_sc_hd__clkbuf_2
Xfanout1264 datapath.PC\[24\] vssd1 vssd1 vccd1 vccd1 net1264 sky130_fd_sc_hd__buf_2
Xfanout1275 screen.counter.ct\[10\] vssd1 vssd1 vccd1 vccd1 net1275 sky130_fd_sc_hd__buf_2
Xfanout1286 net1290 vssd1 vssd1 vccd1 vccd1 net1286 sky130_fd_sc_hd__buf_2
XANTENNA__12449__B1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09314__B1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13947_ clknet_leaf_110_clk _00725_ net1222 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12758__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07876__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11672__A1 _05270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13878_ clknet_leaf_53_clk _00682_ net1183 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[22\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07340__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06983__C _01800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12829_ _05518_ _05732_ vssd1 vssd1 vccd1 vccd1 _06552_ sky130_fd_sc_hd__or2_4
XANTENNA__09617__A1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_150_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_150_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12493__S net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08020_ datapath.rf.registers\[0\]\[10\] net868 _02855_ vssd1 vssd1 vccd1 vccd1 _02856_
+ sky130_fd_sc_hd__o21a_2
XTAP_TAPCELL_ROW_116_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13886__Q datapath.ru.latched_instruction\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11727__A2 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold703 datapath.rf.registers\[19\]\[15\] vssd1 vssd1 vccd1 vccd1 net2051 sky130_fd_sc_hd__dlygate4sd3_1
Xhold714 datapath.rf.registers\[19\]\[18\] vssd1 vssd1 vccd1 vccd1 net2062 sky130_fd_sc_hd__dlygate4sd3_1
Xhold725 datapath.rf.registers\[31\]\[6\] vssd1 vssd1 vccd1 vccd1 net2073 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold736 datapath.rf.registers\[15\]\[9\] vssd1 vssd1 vccd1 vccd1 net2084 sky130_fd_sc_hd__dlygate4sd3_1
Xhold747 datapath.rf.registers\[8\]\[18\] vssd1 vssd1 vccd1 vccd1 net2095 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold758 datapath.rf.registers\[27\]\[22\] vssd1 vssd1 vccd1 vccd1 net2106 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_wire465_X net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09971_ _04746_ _04748_ _04804_ _04745_ _04742_ vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__a311o_1
Xhold769 datapath.rf.registers\[16\]\[26\] vssd1 vssd1 vccd1 vccd1 net2117 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08922_ _03595_ _03757_ net578 vssd1 vssd1 vccd1 vccd1 _03758_ sky130_fd_sc_hd__o21a_1
XANTENNA__07159__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08853_ _03687_ _03688_ net449 vssd1 vssd1 vccd1 vccd1 _03689_ sky130_fd_sc_hd__mux2_1
XANTENNA__11409__Y _05731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout192_A _05659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06906__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07804_ datapath.rf.registers\[5\]\[14\] net945 net933 vssd1 vssd1 vccd1 vccd1 _02640_
+ sky130_fd_sc_hd__and3_1
X_08784_ _03617_ net332 _03613_ vssd1 vssd1 vccd1 vccd1 _03620_ sky130_fd_sc_hd__o21ai_1
XFILLER_85_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09305__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07735_ datapath.rf.registers\[16\]\[16\] net738 net687 datapath.rf.registers\[31\]\[16\]
+ _02570_ vssd1 vssd1 vccd1 vccd1 _02571_ sky130_fd_sc_hd__a221o_1
XFILLER_38_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07666_ datapath.rf.registers\[21\]\[17\] net947 net925 vssd1 vssd1 vccd1 vccd1 _02502_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07331__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09405_ _03444_ _04240_ vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__xor2_1
X_06617_ net1290 net1281 mmio.memload_or_instruction\[22\] vssd1 vssd1 vccd1 vccd1
+ _01456_ sky130_fd_sc_hd__nor3b_2
XANTENNA__10871__C1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout624_A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07597_ datapath.rf.registers\[26\]\[19\] net780 net720 datapath.rf.registers\[20\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__a22o_1
XANTENNA__07619__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09336_ net319 _03942_ vssd1 vssd1 vccd1 vccd1 _04172_ sky130_fd_sc_hd__nor2_1
XFILLER_139_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10916__S net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09267_ _04037_ _04038_ net459 vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout412_X net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_141_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_141_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11601__A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08218_ datapath.rf.registers\[17\]\[6\] net849 net807 datapath.rf.registers\[27\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03054_ sky130_fd_sc_hd__a22o_1
XANTENNA__06842__B2 datapath.ru.latched_instruction\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_5_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09198_ _04028_ _04033_ net376 vssd1 vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__mux2_1
XFILLER_153_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08149_ datapath.rf.registers\[30\]\[7\] net976 net919 vssd1 vssd1 vccd1 vccd1 _02985_
+ sky130_fd_sc_hd__and3_1
XFILLER_146_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09241__C1 _03673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10217__A net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07398__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11160_ net237 net2620 net532 vssd1 vssd1 vccd1 vccd1 _00213_ sky130_fd_sc_hd__mux2_1
XFILLER_122_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout781_X net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout879_X net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10111_ _03744_ _04946_ net1041 vssd1 vssd1 vccd1 vccd1 _04947_ sky130_fd_sc_hd__a21oi_1
X_11091_ net219 net2019 net535 vssd1 vssd1 vccd1 vccd1 _00148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10042_ _04833_ _04877_ vssd1 vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__nor2_1
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold30 columns.count\[3\] vssd1 vssd1 vccd1 vccd1 net1378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 screen.controlBus\[22\] vssd1 vssd1 vccd1 vccd1 net1389 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 mmio.memload_or_instruction\[4\] vssd1 vssd1 vccd1 vccd1 net1400 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold63 net40 vssd1 vssd1 vccd1 vccd1 net1411 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 net47 vssd1 vssd1 vccd1 vccd1 net1422 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold85 screen.controlBus\[16\] vssd1 vssd1 vccd1 vccd1 net1433 sky130_fd_sc_hd__dlygate4sd3_1
X_13801_ clknet_leaf_52_clk _00610_ net1184 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[22\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold96 datapath.multiplication_module.multiplier_i\[1\] vssd1 vssd1 vccd1 vccd1 net1444
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07570__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input18_A DAT_I[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11993_ _06037_ net1438 _06017_ vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__mux2_1
XANTENNA__11482__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13732_ clknet_leaf_18_clk _00542_ net1119 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10457__A2 _05073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07858__B1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10944_ _01466_ net619 _05683_ vssd1 vssd1 vccd1 vccd1 _05684_ sky130_fd_sc_hd__a21oi_4
XFILLER_16_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07322__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13663_ clknet_leaf_12_clk _00473_ net1082 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10875_ datapath.PC\[21\] _05617_ vssd1 vssd1 vccd1 vccd1 _05624_ sky130_fd_sc_hd__xnor2_1
XFILLER_44_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12614_ _06456_ _06457_ _06458_ vssd1 vssd1 vccd1 vccd1 _06459_ sky130_fd_sc_hd__or3_1
X_13594_ clknet_leaf_146_clk _00404_ net1091 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08283__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12545_ datapath.mulitply_result\[6\] datapath.multiplication_module.multiplicand_i\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06401_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_132_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_132_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10826__S net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12476_ _05689_ _05724_ vssd1 vssd1 vccd1 vccd1 _06370_ sky130_fd_sc_hd__or2_1
XANTENNA__11709__A2 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14215_ clknet_leaf_48_clk datapath.multiplication_module.multiplicand_i_n\[26\]
+ net1175 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11427_ net241 net2224 net516 vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__mux2_1
XANTENNA__08035__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_5 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07389__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12382__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14146_ clknet_leaf_37_clk _00903_ net1137 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11358_ net247 net2169 net519 vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__mux2_1
XFILLER_152_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08820__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10309_ net222 _05144_ net1294 vssd1 vssd1 vccd1 vccd1 _05145_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_111_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14077_ clknet_leaf_111_clk _00844_ net1199 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_111_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11289_ net249 net2446 net523 vssd1 vssd1 vccd1 vccd1 _00337_ sky130_fd_sc_hd__mux2_1
XANTENNA__09535__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13028_ _05518_ _06558_ vssd1 vssd1 vccd1 vccd1 _06559_ sky130_fd_sc_hd__or2_1
XFILLER_140_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10145__B2 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08889__A2 _01859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1050 net1051 vssd1 vssd1 vccd1 vccd1 net1050 sky130_fd_sc_hd__clkbuf_2
Xfanout1061 net1066 vssd1 vssd1 vccd1 vccd1 net1061 sky130_fd_sc_hd__buf_2
Xfanout1072 net1074 vssd1 vssd1 vccd1 vccd1 net1072 sky130_fd_sc_hd__clkbuf_4
XFILLER_13_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1083 net1084 vssd1 vssd1 vccd1 vccd1 net1083 sky130_fd_sc_hd__buf_2
Xfanout1094 net1096 vssd1 vssd1 vccd1 vccd1 net1094 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07561__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12488__S net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11392__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07520_ datapath.rf.registers\[7\]\[20\] net818 _02341_ _02346_ _02347_ vssd1 vssd1
+ vccd1 vccd1 _02356_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13173__A datapath.rf.registers\[0\]\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07849__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07451_ _02286_ vssd1 vssd1 vccd1 vccd1 _02287_ sky130_fd_sc_hd__inv_2
XFILLER_23_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07382_ _02217_ vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_33_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09121_ _03836_ _03956_ net374 vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08274__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_123_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_123_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_31_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13112__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09052_ _03883_ _03887_ net353 vssd1 vssd1 vccd1 vccd1 _03888_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_98_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08003_ datapath.rf.registers\[2\]\[10\] net984 net950 vssd1 vssd1 vccd1 vccd1 _02839_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08026__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12951__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold500 datapath.rf.registers\[13\]\[28\] vssd1 vssd1 vccd1 vccd1 net1848 sky130_fd_sc_hd__dlygate4sd3_1
Xhold511 datapath.rf.registers\[29\]\[6\] vssd1 vssd1 vccd1 vccd1 net1859 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10908__B1 _05651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout205_A _05641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold522 datapath.rf.registers\[1\]\[7\] vssd1 vssd1 vccd1 vccd1 net1870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold533 datapath.rf.registers\[15\]\[15\] vssd1 vssd1 vccd1 vccd1 net1881 sky130_fd_sc_hd__dlygate4sd3_1
Xhold544 datapath.rf.registers\[12\]\[13\] vssd1 vssd1 vccd1 vccd1 net1892 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10384__A1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold555 datapath.rf.registers\[17\]\[9\] vssd1 vssd1 vccd1 vccd1 net1903 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold566 datapath.rf.registers\[21\]\[18\] vssd1 vssd1 vccd1 vccd1 net1914 sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 datapath.rf.registers\[3\]\[13\] vssd1 vssd1 vccd1 vccd1 net1925 sky130_fd_sc_hd__dlygate4sd3_1
Xhold588 datapath.rf.registers\[13\]\[12\] vssd1 vssd1 vccd1 vccd1 net1936 sky130_fd_sc_hd__dlygate4sd3_1
X_09954_ _04775_ _04789_ vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__nand2b_1
Xhold599 datapath.rf.registers\[10\]\[29\] vssd1 vssd1 vccd1 vccd1 net1947 sky130_fd_sc_hd__dlygate4sd3_1
X_08905_ datapath.PC\[15\] _03740_ vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__or2_1
XFILLER_98_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09885_ datapath.PC\[24\] datapath.PC\[25\] net1263 datapath.PC\[27\] net594 vssd1
+ vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__o41a_1
Xhold1200 mmio.memload_or_instruction\[26\] vssd1 vssd1 vccd1 vccd1 net2548 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout574_A net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1211 datapath.mulitply_result\[25\] vssd1 vssd1 vccd1 vccd1 net2559 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_146_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1222 datapath.rf.registers\[10\]\[24\] vssd1 vssd1 vccd1 vccd1 net2570 sky130_fd_sc_hd__dlygate4sd3_1
X_08836_ _03171_ net967 _03671_ vssd1 vssd1 vccd1 vccd1 _03672_ sky130_fd_sc_hd__mux2_1
Xhold1233 datapath.rf.registers\[3\]\[9\] vssd1 vssd1 vccd1 vccd1 net2581 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1244 datapath.mulitply_result\[23\] vssd1 vssd1 vccd1 vccd1 net2592 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1255 datapath.rf.registers\[26\]\[25\] vssd1 vssd1 vccd1 vccd1 net2603 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1266 datapath.rf.registers\[25\]\[11\] vssd1 vssd1 vccd1 vccd1 net2614 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1277 datapath.rf.registers\[23\]\[10\] vssd1 vssd1 vccd1 vccd1 net2625 sky130_fd_sc_hd__dlygate4sd3_1
X_08767_ net651 net642 _01606_ vssd1 vssd1 vccd1 vccd1 _03603_ sky130_fd_sc_hd__o21a_1
XFILLER_38_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1288 screen.controlBus\[1\] vssd1 vssd1 vccd1 vccd1 net2636 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1299 datapath.rf.registers\[27\]\[25\] vssd1 vssd1 vccd1 vccd1 net2647 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout839_A net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07718_ datapath.rf.registers\[8\]\[16\] net876 net832 datapath.rf.registers\[30\]\[16\]
+ _02553_ vssd1 vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__a221o_1
XANTENNA__10439__A2 _04338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08698_ _02857_ _02879_ vssd1 vssd1 vccd1 vccd1 _03534_ sky130_fd_sc_hd__nor2_1
XANTENNA__07304__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07649_ _02478_ _02480_ _02482_ _02484_ vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__or4_1
XANTENNA__07512__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout627_X net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10660_ _05472_ _05476_ vssd1 vssd1 vccd1 vccd1 _05479_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_62_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09319_ _04064_ _04154_ net372 vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__mux2_1
XANTENNA__12061__A1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10591_ _02239_ _02283_ _02331_ _02385_ vssd1 vssd1 vccd1 vccd1 _05414_ sky130_fd_sc_hd__or4_1
XANTENNA__12061__B2 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_114_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_114_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_11_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13022__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10072__B1 net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12330_ _04876_ _05624_ net230 vssd1 vssd1 vccd1 vccd1 _06302_ sky130_fd_sc_hd__mux2_1
XANTENNA__06815__B2 datapath.ru.latched_instruction\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout996_X net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08343__C net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10592__D _02587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08017__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12261_ net636 _04838_ vssd1 vssd1 vccd1 vccd1 _06251_ sky130_fd_sc_hd__or2_1
XANTENNA__12861__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14000_ clknet_leaf_114_clk _00777_ net1195 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_11212_ net298 net1938 net526 vssd1 vssd1 vccd1 vccd1 _00262_ sky130_fd_sc_hd__mux2_1
X_12192_ screen.counter.currentCt\[0\] _06167_ vssd1 vssd1 vccd1 vccd1 _06206_ sky130_fd_sc_hd__nand2b_1
Xoutput42 net42 vssd1 vssd1 vccd1 vccd1 ADR_O[11] sky130_fd_sc_hd__buf_2
XFILLER_150_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput53 net53 vssd1 vssd1 vccd1 vccd1 ADR_O[21] sky130_fd_sc_hd__buf_2
X_11143_ net288 net1884 net533 vssd1 vssd1 vccd1 vccd1 _00196_ sky130_fd_sc_hd__mux2_1
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 ADR_O[31] sky130_fd_sc_hd__buf_2
XFILLER_1_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 DAT_O[11] sky130_fd_sc_hd__buf_2
XANTENNA__09517__A0 _02804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput86 net86 vssd1 vssd1 vccd1 vccd1 DAT_O[21] sky130_fd_sc_hd__buf_2
XANTENNA__07791__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07256__A _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput97 net97 vssd1 vssd1 vccd1 vccd1 DAT_O[31] sky130_fd_sc_hd__buf_2
XANTENNA__10127__A1 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11074_ net259 net1663 net536 vssd1 vssd1 vccd1 vccd1 _00131_ sky130_fd_sc_hd__mux2_1
XFILLER_1_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10025_ _04746_ _04805_ vssd1 vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__xor2_2
XFILLER_37_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07543__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11976_ _05323_ _05767_ vssd1 vssd1 vccd1 vccd1 _06021_ sky130_fd_sc_hd__and2_1
XFILLER_60_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13715_ clknet_leaf_35_clk _00525_ net1129 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10927_ datapath.mulitply_result\[28\] net597 net617 vssd1 vssd1 vccd1 vccd1 _05669_
+ sky130_fd_sc_hd__a21o_1
XFILLER_72_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14695_ clknet_leaf_137_clk _01400_ net1089 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_13646_ clknet_leaf_5_clk _00456_ net1056 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10858_ _01453_ net652 _05609_ vssd1 vssd1 vccd1 vccd1 _05610_ sky130_fd_sc_hd__o21a_2
XANTENNA__08256__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12052__A1 _05335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_105_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_105_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13577_ clknet_leaf_62_clk _00387_ net1234 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10789_ _05550_ vssd1 vssd1 vccd1 vccd1 _05551_ sky130_fd_sc_hd__inv_2
XFILLER_40_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06980__D _01666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12528_ _06385_ _06386_ vssd1 vssd1 vccd1 vccd1 _06387_ sky130_fd_sc_hd__nor2_1
XFILLER_145_526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12459_ net164 _05966_ net126 screen.register.currentXbus\[15\] vssd1 vssd1 vccd1
+ vccd1 _00861_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12771__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06989__B _01637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11387__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14129_ clknet_leaf_22_clk _00886_ net1157 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_93_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout309 _06246_ vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__clkbuf_4
XFILLER_141_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07166__A _02001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06951_ net611 net596 vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__nand2_2
XFILLER_39_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09670_ net377 _04155_ _04505_ net330 vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__o211a_1
XFILLER_95_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_863 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06882_ _01629_ _01639_ _01656_ net962 vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__and4_1
XANTENNA__07534__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08731__A1 _02912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08621_ _02333_ _03456_ _03455_ vssd1 vssd1 vccd1 vccd1 _03457_ sky130_fd_sc_hd__o21a_1
XANTENNA__08268__Y _03104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13107__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08709__B _03296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08552_ datapath.rf.registers\[14\]\[0\] net777 _03385_ _03386_ _03387_ vssd1 vssd1
+ vccd1 vccd1 _03388_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_124_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07503_ datapath.rf.registers\[26\]\[20\] net973 net937 vssd1 vssd1 vccd1 vccd1 _02339_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12946__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08483_ _03311_ _03313_ _03314_ _03318_ vssd1 vssd1 vccd1 vccd1 _03319_ sky130_fd_sc_hd__or4_2
XANTENNA__09692__C1 _03614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07434_ _02268_ _02269_ vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__or2_1
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_8_0_clk_X clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07365_ datapath.rf.registers\[19\]\[23\] net974 net927 vssd1 vssd1 vccd1 vccd1 _02201_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12448__A1_N net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09104_ net340 _03811_ _03812_ vssd1 vssd1 vccd1 vccd1 _03940_ sky130_fd_sc_hd__and3_1
X_07296_ datapath.rf.registers\[22\]\[25\] net736 net666 datapath.rf.registers\[15\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__a22o_1
XFILLER_108_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09035_ net608 _03867_ vssd1 vssd1 vccd1 vccd1 _03871_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout1231_A net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold330 datapath.rf.registers\[13\]\[6\] vssd1 vssd1 vccd1 vccd1 net1678 sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 datapath.rf.registers\[12\]\[18\] vssd1 vssd1 vccd1 vccd1 net1689 sky130_fd_sc_hd__dlygate4sd3_1
Xhold352 datapath.rf.registers\[12\]\[21\] vssd1 vssd1 vccd1 vccd1 net1700 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout691_A _01824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11297__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06899__B _01707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold363 datapath.rf.registers\[4\]\[7\] vssd1 vssd1 vccd1 vccd1 net1711 sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 datapath.rf.registers\[7\]\[26\] vssd1 vssd1 vccd1 vccd1 net1722 sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 datapath.rf.registers\[7\]\[19\] vssd1 vssd1 vccd1 vccd1 net1733 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 datapath.rf.registers\[18\]\[27\] vssd1 vssd1 vccd1 vccd1 net1744 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_120_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout810 net812 vssd1 vssd1 vccd1 vccd1 net810 sky130_fd_sc_hd__clkbuf_8
Xfanout821 net823 vssd1 vssd1 vccd1 vccd1 net821 sky130_fd_sc_hd__buf_4
XANTENNA__07773__A2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08970__A1 _03805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout832 net835 vssd1 vssd1 vccd1 vccd1 net832 sky130_fd_sc_hd__clkbuf_8
X_09937_ datapath.PC\[5\] _03124_ vssd1 vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__or2_1
XANTENNA__10109__A1 _04118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout843 net844 vssd1 vssd1 vccd1 vccd1 net843 sky130_fd_sc_hd__buf_4
XANTENNA__07507__C net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13761__RESET_B net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout854 net855 vssd1 vssd1 vccd1 vccd1 net854 sky130_fd_sc_hd__clkbuf_8
Xfanout865 _01726_ vssd1 vssd1 vccd1 vccd1 net865 sky130_fd_sc_hd__clkbuf_4
Xfanout876 net878 vssd1 vssd1 vccd1 vccd1 net876 sky130_fd_sc_hd__clkbuf_8
Xfanout887 net889 vssd1 vssd1 vccd1 vccd1 net887 sky130_fd_sc_hd__buf_4
X_09868_ _04677_ _04696_ _04700_ _04703_ vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__o211a_1
Xhold1030 datapath.rf.registers\[15\]\[19\] vssd1 vssd1 vccd1 vccd1 net2378 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout898 _01626_ vssd1 vssd1 vccd1 vccd1 net898 sky130_fd_sc_hd__buf_2
XFILLER_133_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1041 datapath.rf.registers\[29\]\[13\] vssd1 vssd1 vccd1 vccd1 net2389 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07525__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08819_ net992 _03643_ vssd1 vssd1 vccd1 vccd1 _03655_ sky130_fd_sc_hd__nor2_1
Xhold1052 datapath.rf.registers\[27\]\[10\] vssd1 vssd1 vccd1 vccd1 net2400 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1063 datapath.multiplication_module.multiplicand_i\[14\] vssd1 vssd1 vccd1 vccd1
+ net2411 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1074 datapath.rf.registers\[17\]\[27\] vssd1 vssd1 vccd1 vccd1 net2422 sky130_fd_sc_hd__dlygate4sd3_1
X_09799_ net348 _04251_ net575 vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout744_X net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1085 _00659_ vssd1 vssd1 vccd1 vccd1 net2433 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13017__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11830_ _01423_ net1273 _05299_ _05908_ vssd1 vssd1 vccd1 vccd1 _05909_ sky130_fd_sc_hd__or4b_1
Xhold1096 datapath.rf.registers\[9\]\[25\] vssd1 vssd1 vccd1 vccd1 net2444 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09278__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ net1503 net145 net140 _02331_ vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__a22o_1
XANTENNA__12856__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13500_ clknet_leaf_8_clk _00310_ net1074 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10712_ datapath.multiplication_module.multiplicand_i\[0\] _03321_ net573 vssd1 vssd1
+ vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[1\] sky130_fd_sc_hd__mux2_1
X_14480_ clknet_leaf_57_clk _01185_ net1160 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11692_ _04964_ _05885_ net148 net1452 vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08635__A _01935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13431_ clknet_leaf_126_clk _00241_ net1205 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10643_ _05441_ _05452_ _05461_ vssd1 vssd1 vccd1 vccd1 _05463_ sky130_fd_sc_hd__o21a_1
XANTENNA__08238__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09435__C1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08789__A1 _03296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08354__B net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12585__A2 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13362_ clknet_leaf_30_clk _00172_ net1125 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10574_ _03009_ net560 net464 _03149_ vssd1 vssd1 vccd1 vccd1 _05397_ sky130_fd_sc_hd__and4_1
XANTENNA_clkbuf_leaf_5_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12313_ net890 _04865_ net191 vssd1 vssd1 vccd1 vccd1 _06290_ sky130_fd_sc_hd__a21oi_1
X_13293_ clknet_leaf_125_clk _00103_ net1207 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_12244_ net2440 _06237_ net602 vssd1 vssd1 vccd1 vccd1 _06239_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09466__A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10348__A1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10899__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12175_ _06164_ _06172_ _06178_ vssd1 vssd1 vccd1 vccd1 _06196_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11000__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07764__A2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08961__A1 _03796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11126_ net235 net2629 net428 vssd1 vssd1 vccd1 vccd1 _00181_ sky130_fd_sc_hd__mux2_1
XFILLER_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10124__B _04057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11057_ net235 net2196 net432 vssd1 vssd1 vccd1 vccd1 _00117_ sky130_fd_sc_hd__mux2_1
XANTENNA__07516__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10008_ _04836_ _04841_ _04842_ vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__and3_1
XFILLER_36_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08248__C net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11959_ _05331_ _05782_ _05793_ _06004_ vssd1 vssd1 vccd1 vccd1 _06005_ sky130_fd_sc_hd__or4_1
XANTENNA__08477__B1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12766__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14678_ clknet_leaf_139_clk _01383_ net1099 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13629_ clknet_leaf_149_clk _00439_ net1060 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_17_Left_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07150_ _01984_ _01985_ vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__or2_1
XFILLER_146_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07081_ datapath.rf.registers\[9\]\[29\] net885 net877 datapath.rf.registers\[8\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01917_ sky130_fd_sc_hd__a22o_1
XANTENNA__12328__A2 _04084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09376__A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12514__B _05368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07608__B net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout128 _06369_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_26_Left_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout139 net142 vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__dlymetal6s2s_1
X_07983_ datapath.rf.registers\[31\]\[11\] net689 _02818_ net788 vssd1 vssd1 vccd1
+ vccd1 _02819_ sky130_fd_sc_hd__a211o_1
X_09722_ net630 _04557_ vssd1 vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__nor2_1
X_06934_ datapath.rf.registers\[28\]\[31\] net804 net801 datapath.rf.registers\[3\]\[31\]
+ _01767_ vssd1 vssd1 vccd1 vccd1 _01770_ sky130_fd_sc_hd__a221o_1
XFILLER_68_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09653_ net323 _03974_ vssd1 vssd1 vccd1 vccd1 _04489_ sky130_fd_sc_hd__nor2_1
X_06865_ _01684_ _01686_ _01700_ _01590_ vssd1 vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__o31a_2
XFILLER_28_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout272_A _05564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08180__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08604_ _02826_ _03438_ _02827_ _02727_ _02773_ vssd1 vssd1 vccd1 vccd1 _03440_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_2_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09584_ net354 _04419_ vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__or2_1
X_06796_ net1004 net1020 _01631_ net1028 datapath.ru.latched_instruction\[20\] vssd1
+ vssd1 vccd1 vccd1 _01632_ sky130_fd_sc_hd__a32o_1
XFILLER_70_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_118_Right_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08535_ datapath.rf.registers\[8\]\[0\] net878 _01768_ datapath.rf.registers\[28\]\[0\]
+ _03370_ vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__a221o_1
XANTENNA__08468__B1 _01772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14378__RESET_B net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_35_Left_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08466_ datapath.rf.registers\[27\]\[1\] net975 net939 vssd1 vssd1 vccd1 vccd1 _03302_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07997__C net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07417_ datapath.rf.registers\[26\]\[22\] net836 net826 datapath.rf.registers\[12\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout704_A net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08397_ datapath.rf.registers\[15\]\[2\] net988 net916 vssd1 vssd1 vccd1 vccd1 _03233_
+ sky130_fd_sc_hd__and3_1
XFILLER_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07348_ datapath.rf.registers\[28\]\[24\] net751 net731 datapath.rf.registers\[19\]\[24\]
+ _02173_ vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_21_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07279_ datapath.rf.registers\[9\]\[25\] net886 net828 datapath.rf.registers\[12\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1234_X net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09018_ net323 _03853_ vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__nor2_1
XANTENNA__07994__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10290_ datapath.PC\[7\] _05125_ net1254 vssd1 vssd1 vccd1 vccd1 _05126_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout694_X net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold160 net91 vssd1 vssd1 vccd1 vccd1 net1508 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 datapath.multiplication_module.multiplicand_i\[27\] vssd1 vssd1 vccd1 vccd1
+ net1519 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold182 datapath.multiplication_module.multiplicand_i\[30\] vssd1 vssd1 vccd1 vccd1
+ net1530 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08943__A1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold193 datapath.rf.registers\[7\]\[1\] vssd1 vssd1 vccd1 vccd1 net1541 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_120_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout861_X net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout640 net641 vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__buf_2
XANTENNA_fanout959_X net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout651 _01608_ vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__clkbuf_2
XFILLER_120_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout662 net663 vssd1 vssd1 vccd1 vccd1 net662 sky130_fd_sc_hd__buf_4
X_13980_ clknet_leaf_112_clk net1354 net1198 vssd1 vssd1 vccd1 vccd1 screen.counter.ack2
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout673 net674 vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__buf_4
XFILLER_120_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout684 net686 vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__clkbuf_4
Xfanout695 net697 vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12931_ net287 net1617 net397 vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__mux2_1
XANTENNA__08349__B net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12862_ _05695_ _05720_ vssd1 vssd1 vccd1 vccd1 _06553_ sky130_fd_sc_hd__nand2_1
XFILLER_37_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11813_ datapath.ru.latched_instruction\[19\] net334 net313 _01469_ vssd1 vssd1 vccd1
+ vccd1 _00679_ sky130_fd_sc_hd__a22o_1
X_14601_ clknet_leaf_20_clk _01306_ net1210 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12793_ net183 net1898 net495 vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__mux2_1
XFILLER_15_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09656__C1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11490__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14532_ clknet_leaf_23_clk _01237_ net1156 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11744_ net1480 net144 net139 _03170_ vssd1 vssd1 vccd1 vccd1 _00624_ sky130_fd_sc_hd__a22o_1
XFILLER_42_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07131__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14463_ clknet_leaf_10_clk _01168_ net1081 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_11675_ _05085_ _05885_ net150 net1434 vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__a2bb2o_1
X_13414_ clknet_leaf_17_clk _00224_ net1107 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10626_ _05445_ vssd1 vssd1 vccd1 vccd1 _05446_ sky130_fd_sc_hd__inv_2
XFILLER_139_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14394_ clknet_leaf_3_clk _01099_ net1078 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13345_ clknet_leaf_46_clk _00155_ net1148 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_77_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10557_ _05379_ _00003_ vssd1 vssd1 vccd1 vccd1 keypad.decode.d1 sky130_fd_sc_hd__and2_1
XFILLER_6_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07985__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07709__A _02522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13276_ clknet_leaf_10_clk _00086_ net1080 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10488_ screen.controlBus\[2\] screen.controlBus\[3\] _05317_ vssd1 vssd1 vccd1 vccd1
+ _05318_ sky130_fd_sc_hd__nor3_1
X_12227_ screen.counter.currentCt\[13\] _06227_ vssd1 vssd1 vccd1 vccd1 _06228_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_90_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07198__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07737__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08934__A1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12158_ net1276 _06184_ _06185_ vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_9_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11109_ net287 net1720 net429 vssd1 vssd1 vccd1 vccd1 _00164_ sky130_fd_sc_hd__mux2_1
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12089_ _06121_ _06122_ _06123_ _06127_ vssd1 vssd1 vccd1 vccd1 _06128_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_108_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08162__A2 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06650_ datapath.ru.latched_instruction\[24\] _01464_ _01479_ datapath.ru.latched_instruction\[27\]
+ vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_88_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07731__X _02567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06581_ net1280 vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__inv_2
XANTENNA__12496__S net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08320_ _03154_ _03155_ vssd1 vssd1 vccd1 vccd1 _03156_ sky130_fd_sc_hd__or2_1
XFILLER_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08251_ datapath.rf.registers\[24\]\[5\] net857 net813 datapath.rf.registers\[23\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03087_ sky130_fd_sc_hd__a22o_1
XANTENNA__07610__C net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07202_ datapath.rf.registers\[30\]\[27\] net759 net676 datapath.rf.registers\[29\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02038_ sky130_fd_sc_hd__a22o_1
XANTENNA__12549__A2 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08182_ datapath.rf.registers\[22\]\[7\] net736 net677 datapath.rf.registers\[29\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03018_ sky130_fd_sc_hd__a22o_1
Xteam_04_1304 vssd1 vssd1 vccd1 vccd1 team_04_1304/HI gpio_oeb[13] sky130_fd_sc_hd__conb_1
X_07133_ datapath.rf.registers\[31\]\[28\] net795 net792 datapath.rf.registers\[18\]\[28\]
+ _01968_ vssd1 vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__a221o_1
Xteam_04_1315 vssd1 vssd1 vccd1 vccd1 team_04_1315/HI gpio_out[8] sky130_fd_sc_hd__conb_1
XFILLER_146_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xteam_04_1326 vssd1 vssd1 vccd1 vccd1 team_04_1326/HI gpio_out[30] sky130_fd_sc_hd__conb_1
Xteam_04_1337 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] team_04_1337/LO sky130_fd_sc_hd__conb_1
XANTENNA__13120__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_04_1348 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] team_04_1348/LO sky130_fd_sc_hd__conb_1
XFILLER_145_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07976__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07064_ datapath.rf.registers\[14\]\[30\] net776 net756 datapath.rf.registers\[12\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07728__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout487_A _06552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07966_ _02790_ _02791_ _02801_ vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__or3b_1
XANTENNA__12260__A net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09705_ net357 _04359_ vssd1 vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__or2_1
XANTENNA__06896__C _01656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06917_ net954 net932 vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__and2_4
XTAP_TAPCELL_ROW_52_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07897_ datapath.rf.registers\[16\]\[12\] net863 _01765_ datapath.rf.registers\[13\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02733_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout654_A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_94_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_94_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_83_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09636_ _03428_ _03561_ vssd1 vssd1 vccd1 vccd1 _04472_ sky130_fd_sc_hd__xor2_1
X_06848_ datapath.ru.latched_instruction\[19\] net988 _01664_ datapath.ru.latched_instruction\[8\]
+ _01683_ vssd1 vssd1 vccd1 vccd1 _01684_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07900__A2 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_43_Left_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09567_ net324 _04080_ _04402_ net642 vssd1 vssd1 vccd1 vccd1 _04403_ sky130_fd_sc_hd__o211a_1
X_06779_ net1005 net1021 _01615_ vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__and3_1
XANTENNA__10919__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout821_A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08456__Y _03292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11604__A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08518_ datapath.rf.registers\[2\]\[1\] net914 net909 vssd1 vssd1 vccd1 vccd1 _03354_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_26_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09498_ _03642_ _04314_ _04328_ _03614_ vssd1 vssd1 vccd1 vccd1 _04334_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_156_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08449_ datapath.rf.registers\[7\]\[2\] net674 net662 datapath.rf.registers\[5\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03285_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_156_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout707_X net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11460_ net1840 net244 net406 vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__mux2_1
XFILLER_23_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10411_ net906 _03548_ net626 _03546_ _05246_ vssd1 vssd1 vccd1 vccd1 _05247_ sky130_fd_sc_hd__a221o_1
X_11391_ net2138 net252 net411 vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13030__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13130_ net1670 net286 net385 vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__mux2_1
X_10342_ _04538_ _04562_ vssd1 vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__nor2_1
XFILLER_152_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08351__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13061_ _05696_ _06558_ vssd1 vssd1 vccd1 vccd1 _06560_ sky130_fd_sc_hd__nor2_1
X_10273_ net1267 net466 net1042 _05108_ vssd1 vssd1 vccd1 vccd1 _05109_ sky130_fd_sc_hd__o211a_1
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12012_ _06021_ _06025_ _06050_ _06055_ vssd1 vssd1 vccd1 vccd1 _06056_ sky130_fd_sc_hd__or4_1
XANTENNA__07719__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10723__A1 _02912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11485__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout470 net473 vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__buf_6
Xfanout481 _06556_ vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__clkbuf_4
XFILLER_120_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout492 _06551_ vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__clkbuf_8
X_13963_ clknet_leaf_104_clk _00741_ net1224 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_85_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_clk sky130_fd_sc_hd__clkbuf_8
X_12914_ net2102 net219 net482 vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__mux2_1
X_13894_ clknet_leaf_43_clk keypad.decode.d1 net1150 vssd1 vssd1 vccd1 vccd1 keypad.decode.d2
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12845_ net250 net1967 net487 vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07711__B net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12776_ net263 net2277 net496 vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__mux2_1
XANTENNA__07104__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08301__C1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08447__A3 _01831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08526__C net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11727_ net14 net1033 net1023 net2199 vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__o22a_1
XFILLER_148_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08852__A0 _02312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14515_ clknet_leaf_35_clk _01220_ net1130 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11658_ net2646 _05875_ _05878_ vssd1 vssd1 vccd1 vccd1 _00551_ sky130_fd_sc_hd__a21o_1
XANTENNA__09919__A _01585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14446_ clknet_leaf_1_clk _01151_ net1056 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_156_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13864__RESET_B net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10609_ net38 _05379_ _05380_ net37 vssd1 vssd1 vccd1 vccd1 _05429_ sky130_fd_sc_hd__and4b_1
X_14377_ clknet_leaf_91_clk _01082_ net1233 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_127_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11589_ _05760_ _05812_ vssd1 vssd1 vccd1 vccd1 _05813_ sky130_fd_sc_hd__nor2_1
Xhold907 datapath.rf.registers\[29\]\[18\] vssd1 vssd1 vccd1 vccd1 net2255 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07958__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10411__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13328_ clknet_leaf_24_clk _00138_ net1158 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold918 datapath.rf.registers\[8\]\[25\] vssd1 vssd1 vccd1 vccd1 net2266 sky130_fd_sc_hd__dlygate4sd3_1
Xhold929 datapath.rf.registers\[23\]\[12\] vssd1 vssd1 vccd1 vccd1 net2277 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10962__A1 _01500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap659 _05364_ vssd1 vssd1 vccd1 vccd1 net659 sky130_fd_sc_hd__clkbuf_4
XFILLER_143_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13259_ clknet_leaf_55_clk _00069_ net1179 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09654__A net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10714__A1 _03204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11395__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07820_ datapath.rf.registers\[24\]\[14\] net857 net827 datapath.rf.registers\[12\]\[14\]
+ _02655_ vssd1 vssd1 vccd1 vccd1 _02656_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_4_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08383__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07591__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07751_ _02576_ _02582_ _02586_ net782 datapath.rf.registers\[0\]\[16\] vssd1 vssd1
+ vccd1 vccd1 _02587_ sky130_fd_sc_hd__o32a_4
XANTENNA_clkbuf_leaf_92_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_76_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_93_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06702_ datapath.ru.latched_instruction\[20\] datapath.ru.latched_instruction\[21\]
+ datapath.ru.latched_instruction\[22\] datapath.ru.latched_instruction\[23\] vssd1
+ vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__or4_1
XANTENNA__08135__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07682_ _02514_ _02515_ _02516_ _02517_ vssd1 vssd1 vccd1 vccd1 _02518_ sky130_fd_sc_hd__or4_1
XANTENNA__07343__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09421_ _02661_ _02705_ net442 vssd1 vssd1 vccd1 vccd1 _04257_ sky130_fd_sc_hd__mux2_1
X_06633_ datapath.ru.latched_instruction\[30\] _01466_ _01468_ _01471_ _01465_ vssd1
+ vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__o2111a_1
XFILLER_80_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13115__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08717__B _03228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09352_ _04185_ _04186_ net454 vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__a21o_1
X_06564_ datapath.ru.n_memwrite vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_23_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08303_ datapath.rf.registers\[16\]\[4\] net860 net826 datapath.rf.registers\[12\]\[4\]
+ _03138_ vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__a221o_1
XFILLER_139_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_150_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08843__A0 _03419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08436__C _01823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09283_ _02544_ _02545_ vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__and2b_2
XANTENNA__12954__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout235_A _05616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08234_ datapath.rf.registers\[19\]\[6\] net730 net726 datapath.rf.registers\[25\]\[6\]
+ _03069_ vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_30_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09399__B2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08165_ datapath.rf.registers\[4\]\[7\] net865 _02995_ _02996_ _03000_ vssd1 vssd1
+ vccd1 vccd1 _03001_ sky130_fd_sc_hd__a2111oi_1
XANTENNA_fanout402_A _06549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1144_A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07116_ datapath.rf.registers\[3\]\[29\] net770 net669 datapath.rf.registers\[21\]\[29\]
+ _01951_ vssd1 vssd1 vccd1 vccd1 _01952_ sky130_fd_sc_hd__a221o_1
X_08096_ _02919_ _02925_ _02931_ vssd1 vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__nor3_1
XFILLER_146_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08171__C net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload80 clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 clkload80/Y sky130_fd_sc_hd__bufinv_16
XANTENNA_clkbuf_leaf_45_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07047_ datapath.rf.registers\[16\]\[30\] net862 net858 datapath.rf.registers\[24\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__a22o_1
Xclkload91 clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 clkload91/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09564__A net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10705__A1 _02876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout771_A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout392_X net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout869_A net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08374__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08998_ _01888_ _01934_ net442 vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_149_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07582__B1 _02417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07949_ datapath.rf.registers\[6\]\[11\] net952 net934 vssd1 vssd1 vccd1 vccd1 _02785_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout657_X net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_67_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08126__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_103_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10960_ datapath.PC\[0\] _05237_ net897 vssd1 vssd1 vccd1 vccd1 _05698_ sky130_fd_sc_hd__mux2_1
XFILLER_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09619_ _04454_ vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__inv_2
X_10891_ _05636_ _05637_ vssd1 vssd1 vccd1 vccd1 _05638_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout824_X net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13025__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12630_ datapath.mulitply_result\[20\] datapath.multiplication_module.multiplicand_i\[20\]
+ vssd1 vssd1 vccd1 vccd1 _06472_ sky130_fd_sc_hd__or2_1
XFILLER_71_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_118_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08346__C net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12561_ net500 _06413_ _06414_ net504 net2081 vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__a32o_1
XANTENNA__12864__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11512_ _05361_ _05353_ _05736_ vssd1 vssd1 vccd1 vccd1 _05737_ sky130_fd_sc_hd__mux2_1
X_14300_ clknet_leaf_94_clk _01005_ net1217 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[20\]
+ sky130_fd_sc_hd__dfrtp_2
X_12492_ net251 net2573 net506 vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__mux2_1
XFILLER_156_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14231_ clknet_leaf_42_clk _00952_ net1144 vssd1 vssd1 vccd1 vccd1 columns.count\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11443_ _05696_ _05732_ vssd1 vssd1 vccd1 vccd1 _05733_ sky130_fd_sc_hd__nor2_4
XANTENNA__06860__A2 _01610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10237__X _05073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire189 _05203_ vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__buf_1
X_14162_ clknet_leaf_65_clk _00917_ net1235 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11374_ net170 net1573 net518 vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__mux2_1
XANTENNA__10944__A1 _01466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13113_ net220 net1872 net470 vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__mux2_1
X_10325_ net1040 _05158_ _05160_ net635 vssd1 vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__a211o_1
XFILLER_125_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14093_ clknet_leaf_110_clk _00859_ net1201 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_113_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13044_ net247 net2535 net474 vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__mux2_1
X_10256_ _04835_ _04851_ _04854_ vssd1 vssd1 vccd1 vccd1 _05092_ sky130_fd_sc_hd__o21a_1
XFILLER_3_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09905__C _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1210 net1213 vssd1 vssd1 vccd1 vccd1 net1210 sky130_fd_sc_hd__clkbuf_4
Xfanout1221 net1222 vssd1 vssd1 vccd1 vccd1 net1221 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08365__A2 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1232 net1251 vssd1 vssd1 vccd1 vccd1 net1232 sky130_fd_sc_hd__clkbuf_4
X_10187_ _04146_ _05022_ vssd1 vssd1 vccd1 vccd1 _05023_ sky130_fd_sc_hd__nand2_1
XANTENNA__10413__A net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1243 net1244 vssd1 vssd1 vccd1 vccd1 net1243 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10172__A2 net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1254 net1257 vssd1 vssd1 vccd1 vccd1 net1254 sky130_fd_sc_hd__clkbuf_4
XFILLER_94_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1265 datapath.PC\[22\] vssd1 vssd1 vccd1 vccd1 net1265 sky130_fd_sc_hd__buf_2
Xfanout1276 screen.counter.ct\[9\] vssd1 vssd1 vccd1 vccd1 net1276 sky130_fd_sc_hd__buf_2
XFILLER_66_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1287 net1289 vssd1 vssd1 vccd1 vccd1 net1287 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_58_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08117__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_11_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_11_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_93_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09921__B _01786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13946_ clknet_leaf_111_clk _00724_ net1202 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07325__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_85_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13877_ clknet_leaf_53_clk _00681_ net1183 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[21\]
+ sky130_fd_sc_hd__dfrtp_4
X_12828_ net1860 net169 net491 vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__mux2_1
XFILLER_62_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12774__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12759_ net2092 net178 net404 vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__mux2_1
XFILLER_30_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14429_ clknet_leaf_147_clk _01134_ net1088 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_144_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold704 datapath.rf.registers\[29\]\[8\] vssd1 vssd1 vccd1 vccd1 net2052 sky130_fd_sc_hd__dlygate4sd3_1
Xhold715 datapath.rf.registers\[2\]\[16\] vssd1 vssd1 vccd1 vccd1 net2063 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold726 datapath.rf.registers\[18\]\[17\] vssd1 vssd1 vccd1 vccd1 net2074 sky130_fd_sc_hd__dlygate4sd3_1
Xhold737 datapath.rf.registers\[29\]\[7\] vssd1 vssd1 vccd1 vccd1 net2085 sky130_fd_sc_hd__dlygate4sd3_1
X_09970_ _04746_ _04748_ _04804_ _04745_ vssd1 vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__a31o_1
Xhold748 datapath.rf.registers\[23\]\[1\] vssd1 vssd1 vccd1 vccd1 net2096 sky130_fd_sc_hd__dlygate4sd3_1
Xhold759 datapath.rf.registers\[5\]\[28\] vssd1 vssd1 vccd1 vccd1 net2107 sky130_fd_sc_hd__dlygate4sd3_1
X_08921_ _03489_ _03594_ _03487_ vssd1 vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__a21oi_1
XFILLER_112_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08356__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08852_ _02312_ _02365_ net444 vssd1 vssd1 vccd1 vccd1 _03688_ sky130_fd_sc_hd__mux2_1
XFILLER_97_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07803_ datapath.rf.registers\[23\]\[14\] net940 net923 vssd1 vssd1 vccd1 vccd1 _02639_
+ sky130_fd_sc_hd__and3_1
XFILLER_85_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08783_ net971 _03172_ _03615_ vssd1 vssd1 vccd1 vccd1 _03619_ sky130_fd_sc_hd__mux2_2
XANTENNA__12949__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_49_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_66_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08108__A2 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07734_ datapath.rf.registers\[26\]\[16\] net778 net675 datapath.rf.registers\[29\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__a22o_1
XANTENNA__08287__X _03123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07665_ datapath.rf.registers\[23\]\[17\] net941 net925 vssd1 vssd1 vccd1 vccd1 _02501_
+ sky130_fd_sc_hd__and3_1
XFILLER_53_644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09404_ _02727_ _03441_ vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__and2b_1
X_06616_ datapath.ru.latched_instruction\[17\] _01452_ _01454_ datapath.ru.latched_instruction\[18\]
+ vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__o22ai_1
XPHY_EDGE_ROW_9_Left_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07596_ datapath.rf.registers\[24\]\[19\] net768 net712 datapath.rf.registers\[11\]\[19\]
+ _02431_ vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__a221o_1
XANTENNA__14054__CLK clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13786__RESET_B net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08816__A0 _01666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09335_ net906 _03518_ vssd1 vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout1261_A net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07095__A2 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09266_ _04100_ _04101_ net454 vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__a21o_1
X_08217_ datapath.rf.registers\[25\]\[6\] net841 net804 datapath.rf.registers\[28\]\[6\]
+ _03052_ vssd1 vssd1 vccd1 vccd1 _03053_ sky130_fd_sc_hd__a221o_1
XANTENNA__08029__D1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09197_ _03876_ _04031_ net374 vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__mux2_1
XFILLER_153_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout405_X net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08148_ _02960_ _02983_ vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__and2_1
XANTENNA__10387__C1 _03614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout986_A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08079_ datapath.rf.registers\[24\]\[9\] net768 net689 datapath.rf.registers\[31\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02915_ sky130_fd_sc_hd__a22o_1
XFILLER_150_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10110_ datapath.PC\[19\] _03743_ vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__nand2_1
XFILLER_1_924 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09294__A _02466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11090_ net239 net1992 net536 vssd1 vssd1 vccd1 vccd1 _00147_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout774_X net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10041_ _04874_ _04876_ vssd1 vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__nand2_1
Xhold20 keypad.decode.d2 vssd1 vssd1 vccd1 vccd1 net1368 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold31 screen.counter.currentCt\[22\] vssd1 vssd1 vccd1 vccd1 net1379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 screen.controlBus\[29\] vssd1 vssd1 vccd1 vccd1 net1390 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold53 screen.controlBus\[13\] vssd1 vssd1 vccd1 vccd1 net1401 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12859__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold64 screen.controlBus\[27\] vssd1 vssd1 vccd1 vccd1 net1412 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout941_X net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold75 net60 vssd1 vssd1 vccd1 vccd1 net1423 sky130_fd_sc_hd__dlygate4sd3_1
X_13800_ clknet_leaf_73_clk _00609_ net1184 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[21\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold86 net66 vssd1 vssd1 vccd1 vccd1 net1434 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold97 net104 vssd1 vssd1 vccd1 vccd1 net1445 sky130_fd_sc_hd__dlygate4sd3_1
X_11992_ _06023_ _06026_ _06036_ vssd1 vssd1 vccd1 vccd1 _06037_ sky130_fd_sc_hd__or3_1
XFILLER_72_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13731_ clknet_leaf_119_clk _00541_ net1191 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10943_ _01429_ net615 _05682_ net654 vssd1 vssd1 vccd1 vccd1 _05683_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_67_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07261__B net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13662_ clknet_leaf_147_clk _00472_ net1064 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10874_ net231 net2016 net542 vssd1 vssd1 vccd1 vccd1 _00022_ sky130_fd_sc_hd__mux2_1
XFILLER_45_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12613_ datapath.mulitply_result\[17\] datapath.multiplication_module.multiplicand_i\[17\]
+ vssd1 vssd1 vccd1 vccd1 _06458_ sky130_fd_sc_hd__nor2_1
X_13593_ clknet_leaf_32_clk _00403_ net1122 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09469__A _02856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12544_ datapath.mulitply_result\[6\] datapath.multiplication_module.multiplicand_i\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06400_ sky130_fd_sc_hd__nand2_1
XANTENNA__07086__A2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12475_ net164 _05998_ net126 screen.register.currentXbus\[31\] vssd1 vssd1 vccd1
+ vccd1 _00877_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_138_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12367__B1 _05002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14214_ clknet_leaf_48_clk datapath.multiplication_module.multiplicand_i_n\[25\]
+ net1175 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11426_ net245 net1867 net514 vssd1 vssd1 vccd1 vccd1 _00466_ sky130_fd_sc_hd__mux2_1
XANTENNA_6 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09232__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14145_ clknet_leaf_138_clk _00902_ net1098 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_11357_ net253 net2462 net518 vssd1 vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__mux2_1
XFILLER_152_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07794__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10308_ _04857_ _05143_ vssd1 vssd1 vccd1 vccd1 _05144_ sky130_fd_sc_hd__or2_1
XFILLER_3_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14076_ clknet_leaf_121_clk _00843_ net1199 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11288_ net252 net2330 net522 vssd1 vssd1 vccd1 vccd1 _00336_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13027_ _05514_ _05690_ vssd1 vssd1 vccd1 vccd1 _06558_ sky130_fd_sc_hd__or2_1
X_10239_ _04839_ _04840_ vssd1 vssd1 vccd1 vccd1 _05075_ sky130_fd_sc_hd__and2b_1
Xfanout1040 net1042 vssd1 vssd1 vccd1 vccd1 net1040 sky130_fd_sc_hd__clkbuf_4
XFILLER_67_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1051 _01437_ vssd1 vssd1 vccd1 vccd1 net1051 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07010__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1062 net1066 vssd1 vssd1 vccd1 vccd1 net1062 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12769__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1073 net1074 vssd1 vssd1 vccd1 vccd1 net1073 sky130_fd_sc_hd__clkbuf_4
Xfanout1084 net1121 vssd1 vssd1 vccd1 vccd1 net1084 sky130_fd_sc_hd__buf_2
Xfanout1095 net1096 vssd1 vssd1 vccd1 vccd1 net1095 sky130_fd_sc_hd__clkbuf_4
XFILLER_75_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13929_ clknet_leaf_110_clk _00707_ net1201 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_81_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10289__S net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10302__C1 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08510__A2 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07171__B net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07450_ net563 _02284_ vssd1 vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__nand2_1
X_07381_ _02207_ _02216_ datapath.rf.registers\[0\]\[23\] net866 vssd1 vssd1 vccd1
+ vccd1 _02217_ sky130_fd_sc_hd__o2bb2a_4
X_09120_ _03875_ _03955_ net367 vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09471__A0 _02961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12070__A2 _05773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09051_ net456 _03843_ _03844_ _03886_ vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__a31oi_1
XFILLER_30_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08002_ datapath.rf.registers\[22\]\[10\] net952 net925 vssd1 vssd1 vccd1 vccd1 _02838_
+ sky130_fd_sc_hd__and3_1
Xhold501 datapath.rf.registers\[21\]\[25\] vssd1 vssd1 vccd1 vccd1 net1849 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10908__A1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold512 datapath.rf.registers\[1\]\[31\] vssd1 vssd1 vccd1 vccd1 net1860 sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 datapath.rf.registers\[24\]\[13\] vssd1 vssd1 vccd1 vccd1 net1871 sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 datapath.rf.registers\[31\]\[18\] vssd1 vssd1 vccd1 vccd1 net1882 sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 datapath.rf.registers\[20\]\[7\] vssd1 vssd1 vccd1 vccd1 net1893 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold556 datapath.rf.registers\[30\]\[11\] vssd1 vssd1 vccd1 vccd1 net1904 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07785__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold567 datapath.multiplication_module.multiplicand_i\[6\] vssd1 vssd1 vccd1 vccd1
+ net1915 sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 datapath.rf.registers\[31\]\[9\] vssd1 vssd1 vccd1 vccd1 net1926 sky130_fd_sc_hd__dlygate4sd3_1
Xhold589 datapath.rf.registers\[1\]\[25\] vssd1 vssd1 vccd1 vccd1 net1937 sky130_fd_sc_hd__dlygate4sd3_1
X_09953_ datapath.PC\[4\] _03150_ vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__or2_1
XFILLER_106_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08329__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08904_ datapath.PC\[14\] _03739_ vssd1 vssd1 vccd1 vccd1 _03740_ sky130_fd_sc_hd__or2_1
X_09884_ net1263 net594 vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__nand2_1
XFILLER_58_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07537__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1107_A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07914__X _02750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1201 datapath.rf.registers\[2\]\[8\] vssd1 vssd1 vccd1 vccd1 net2549 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_4_0_clk_X clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07001__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1212 screen.counter.currentCt\[6\] vssd1 vssd1 vccd1 vccd1 net2560 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09842__A net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1223 datapath.rf.registers\[14\]\[29\] vssd1 vssd1 vccd1 vccd1 net2571 sky130_fd_sc_hd__dlygate4sd3_1
X_08835_ _01609_ net606 _03669_ vssd1 vssd1 vccd1 vccd1 _03671_ sky130_fd_sc_hd__or3_4
Xhold1234 datapath.rf.registers\[24\]\[7\] vssd1 vssd1 vccd1 vccd1 net2582 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1245 screen.counter.currentCt\[9\] vssd1 vssd1 vccd1 vccd1 net2593 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1256 screen.counter.ct\[22\] vssd1 vssd1 vccd1 vccd1 net2604 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1267 datapath.mulitply_result\[19\] vssd1 vssd1 vccd1 vccd1 net2615 sky130_fd_sc_hd__dlygate4sd3_1
X_08766_ net642 _03601_ vssd1 vssd1 vccd1 vccd1 _03602_ sky130_fd_sc_hd__or2_1
Xhold1278 mmio.memload_or_instruction\[24\] vssd1 vssd1 vccd1 vccd1 net2626 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1289 datapath.rf.registers\[24\]\[12\] vssd1 vssd1 vccd1 vccd1 net2637 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08458__A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07717_ datapath.rf.registers\[10\]\[16\] net879 net853 datapath.rf.registers\[19\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02553_ sky130_fd_sc_hd__a22o_1
X_08697_ _03532_ vssd1 vssd1 vccd1 vccd1 _03533_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_49_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout734_A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07648_ datapath.rf.registers\[25\]\[18\] net726 net714 datapath.rf.registers\[4\]\[18\]
+ _02483_ vssd1 vssd1 vccd1 vccd1 _02484_ sky130_fd_sc_hd__a221o_1
XFILLER_25_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout901_A net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout522_X net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07579_ datapath.rf.registers\[8\]\[19\] net878 _02388_ _02389_ _02401_ vssd1 vssd1
+ vccd1 vccd1 _02415_ sky130_fd_sc_hd__a2111oi_1
XTAP_TAPCELL_ROW_62_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09318_ net369 _04152_ _04153_ vssd1 vssd1 vccd1 vccd1 _04154_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_62_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07068__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10590_ _05411_ _05412_ vssd1 vssd1 vccd1 vccd1 _05413_ sky130_fd_sc_hd__or2_1
XFILLER_40_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09462__B1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08193__A _01598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10072__A1 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09249_ _02441_ _02442_ vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__nand2_2
X_12260_ net636 _04338_ vssd1 vssd1 vccd1 vccd1 _06250_ sky130_fd_sc_hd__nand2_1
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout891_X net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08984__A1_N net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11211_ net302 net1954 net528 vssd1 vssd1 vccd1 vccd1 _00261_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout989_X net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12191_ _06167_ screen.counter.currentCt\[0\] vssd1 vssd1 vccd1 vccd1 _06205_ sky130_fd_sc_hd__and2b_1
XFILLER_134_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12443__A net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10375__A2 net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput43 net43 vssd1 vssd1 vccd1 vccd1 ADR_O[12] sky130_fd_sc_hd__buf_2
X_11142_ net261 net2631 net532 vssd1 vssd1 vccd1 vccd1 _00195_ sky130_fd_sc_hd__mux2_1
XFILLER_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput54 net54 vssd1 vssd1 vccd1 vccd1 ADR_O[22] sky130_fd_sc_hd__buf_2
XFILLER_150_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 ADR_O[3] sky130_fd_sc_hd__buf_2
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 DAT_O[12] sky130_fd_sc_hd__buf_2
XANTENNA__09517__A1 _02856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput87 net87 vssd1 vssd1 vccd1 vccd1 DAT_O[22] sky130_fd_sc_hd__buf_2
XFILLER_1_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11073_ net208 net1955 net536 vssd1 vssd1 vccd1 vccd1 _00130_ sky130_fd_sc_hd__mux2_1
XANTENNA__07256__B _02091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput98 net98 vssd1 vssd1 vccd1 vccd1 DAT_O[3] sky130_fd_sc_hd__buf_2
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07528__B1 _02363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input30_A DAT_I[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10024_ _04856_ _04859_ _04855_ vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__and3b_1
XANTENNA__07824__X _02660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11493__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11975_ _05758_ _05852_ vssd1 vssd1 vccd1 vccd1 _06020_ sky130_fd_sc_hd__nor2_1
XANTENNA__10835__A0 _04207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13714_ clknet_leaf_32_clk _00524_ net1123 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10926_ _03827_ _05667_ net901 vssd1 vssd1 vccd1 vccd1 _05668_ sky130_fd_sc_hd__mux2_2
X_14694_ clknet_leaf_11_clk _01399_ net1083 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07700__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10857_ datapath.mulitply_result\[18\] net597 _05608_ net617 vssd1 vssd1 vccd1 vccd1
+ _05609_ sky130_fd_sc_hd__a211o_1
X_13645_ clknet_leaf_124_clk _00455_ net1207 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09453__A0 _02751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07059__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13576_ clknet_leaf_61_clk _00386_ net1165 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10788_ _05548_ _05549_ vssd1 vssd1 vccd1 vccd1 _05550_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_30_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12527_ datapath.mulitply_result\[3\] datapath.multiplication_module.multiplicand_i\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06386_ sky130_fd_sc_hd__nor2_1
XANTENNA__10138__A net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12458_ net165 _05964_ net127 screen.register.currentXbus\[14\] vssd1 vssd1 vccd1
+ vccd1 _00860_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08831__A _03636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06903__X _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09756__A1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11409_ _05517_ _05710_ vssd1 vssd1 vccd1 vccd1 _05731_ sky130_fd_sc_hd__nand2_4
X_12389_ _05946_ net159 vssd1 vssd1 vccd1 vccd1 _06342_ sky130_fd_sc_hd__nor2_1
XFILLER_114_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08550__B net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07767__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06989__C _01647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07231__A2 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14128_ clknet_leaf_27_clk _00885_ net1134 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_06950_ net610 net596 vssd1 vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__and2_2
XFILLER_140_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14059_ clknet_leaf_121_clk _00826_ net1199 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07519__B1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12499__S net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06881_ _01656_ net962 vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__and2_2
XANTENNA__08192__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08620_ _02365_ _02386_ vssd1 vssd1 vccd1 vccd1 _03456_ sky130_fd_sc_hd__nand2_1
XFILLER_95_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06742__A1 _01500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08551_ datapath.rf.registers\[17\]\[0\] _01800_ net907 vssd1 vssd1 vccd1 vccd1 _03387_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_38_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_124_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07502_ datapath.rf.registers\[2\]\[20\] net982 net949 vssd1 vssd1 vccd1 vccd1 _02338_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_141_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08482_ _03315_ _03316_ _03317_ vssd1 vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__or3_1
XANTENNA__07298__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07433_ datapath.rf.registers\[26\]\[22\] net778 net722 datapath.rf.registers\[18\]\[22\]
+ _02267_ vssd1 vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout148_A net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13123__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12579__B1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07364_ datapath.rf.registers\[29\]\[23\] net974 net917 vssd1 vssd1 vccd1 vccd1 _02200_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_44_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_99_Left_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09103_ net338 _03936_ _03938_ _03673_ vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__o211a_1
XANTENNA__12962__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07295_ datapath.rf.registers\[16\]\[25\] net740 net712 datapath.rf.registers\[11\]\[25\]
+ _02130_ vssd1 vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1057_A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09034_ _03590_ _03866_ net578 vssd1 vssd1 vccd1 vccd1 _03870_ sky130_fd_sc_hd__o21a_1
Xhold320 datapath.rf.registers\[14\]\[2\] vssd1 vssd1 vccd1 vccd1 net1668 sky130_fd_sc_hd__dlygate4sd3_1
Xhold331 datapath.rf.registers\[7\]\[5\] vssd1 vssd1 vccd1 vccd1 net1679 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12263__A net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1224_A net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold342 datapath.rf.registers\[9\]\[17\] vssd1 vssd1 vccd1 vccd1 net1690 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08460__B _03294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold353 datapath.rf.registers\[24\]\[2\] vssd1 vssd1 vccd1 vccd1 net1701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 datapath.rf.registers\[7\]\[13\] vssd1 vssd1 vccd1 vccd1 net1712 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06899__C net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold375 datapath.rf.registers\[6\]\[7\] vssd1 vssd1 vccd1 vccd1 net1723 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout684_A net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout800 _01772_ vssd1 vssd1 vccd1 vccd1 net800 sky130_fd_sc_hd__clkbuf_8
Xhold386 datapath.rf.registers\[27\]\[2\] vssd1 vssd1 vccd1 vccd1 net1734 sky130_fd_sc_hd__dlygate4sd3_1
Xhold397 datapath.rf.registers\[12\]\[26\] vssd1 vssd1 vccd1 vccd1 net1745 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout811 net812 vssd1 vssd1 vccd1 vccd1 net811 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout822 net823 vssd1 vssd1 vccd1 vccd1 net822 sky130_fd_sc_hd__clkbuf_4
X_09936_ datapath.PC\[5\] _03124_ vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__nand2_1
Xfanout833 net835 vssd1 vssd1 vccd1 vccd1 net833 sky130_fd_sc_hd__clkbuf_4
Xfanout844 _01738_ vssd1 vssd1 vccd1 vccd1 net844 sky130_fd_sc_hd__buf_4
Xfanout855 _01733_ vssd1 vssd1 vccd1 vccd1 net855 sky130_fd_sc_hd__clkbuf_8
Xfanout866 net867 vssd1 vssd1 vccd1 vccd1 net866 sky130_fd_sc_hd__buf_6
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout877 net878 vssd1 vssd1 vccd1 vccd1 net877 sky130_fd_sc_hd__buf_4
X_09867_ _03032_ _04701_ _04702_ _04675_ vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout851_A _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout472_X net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout888 net889 vssd1 vssd1 vccd1 vccd1 net888 sky130_fd_sc_hd__clkbuf_2
Xhold1020 datapath.rf.registers\[30\]\[4\] vssd1 vssd1 vccd1 vccd1 net2368 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout899 net903 vssd1 vssd1 vccd1 vccd1 net899 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08183__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout949_A net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1031 datapath.mulitply_result\[13\] vssd1 vssd1 vccd1 vccd1 net2379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1042 datapath.rf.registers\[11\]\[16\] vssd1 vssd1 vccd1 vccd1 net2390 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07804__B net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1053 datapath.rf.registers\[30\]\[16\] vssd1 vssd1 vccd1 vccd1 net2401 sky130_fd_sc_hd__dlygate4sd3_1
X_08818_ net612 _03417_ _03644_ _03384_ vssd1 vssd1 vccd1 vccd1 _03654_ sky130_fd_sc_hd__a211o_1
X_09798_ net311 _04632_ _04633_ _03641_ vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__o22a_1
Xhold1064 datapath.rf.registers\[7\]\[11\] vssd1 vssd1 vccd1 vccd1 net2412 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1075 datapath.rf.registers\[19\]\[31\] vssd1 vssd1 vccd1 vccd1 net2423 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1086 datapath.rf.registers\[22\]\[3\] vssd1 vssd1 vccd1 vccd1 net2434 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1097 datapath.rf.registers\[13\]\[30\] vssd1 vssd1 vccd1 vccd1 net2445 sky130_fd_sc_hd__dlygate4sd3_1
X_08749_ _03507_ _03508_ _03582_ _03505_ _03503_ vssd1 vssd1 vccd1 vccd1 _03585_ sky130_fd_sc_hd__a311o_1
XANTENNA_fanout737_X net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11760_ net1491 net143 net138 _02385_ vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__a22o_1
XANTENNA__12282__A2 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10711_ net558 _05368_ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[0\]
+ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11691_ _04997_ net153 net148 net1439 vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout904_X net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13033__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10642_ _05428_ _05450_ vssd1 vssd1 vccd1 vccd1 _05462_ sky130_fd_sc_hd__nor2_1
X_13430_ clknet_leaf_141_clk _00240_ net1096 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08354__C net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08789__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13361_ clknet_leaf_39_clk _00171_ net1141 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12872__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10573_ _05394_ _05395_ vssd1 vssd1 vccd1 vccd1 _05396_ sky130_fd_sc_hd__or2_1
XFILLER_6_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09747__A _04239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12312_ datapath.PC\[15\] net308 _06289_ vssd1 vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__a21o_1
XANTENNA__07461__A2 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13292_ clknet_leaf_15_clk _00102_ net1103 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_108_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11488__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12243_ screen.counter.currentCt\[19\] _06237_ vssd1 vssd1 vccd1 vccd1 _06238_ sky130_fd_sc_hd__and2_1
XANTENNA__07749__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12174_ net1271 net1272 _06192_ screen.counter.ct\[16\] vssd1 vssd1 vccd1 vccd1 _06195_
+ sky130_fd_sc_hd__a31o_1
XFILLER_150_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11125_ net220 net1756 net426 vssd1 vssd1 vccd1 vccd1 _00180_ sky130_fd_sc_hd__mux2_1
XFILLER_95_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11056_ net220 net2095 net430 vssd1 vssd1 vccd1 vccd1 _00116_ sky130_fd_sc_hd__mux2_1
XFILLER_95_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08369__Y _03205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08174__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10007_ _04841_ _04842_ vssd1 vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__nand2_1
XANTENNA__07714__B net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07921__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11958_ _05325_ _05328_ _06003_ vssd1 vssd1 vccd1 vccd1 _06004_ sky130_fd_sc_hd__and3_1
XFILLER_32_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10909_ net196 net1999 net543 vssd1 vssd1 vccd1 vccd1 _00027_ sky130_fd_sc_hd__mux2_1
X_14677_ clknet_leaf_18_clk _01382_ net1108 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11889_ net136 _05956_ _05955_ vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__o21ai_1
X_13628_ clknet_leaf_10_clk _00438_ net1080 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07437__C1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12782__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13559_ clknet_leaf_127_clk _00369_ net1208 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07988__B1 _02820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07080_ datapath.rf.registers\[25\]\[29\] net842 net811 datapath.rf.registers\[13\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__a22o_1
XANTENNA__11398__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07448__Y _02284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07204__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout129 _06369_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__buf_1
XFILLER_86_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07982_ datapath.rf.registers\[4\]\[11\] net716 net696 datapath.rf.registers\[8\]\[11\]
+ _02806_ vssd1 vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__a221o_1
XFILLER_114_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06933_ net984 net928 vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__and2_1
X_09721_ _03437_ _03536_ vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__xnor2_1
XFILLER_113_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13118__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09901__A1 _04727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06864_ _01689_ _01691_ _01697_ _01699_ vssd1 vssd1 vccd1 vccd1 _01700_ sky130_fd_sc_hd__or4_1
X_09652_ net905 _03563_ net627 _03540_ _04487_ vssd1 vssd1 vccd1 vccd1 _04488_ sky130_fd_sc_hd__a221o_1
XFILLER_82_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07912__B1 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08603_ _02826_ _03438_ _02827_ vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__a21oi_1
X_09583_ _04340_ _04353_ net457 vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__mux2_1
X_06795_ datapath.ru.latched_instruction\[20\] _01493_ net1014 vssd1 vssd1 vccd1 vccd1
+ _01631_ sky130_fd_sc_hd__mux2_1
XANTENNA__12957__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout265_A _05575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08534_ datapath.rf.registers\[25\]\[0\] net843 _01743_ datapath.rf.registers\[26\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03370_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_46_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10275__A1 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08465_ datapath.rf.registers\[7\]\[1\] _01758_ net816 datapath.rf.registers\[21\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03301_ sky130_fd_sc_hd__a22o_1
XFILLER_50_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout432_A net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1174_A net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07416_ datapath.rf.registers\[28\]\[22\] net804 net793 datapath.rf.registers\[31\]\[22\]
+ _02251_ vssd1 vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__a221o_1
XFILLER_11_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12016__A2 _05773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09417__B1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08396_ datapath.rf.registers\[28\]\[2\] net930 _01744_ vssd1 vssd1 vccd1 vccd1 _03232_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07691__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07347_ datapath.rf.registers\[22\]\[24\] net735 net669 datapath.rf.registers\[21\]\[24\]
+ _02182_ vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__a221o_1
XFILLER_6_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07979__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07443__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07278_ net874 _02111_ _02112_ _02113_ vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_154_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12264__Y _06254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout899_A net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09017_ _03851_ _03852_ net338 vssd1 vssd1 vccd1 vccd1 _03853_ sky130_fd_sc_hd__mux2_1
XFILLER_124_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10506__A _05335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11101__S net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold150 net49 vssd1 vssd1 vccd1 vccd1 net1498 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold161 datapath.multiplication_module.multiplier_i\[4\] vssd1 vssd1 vccd1 vccd1
+ net1509 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 screen.counter.currentCt\[20\] vssd1 vssd1 vccd1 vccd1 net1520 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold183 datapath.rf.registers\[0\]\[15\] vssd1 vssd1 vccd1 vccd1 net1531 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout687_X net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold194 datapath.rf.registers\[14\]\[21\] vssd1 vssd1 vccd1 vccd1 net1542 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12721__A _05894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout630 _01706_ vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__buf_4
Xfanout641 _01627_ vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__clkbuf_2
Xfanout652 net653 vssd1 vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__buf_2
X_09919_ _01585_ net899 net992 vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__and3_1
XFILLER_144_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout663 _01835_ vssd1 vssd1 vccd1 vccd1 net663 sky130_fd_sc_hd__buf_2
Xfanout674 _01830_ vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08156__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout854_X net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout685 net686 vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__clkbuf_8
XFILLER_19_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_70_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12930_ net260 net1601 net397 vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__mux2_1
Xfanout696 net697 vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__buf_4
XFILLER_37_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07903__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08349__C _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12861_ net169 net2325 net487 vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__mux2_1
XANTENNA__12867__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14600_ clknet_leaf_65_clk _01305_ net1235 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11812_ datapath.ru.latched_instruction\[18\] net333 net314 _01453_ vssd1 vssd1 vccd1
+ vccd1 _00678_ sky130_fd_sc_hd__a22o_1
X_12792_ net176 net2346 net497 vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__mux2_1
XFILLER_15_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14531_ clknet_leaf_138_clk _01236_ net1100 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_42_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11743_ net1469 net145 net141 _03227_ vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__a22o_1
XFILLER_42_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14462_ clknet_leaf_149_clk _01167_ net1060 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_42_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11674_ _05281_ net154 net150 net1409 vssd1 vssd1 vccd1 vccd1 _00559_ sky130_fd_sc_hd__a22o_1
X_13413_ clknet_leaf_121_clk _00223_ net1192 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10625_ net122 net121 net124 net123 vssd1 vssd1 vccd1 vccd1 _05445_ sky130_fd_sc_hd__or4b_4
X_14393_ clknet_leaf_9_clk _01098_ net1072 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11766__B2 _02090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07549__X _02385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10556_ _05380_ _05382_ vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__nand2_1
X_13344_ clknet_leaf_135_clk _00154_ net1089 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_40_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14017__RESET_B net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13275_ clknet_leaf_45_clk _00085_ net1146 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10487_ screen.controlBus\[7\] screen.controlBus\[6\] _05316_ vssd1 vssd1 vccd1 vccd1
+ _05317_ sky130_fd_sc_hd__or3_1
XANTENNA__11011__S net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09764__X _04600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_12_0_clk_X clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12226_ _06168_ _06226_ _06227_ vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_90_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10135__B _04023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10850__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12157_ _06155_ net601 net1276 vssd1 vssd1 vccd1 vccd1 _06185_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_9_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11108_ net261 net2072 net429 vssd1 vssd1 vccd1 vccd1 _00163_ sky130_fd_sc_hd__mux2_1
X_12088_ screen.register.currentXbus\[14\] _05768_ _05772_ screen.register.currentXbus\[30\]
+ vssd1 vssd1 vccd1 vccd1 _06127_ sky130_fd_sc_hd__a22o_1
XFILLER_84_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11039_ net261 net1831 net433 vssd1 vssd1 vccd1 vccd1 _00099_ sky130_fd_sc_hd__mux2_1
XFILLER_77_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12777__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06580_ screen.register.cFill2 vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_121_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06628__X _01467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06775__S net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08250_ datapath.rf.registers\[16\]\[5\] net861 net815 datapath.rf.registers\[21\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03086_ sky130_fd_sc_hd__a22o_1
XANTENNA__07673__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07201_ datapath.rf.registers\[14\]\[27\] net775 net743 datapath.rf.registers\[2\]\[27\]
+ _02034_ vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__a221o_1
XFILLER_32_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08181_ datapath.rf.registers\[16\]\[7\] net740 net673 datapath.rf.registers\[7\]\[7\]
+ _03016_ vssd1 vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__a221o_1
XANTENNA__11757__B2 _02542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07132_ datapath.rf.registers\[24\]\[28\] net859 net812 datapath.rf.registers\[13\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__a22o_1
XFILLER_145_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xteam_04_1305 vssd1 vssd1 vccd1 vccd1 team_04_1305/HI gpio_oeb[14] sky130_fd_sc_hd__conb_1
XANTENNA__07425__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08291__A net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xteam_04_1316 vssd1 vssd1 vccd1 vccd1 team_04_1316/HI gpio_out[20] sky130_fd_sc_hd__conb_1
XFILLER_146_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xteam_04_1327 vssd1 vssd1 vccd1 vccd1 team_04_1327/HI gpio_out[31] sky130_fd_sc_hd__conb_1
Xteam_04_1338 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] team_04_1338/LO sky130_fd_sc_hd__conb_1
X_07063_ datapath.rf.registers\[19\]\[30\] net732 net689 datapath.rf.registers\[31\]\[30\]
+ _01898_ vssd1 vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__a221o_1
XANTENNA__10326__A _04207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09178__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08386__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_151_Right_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08925__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06810__Y _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07965_ datapath.rf.registers\[30\]\[11\] net834 _02775_ _02776_ _02789_ vssd1 vssd1
+ vccd1 vccd1 _02801_ sky130_fd_sc_hd__a2111oi_1
XANTENNA_fanout382_A net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08138__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12260__B _04338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09704_ _03568_ _04539_ net580 vssd1 vssd1 vccd1 vccd1 _04540_ sky130_fd_sc_hd__o21ai_1
X_06916_ _01731_ _01734_ _01736_ _01751_ vssd1 vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_52_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07896_ datapath.rf.registers\[6\]\[12\] net825 net814 datapath.rf.registers\[23\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__a22o_1
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_4_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09635_ _03559_ _03561_ vssd1 vssd1 vccd1 vccd1 _04471_ sky130_fd_sc_hd__xnor2_1
XFILLER_56_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06847_ datapath.ru.latched_instruction\[28\] _01600_ _01602_ datapath.ru.latched_instruction\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01683_ sky130_fd_sc_hd__a22o_1
XFILLER_71_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout647_A _01609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06778_ datapath.ru.latched_instruction\[13\] _01446_ net1016 vssd1 vssd1 vccd1 vccd1
+ _01615_ sky130_fd_sc_hd__mux2_1
X_09566_ net906 _03556_ net626 _03543_ _04401_ vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__a221oi_1
XFILLER_82_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07370__A net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11604__B net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08517_ datapath.rf.registers\[28\]\[1\] net964 net911 _01795_ vssd1 vssd1 vccd1
+ vccd1 _03353_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout814_A _01760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout435_X net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09497_ _03637_ _04329_ _04332_ vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1177_X net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_156_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08448_ datapath.rf.registers\[30\]\[2\] net761 net678 datapath.rf.registers\[29\]\[2\]
+ _03283_ vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_156_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08379_ datapath.rf.registers\[30\]\[3\] net761 net716 datapath.rf.registers\[4\]\[3\]
+ _03214_ vssd1 vssd1 vccd1 vccd1 _03215_ sky130_fd_sc_hd__a221o_1
XFILLER_109_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11748__B2 _02980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10410_ net559 _03359_ net623 vssd1 vssd1 vccd1 vccd1 _05246_ sky130_fd_sc_hd__a21oi_1
XFILLER_136_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07416__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11390_ datapath.rf.registers\[13\]\[13\] _05582_ net411 vssd1 vssd1 vccd1 vccd1
+ _00431_ sky130_fd_sc_hd__mux2_1
XFILLER_137_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10341_ datapath.PC\[14\] net1255 _05174_ _05176_ vssd1 vssd1 vccd1 vccd1 _05177_
+ sky130_fd_sc_hd__o22a_1
XFILLER_136_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13060_ net171 net2221 net474 vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__mux2_1
X_10272_ net466 _04537_ vssd1 vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__nand2_1
XFILLER_140_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout971_X net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12011_ _05840_ _06052_ _06054_ net1001 vssd1 vssd1 vccd1 vccd1 _06055_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_72_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08377__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08129__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout460 net462 vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__buf_2
Xfanout471 net473 vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__clkbuf_8
XFILLER_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout482 _06554_ vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__buf_6
XANTENNA__07264__B net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13962_ clknet_leaf_107_clk _00740_ net1223 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[5\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout493 _06551_ vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12913_ net1769 net241 net484 vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__mux2_1
X_13893_ clknet_leaf_49_clk keypad.decode.button_n\[4\] net1176 vssd1 vssd1 vccd1
+ vccd1 button\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_46_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12844_ net252 net2511 net486 vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07711__C net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12775_ net267 net2274 net496 vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__mux2_1
XANTENNA__08301__B1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11006__S net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14514_ clknet_leaf_33_clk _01219_ net1123 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11726_ net12 net1035 net1025 mmio.memload_or_instruction\[19\] vssd1 vssd1 vccd1
+ vccd1 _00607_ sky130_fd_sc_hd__a22o_1
XFILLER_15_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08852__A1 _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14445_ clknet_leaf_124_clk _01150_ net1207 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11657_ button\[2\] _05874_ vssd1 vssd1 vccd1 vccd1 _05878_ sky130_fd_sc_hd__and2_1
XANTENNA__09919__B net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10608_ net38 _05379_ _05381_ vssd1 vssd1 vccd1 vccd1 _05428_ sky130_fd_sc_hd__and3_2
X_14376_ clknet_leaf_64_clk _01081_ net1236 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06624__A mmio.memload_or_instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11588_ _05807_ _05808_ _05811_ vssd1 vssd1 vccd1 vccd1 _05812_ sky130_fd_sc_hd__or3_1
XANTENNA__10411__A1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13327_ clknet_leaf_27_clk _00137_ net1132 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold908 datapath.rf.registers\[19\]\[0\] vssd1 vssd1 vccd1 vccd1 net2256 sky130_fd_sc_hd__dlygate4sd3_1
Xhold919 datapath.rf.registers\[0\]\[1\] vssd1 vssd1 vccd1 vccd1 net2267 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08080__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10539_ datapath.multiplication_module.mul_prev net615 vssd1 vssd1 vccd1 vccd1 _05367_
+ sky130_fd_sc_hd__nor2_2
XANTENNA__10962__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13258_ clknet_leaf_61_clk _00068_ net1166 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08368__B1 _03203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12209_ _06215_ _06216_ vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__nor2_1
XFILLER_97_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09654__B _04486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13189_ net2179 vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__clkbuf_1
XFILLER_111_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09317__C1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07750_ _02571_ _02572_ _02584_ _02585_ vssd1 vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__or4_1
X_06701_ _01488_ _01509_ _01539_ vssd1 vssd1 vccd1 vccd1 _01540_ sky130_fd_sc_hd__or3_1
XFILLER_38_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07681_ datapath.rf.registers\[6\]\[17\] net825 _02498_ _02503_ _02504_ vssd1 vssd1
+ vccd1 vccd1 _02517_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11675__B1 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08540__B1 _01772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06632_ net1287 net1282 datapath.ru.latched_instruction\[19\] mmio.memload_or_instruction\[19\]
+ vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__or4b_1
X_09420_ net328 _04028_ _03623_ vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__o21a_1
XFILLER_18_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07190__A _02025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06563_ columns.count\[4\] vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__inv_2
X_09351_ _04185_ _04186_ vssd1 vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__nand2_1
XFILLER_80_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08302_ datapath.rf.registers\[2\]\[4\] net887 net790 datapath.rf.registers\[18\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__a22o_1
X_09282_ net556 _04088_ _04117_ _04086_ net632 vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__a32o_2
XTAP_TAPCELL_ROW_138_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07646__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08843__A1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08233_ datapath.rf.registers\[4\]\[6\] net714 net691 datapath.rf.registers\[13\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03069_ sky130_fd_sc_hd__a22o_1
XFILLER_138_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout130_A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13131__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07189__X _02025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08164_ _02997_ _02998_ _02999_ vssd1 vssd1 vccd1 vccd1 _03000_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_151_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07115_ datapath.rf.registers\[2\]\[29\] net743 net684 datapath.rf.registers\[27\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__a22o_1
XFILLER_109_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12970__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08095_ datapath.rf.registers\[22\]\[9\] net736 net708 datapath.rf.registers\[10\]\[9\]
+ _02914_ vssd1 vssd1 vccd1 vccd1 _02931_ sky130_fd_sc_hd__a221o_1
XANTENNA__08071__A2 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload70 clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 clkload70/Y sky130_fd_sc_hd__inv_8
XANTENNA_fanout1137_A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07046_ datapath.rf.registers\[9\]\[30\] net886 net854 datapath.rf.registers\[19\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__a22o_1
Xclkload81 clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 clkload81/Y sky130_fd_sc_hd__inv_6
Xclkload92 clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 clkload92/X sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout597_A net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08997_ net370 _03632_ vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout385_X net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout764_A net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07948_ datapath.rf.registers\[23\]\[11\] net941 net924 vssd1 vssd1 vccd1 vccd1 _02784_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout931_A net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07879_ datapath.rf.registers\[4\]\[13\] net715 net669 datapath.rf.registers\[21\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1294_X net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08531__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09618_ _04450_ _04452_ _04453_ _04430_ net631 vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__a32o_1
X_10890_ datapath.PC\[23\] _05629_ vssd1 vssd1 vccd1 vccd1 _05637_ sky130_fd_sc_hd__nor2_1
XANTENNA__07885__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08196__A _03009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09549_ net375 _03985_ _04384_ vssd1 vssd1 vccd1 vccd1 _04385_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout817_X net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07637__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12560_ _06410_ _06411_ _06412_ vssd1 vssd1 vccd1 vccd1 _06414_ sky130_fd_sc_hd__o21ai_1
XFILLER_140_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11511_ _05331_ _05349_ vssd1 vssd1 vccd1 vccd1 _05736_ sky130_fd_sc_hd__nand2_1
XFILLER_11_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12491_ net256 net2488 net508 vssd1 vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__mux2_1
XANTENNA__13041__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14230_ clknet_leaf_42_clk _00951_ net1144 vssd1 vssd1 vccd1 vccd1 columns.count\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07099__X _01935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11442_ _05712_ _05724_ vssd1 vssd1 vccd1 vccd1 _05732_ sky130_fd_sc_hd__or2_1
XFILLER_125_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11373_ net173 net1675 net519 vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__mux2_1
XANTENNA__12880__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14161_ clknet_leaf_65_clk _00916_ net1235 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08062__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10944__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10324_ _03741_ _05159_ net1040 vssd1 vssd1 vccd1 vccd1 _05160_ sky130_fd_sc_hd__a21oi_1
X_13112_ net241 net2023 net471 vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__mux2_1
X_14092_ clknet_leaf_110_clk _00858_ net1202 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11496__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10255_ _04564_ _05086_ _05090_ net223 vssd1 vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__a211oi_1
X_13043_ net253 net1741 net474 vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__mux2_1
XFILLER_3_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1200 net1203 vssd1 vssd1 vccd1 vccd1 net1200 sky130_fd_sc_hd__buf_2
Xfanout1211 net1213 vssd1 vssd1 vccd1 vccd1 net1211 sky130_fd_sc_hd__clkbuf_4
XFILLER_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10186_ net466 _05021_ _04999_ vssd1 vssd1 vccd1 vccd1 _05022_ sky130_fd_sc_hd__a21o_1
Xfanout1222 net1231 vssd1 vssd1 vccd1 vccd1 net1222 sky130_fd_sc_hd__clkbuf_4
XFILLER_120_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1233 net1234 vssd1 vssd1 vccd1 vccd1 net1233 sky130_fd_sc_hd__buf_2
Xfanout1244 net1250 vssd1 vssd1 vccd1 vccd1 net1244 sky130_fd_sc_hd__buf_4
Xfanout1255 net1256 vssd1 vssd1 vccd1 vccd1 net1255 sky130_fd_sc_hd__clkbuf_4
XFILLER_121_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1266 datapath.PC\[12\] vssd1 vssd1 vccd1 vccd1 net1266 sky130_fd_sc_hd__buf_2
Xfanout1277 screen.counter.ct\[8\] vssd1 vssd1 vccd1 vccd1 net1277 sky130_fd_sc_hd__clkbuf_2
Xfanout1288 net1289 vssd1 vssd1 vccd1 vccd1 net1288 sky130_fd_sc_hd__clkbuf_2
Xfanout290 net291 vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__clkbuf_2
X_13945_ clknet_leaf_111_clk _00723_ net1202 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08522__B1 _03324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload6_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13876_ clknet_leaf_52_clk _00680_ net1184 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_35_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07876__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12827_ net2287 net175 net492 vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__mux2_1
XANTENNA__07089__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12082__B1 _06018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12758_ net1704 net187 net403 vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__mux2_1
XFILLER_61_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08834__A _01586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11709_ net24 net1035 net1025 net1448 vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_62_Left_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12689_ net499 _06520_ _06521_ net503 net2057 vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__a32o_1
XFILLER_129_931 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14428_ clknet_leaf_7_clk _01133_ net1073 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_116_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12790__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold705 datapath.rf.registers\[4\]\[13\] vssd1 vssd1 vccd1 vccd1 net2053 sky130_fd_sc_hd__dlygate4sd3_1
X_14359_ clknet_leaf_127_clk _01064_ net1211 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold716 datapath.rf.registers\[30\]\[9\] vssd1 vssd1 vccd1 vccd1 net2064 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10935__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold727 datapath.mulitply_result\[9\] vssd1 vssd1 vccd1 vccd1 net2075 sky130_fd_sc_hd__dlygate4sd3_1
Xhold738 datapath.rf.registers\[30\]\[28\] vssd1 vssd1 vccd1 vccd1 net2086 sky130_fd_sc_hd__dlygate4sd3_1
Xhold749 datapath.rf.registers\[2\]\[0\] vssd1 vssd1 vccd1 vccd1 net2097 sky130_fd_sc_hd__dlygate4sd3_1
X_08920_ net637 _03480_ _03727_ vssd1 vssd1 vccd1 vccd1 _03756_ sky130_fd_sc_hd__nand3_1
XANTENNA__07013__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10699__A1 _03170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08851_ _02218_ net444 _03686_ vssd1 vssd1 vccd1 vccd1 _03687_ sky130_fd_sc_hd__o21a_1
XFILLER_112_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_71_Left_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07802_ datapath.rf.registers\[4\]\[14\] net958 net933 vssd1 vssd1 vccd1 vccd1 _02638_
+ sky130_fd_sc_hd__and3_1
XFILLER_111_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08782_ net967 _03171_ _03615_ vssd1 vssd1 vccd1 vccd1 _03618_ sky130_fd_sc_hd__mux2_1
XFILLER_38_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09305__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07733_ datapath.rf.registers\[30\]\[16\] net758 net750 datapath.rf.registers\[28\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__a22o_1
XFILLER_53_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13126__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout178_A _05670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07664_ datapath.rf.registers\[19\]\[17\] net973 net927 vssd1 vssd1 vccd1 vccd1 _02500_
+ sky130_fd_sc_hd__and3_1
XFILLER_26_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09403_ net555 _04211_ _04212_ _04238_ _04209_ vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__a41o_2
X_06615_ net1286 net1285 mmio.memload_or_instruction\[18\] vssd1 vssd1 vccd1 vccd1
+ _01454_ sky130_fd_sc_hd__or3b_1
XFILLER_53_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12965__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07595_ datapath.rf.registers\[22\]\[19\] net736 net662 datapath.rf.registers\[5\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__a22o_1
XFILLER_111_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1087_A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09334_ _02567_ _02588_ net625 vssd1 vssd1 vccd1 vccd1 _04170_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07619__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08816__A1 _03358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_80_Left_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_0_0_clk_X clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09265_ net551 net547 _02418_ vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout133_X net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout512_A _05735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1254_A net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08463__B net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08216_ datapath.rf.registers\[13\]\[6\] net810 net793 datapath.rf.registers\[31\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__a22o_1
X_09196_ _04031_ vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__inv_2
XANTENNA__13755__RESET_B net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08147_ net611 _02980_ _02982_ vssd1 vssd1 vccd1 vccd1 _02983_ sky130_fd_sc_hd__o21ai_2
XANTENNA_fanout1042_X net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07252__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08078_ datapath.rf.registers\[12\]\[9\] net756 net673 datapath.rf.registers\[7\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02914_ sky130_fd_sc_hd__a22o_1
XFILLER_1_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout881_A _01721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07029_ datapath.rf.registers\[11\]\[30\] net987 net938 vssd1 vssd1 vccd1 vccd1 _01865_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout979_A net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10073__X _04909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10040_ _04815_ _04875_ vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07004__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold10 keypad.debounce.debounce\[1\] vssd1 vssd1 vccd1 vccd1 net1358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 keypad.debounce.debounce\[7\] vssd1 vssd1 vccd1 vccd1 net1369 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout767_X net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold32 screen.controlBus\[11\] vssd1 vssd1 vccd1 vccd1 net1380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 net110 vssd1 vssd1 vccd1 vccd1 net1391 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 net61 vssd1 vssd1 vccd1 vccd1 net1402 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 screen.controlBus\[20\] vssd1 vssd1 vccd1 vccd1 net1413 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 screen.controlBus\[31\] vssd1 vssd1 vccd1 vccd1 net1424 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 net114 vssd1 vssd1 vccd1 vccd1 net1435 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout934_X net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11991_ _05335_ _05825_ _06030_ net1010 _06035_ vssd1 vssd1 vccd1 vccd1 _06036_ sky130_fd_sc_hd__a221o_1
Xhold98 datapath.multiplication_module.multiplier_i\[10\] vssd1 vssd1 vccd1 vccd1
+ net1446 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12300__B2 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13036__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13730_ clknet_leaf_151_clk _00540_ net1056 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10942_ net901 _04664_ _05681_ vssd1 vssd1 vccd1 vccd1 _05682_ sky130_fd_sc_hd__o21ai_4
XANTENNA__07858__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07261__C net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13661_ clknet_leaf_147_clk _00471_ net1060 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_119_Left_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10873_ _01493_ net617 _05621_ _05622_ vssd1 vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__a22o_2
XANTENNA__12875__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12612_ datapath.mulitply_result\[17\] datapath.multiplication_module.multiplicand_i\[17\]
+ vssd1 vssd1 vccd1 vccd1 _06457_ sky130_fd_sc_hd__and2_1
XFILLER_25_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13592_ clknet_leaf_6_clk _00402_ net1068 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12543_ net500 _06398_ _06399_ net504 net2125 vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__a32o_1
XANTENNA__08283__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07491__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12474_ net164 _05996_ net126 screen.register.currentXbus\[30\] vssd1 vssd1 vccd1
+ vccd1 _00876_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_clkbuf_leaf_91_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14213_ clknet_leaf_48_clk datapath.multiplication_module.multiplicand_i_n\[24\]
+ net1177 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_11425_ net247 net2049 net515 vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__mux2_1
XFILLER_126_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08035__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_7 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07243__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14144_ clknet_leaf_10_clk _00901_ net1080 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_128_Left_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11356_ net255 net1810 net518 vssd1 vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__mux2_1
XANTENNA__06902__A net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10307_ _04855_ _04856_ vssd1 vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__and2b_1
X_14075_ clknet_leaf_121_clk _00842_ net1199 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11287_ net255 net2160 net524 vssd1 vssd1 vccd1 vccd1 _00335_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13026_ net1853 net170 net390 vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__mux2_1
XANTENNA__09535__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10238_ _04909_ _05073_ vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__or2_1
Xfanout1030 net1032 vssd1 vssd1 vccd1 vccd1 net1030 sky130_fd_sc_hd__buf_4
Xfanout1041 net1042 vssd1 vssd1 vccd1 vccd1 net1041 sky130_fd_sc_hd__clkbuf_2
X_10169_ net1043 _03742_ vssd1 vssd1 vccd1 vccd1 _05005_ sky130_fd_sc_hd__nand2_1
Xfanout1052 net1058 vssd1 vssd1 vccd1 vccd1 net1052 sky130_fd_sc_hd__clkbuf_4
Xfanout1063 net1066 vssd1 vssd1 vccd1 vccd1 net1063 sky130_fd_sc_hd__clkbuf_2
XFILLER_67_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1074 net1075 vssd1 vssd1 vccd1 vccd1 net1074 sky130_fd_sc_hd__buf_2
Xfanout1085 net1092 vssd1 vssd1 vccd1 vccd1 net1085 sky130_fd_sc_hd__clkbuf_4
Xfanout1096 net1101 vssd1 vssd1 vccd1 vccd1 net1096 sky130_fd_sc_hd__clkbuf_2
XFILLER_35_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13928_ clknet_leaf_110_clk _00706_ net1202 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07452__B net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_137_Left_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07849__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14213__RESET_B net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13859_ clknet_leaf_53_clk _00663_ net1183 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07171__C net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12785__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_44_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12055__B1 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07380_ _02211_ _02213_ _02214_ _02215_ vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__nor4_1
XFILLER_31_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08274__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09471__A1 _03009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09050_ net459 _03884_ _03885_ vssd1 vssd1 vccd1 vccd1 _03886_ sky130_fd_sc_hd__and3_1
XANTENNA__07482__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_59_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08001_ datapath.rf.registers\[5\]\[10\] net947 net935 vssd1 vssd1 vccd1 vccd1 _02837_
+ sky130_fd_sc_hd__and3_1
XFILLER_117_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08026__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold502 datapath.rf.registers\[31\]\[3\] vssd1 vssd1 vccd1 vccd1 net1850 sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 datapath.rf.registers\[29\]\[3\] vssd1 vssd1 vccd1 vccd1 net1861 sky130_fd_sc_hd__dlygate4sd3_1
Xhold524 datapath.rf.registers\[28\]\[18\] vssd1 vssd1 vccd1 vccd1 net1872 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold535 datapath.rf.registers\[6\]\[16\] vssd1 vssd1 vccd1 vccd1 net1883 sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 datapath.rf.registers\[28\]\[25\] vssd1 vssd1 vccd1 vccd1 net1894 sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 datapath.rf.registers\[23\]\[30\] vssd1 vssd1 vccd1 vccd1 net1905 sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 columns.count\[5\] vssd1 vssd1 vccd1 vccd1 net1916 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold579 datapath.rf.registers\[13\]\[20\] vssd1 vssd1 vccd1 vccd1 net1927 sky130_fd_sc_hd__dlygate4sd3_1
X_09952_ _04777_ _04787_ _04776_ vssd1 vssd1 vccd1 vccd1 _04788_ sky130_fd_sc_hd__a21o_1
XFILLER_131_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08903_ net1266 datapath.PC\[13\] _03738_ vssd1 vssd1 vccd1 vccd1 _03739_ sky130_fd_sc_hd__or3_1
XANTENNA_clkbuf_leaf_117_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09883_ _04717_ _04718_ vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout295_A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1202 screen.register.currentYbus\[3\] vssd1 vssd1 vccd1 vccd1 net2550 sky130_fd_sc_hd__dlygate4sd3_1
X_08834_ _01586_ net897 vssd1 vssd1 vccd1 vccd1 _03670_ sky130_fd_sc_hd__nor2_2
XFILLER_58_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09842__B _03419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1213 screen.register.currentYbus\[17\] vssd1 vssd1 vccd1 vccd1 net2561 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1224 datapath.rf.registers\[26\]\[0\] vssd1 vssd1 vccd1 vccd1 net2572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1235 datapath.rf.registers\[18\]\[11\] vssd1 vssd1 vccd1 vccd1 net2583 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1246 datapath.rf.registers\[8\]\[0\] vssd1 vssd1 vccd1 vccd1 net2594 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1257 datapath.rf.registers\[24\]\[25\] vssd1 vssd1 vccd1 vccd1 net2605 sky130_fd_sc_hd__dlygate4sd3_1
X_08765_ _01601_ _01603_ _01604_ vssd1 vssd1 vccd1 vccd1 _03601_ sky130_fd_sc_hd__and3b_2
Xhold1268 datapath.rf.registers\[29\]\[22\] vssd1 vssd1 vccd1 vccd1 net2616 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1279 datapath.rf.registers\[28\]\[12\] vssd1 vssd1 vccd1 vccd1 net2627 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07362__B net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07716_ datapath.rf.registers\[12\]\[16\] net826 net801 datapath.rf.registers\[3\]\[16\]
+ _02547_ vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__a221o_1
XFILLER_26_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08696_ _02805_ _02825_ vssd1 vssd1 vccd1 vccd1 _03532_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_49_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07647_ datapath.rf.registers\[11\]\[18\] net710 net671 datapath.rf.registers\[7\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02483_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout250_X net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout727_A _01812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07578_ _02397_ _02411_ _02412_ _02413_ vssd1 vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__or4_1
XFILLER_139_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09317_ _02418_ net440 _04151_ net369 vssd1 vssd1 vccd1 vccd1 _04153_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_62_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08265__A2 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout515_X net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09462__A1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08193__B _01784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1257_X net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11104__S net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07473__B1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09248_ net632 _04058_ _04060_ _04083_ vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__a22o_2
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08017__A2 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_10_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_10_0_clk sky130_fd_sc_hd__clkbuf_8
X_09179_ net905 _03502_ _04014_ vssd1 vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__a21oi_1
XFILLER_147_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07225__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11210_ net288 net2381 net529 vssd1 vssd1 vccd1 vccd1 _00260_ sky130_fd_sc_hd__mux2_1
X_12190_ net2604 _06179_ _06204_ vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__a21o_1
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout884_X net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11141_ net209 net2572 net532 vssd1 vssd1 vccd1 vccd1 _00194_ sky130_fd_sc_hd__mux2_1
Xoutput44 net44 vssd1 vssd1 vccd1 vccd1 ADR_O[13] sky130_fd_sc_hd__buf_2
Xoutput55 net55 vssd1 vssd1 vccd1 vccd1 ADR_O[23] sky130_fd_sc_hd__buf_2
XFILLER_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 ADR_O[4] sky130_fd_sc_hd__buf_2
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 DAT_O[13] sky130_fd_sc_hd__buf_2
X_11072_ _05518_ _05713_ vssd1 vssd1 vccd1 vccd1 _05714_ sky130_fd_sc_hd__or2_1
Xoutput88 net88 vssd1 vssd1 vccd1 vccd1 DAT_O[23] sky130_fd_sc_hd__buf_2
XFILLER_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput99 net99 vssd1 vssd1 vccd1 vccd1 DAT_O[4] sky130_fd_sc_hd__buf_2
XANTENNA__12730__Y _06549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10023_ _04803_ _04858_ vssd1 vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08649__A _01980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input23_A DAT_I[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11974_ net1006 _05770_ vssd1 vssd1 vccd1 vccd1 _06019_ sky130_fd_sc_hd__nor2_2
XANTENNA__09150__A0 _02217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13713_ clknet_leaf_35_clk _00523_ net1127 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10925_ _05665_ _05666_ vssd1 vssd1 vccd1 vccd1 _05667_ sky130_fd_sc_hd__nor2_1
X_14693_ clknet_leaf_119_clk _01398_ net1191 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13644_ clknet_leaf_15_clk _00454_ net1103 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10856_ _04600_ _05607_ net901 vssd1 vssd1 vccd1 vccd1 _05608_ sky130_fd_sc_hd__mux2_2
X_13575_ clknet_leaf_145_clk _00385_ net1086 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08256__A2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09453__A1 _02805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10787_ datapath.PC\[8\] _05542_ vssd1 vssd1 vccd1 vccd1 _05549_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_30_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11014__S net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12526_ datapath.mulitply_result\[3\] datapath.multiplication_module.multiplicand_i\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06385_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_97_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12457_ net164 _05962_ net126 screen.register.currentXbus\[13\] vssd1 vssd1 vccd1
+ vccd1 _00859_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10853__S net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08008__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08390__Y _03226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11408_ net2043 net168 net410 vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__mux2_1
XANTENNA__07216__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12388_ net1527 net133 _06341_ vssd1 vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__a21o_1
XANTENNA__08964__A0 _02750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08550__C _01823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14127_ clknet_leaf_0_clk _00884_ net1054 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11339_ net1724 net174 net416 vssd1 vssd1 vccd1 vccd1 _00384_ sky130_fd_sc_hd__mux2_1
XANTENNA__06989__D _01666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10771__B1 _05534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14058_ clknet_leaf_95_clk _00825_ net1216 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13009_ net1562 net253 net390 vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__mux2_1
X_06880_ net981 net943 vssd1 vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__and2_4
XTAP_TAPCELL_ROW_128_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07463__A net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_145_Left_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08550_ datapath.rf.registers\[13\]\[0\] net969 _01823_ vssd1 vssd1 vccd1 vccd1 _03386_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12276__B1 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07501_ datapath.rf.registers\[18\]\[20\] net973 net949 vssd1 vssd1 vccd1 vccd1 _02337_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_141_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08481_ datapath.rf.registers\[10\]\[1\] net881 net794 datapath.rf.registers\[31\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03317_ sky130_fd_sc_hd__a22o_1
XFILLER_63_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07432_ datapath.rf.registers\[24\]\[22\] net766 net730 datapath.rf.registers\[19\]\[22\]
+ _02265_ vssd1 vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__a221o_1
XANTENNA__12579__A1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07363_ datapath.rf.registers\[7\]\[23\] net940 net932 vssd1 vssd1 vccd1 vccd1 _02199_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_44_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09102_ net344 _03782_ _03937_ net320 vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__a211o_1
XANTENNA__08429__A1_N _01637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_154_Left_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07294_ datapath.rf.registers\[2\]\[25\] net744 net677 datapath.rf.registers\[29\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__a22o_1
XANTENNA__08581__X _03417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09033_ _03590_ _03866_ vssd1 vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout308_A _06246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold310 datapath.rf.registers\[16\]\[6\] vssd1 vssd1 vccd1 vccd1 net1658 sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 datapath.rf.registers\[7\]\[28\] vssd1 vssd1 vccd1 vccd1 net1669 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12263__B net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08955__A0 _02467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold332 datapath.multiplication_module.multiplicand_i\[7\] vssd1 vssd1 vccd1 vccd1
+ net1680 sky130_fd_sc_hd__dlygate4sd3_1
Xhold343 datapath.rf.registers\[14\]\[24\] vssd1 vssd1 vccd1 vccd1 net1691 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10211__C1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07357__B net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold354 datapath.rf.registers\[3\]\[20\] vssd1 vssd1 vccd1 vccd1 net1702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 datapath.rf.registers\[16\]\[4\] vssd1 vssd1 vccd1 vccd1 net1713 sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 datapath.rf.registers\[12\]\[30\] vssd1 vssd1 vccd1 vccd1 net1724 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10762__B1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1217_A net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold387 datapath.rf.registers\[28\]\[19\] vssd1 vssd1 vccd1 vccd1 net1735 sky130_fd_sc_hd__dlygate4sd3_1
Xhold398 datapath.rf.registers\[14\]\[6\] vssd1 vssd1 vccd1 vccd1 net1746 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout801 net802 vssd1 vssd1 vccd1 vccd1 net801 sky130_fd_sc_hd__clkbuf_8
Xfanout812 _01765_ vssd1 vssd1 vccd1 vccd1 net812 sky130_fd_sc_hd__clkbuf_8
X_09935_ _04769_ _04770_ vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__nand2b_1
Xfanout823 _01755_ vssd1 vssd1 vccd1 vccd1 net823 sky130_fd_sc_hd__buf_4
Xfanout834 net835 vssd1 vssd1 vccd1 vccd1 net834 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout677_A net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout845 _01737_ vssd1 vssd1 vccd1 vccd1 net845 sky130_fd_sc_hd__buf_4
Xfanout856 net859 vssd1 vssd1 vccd1 vccd1 net856 sky130_fd_sc_hd__buf_4
Xfanout867 _01724_ vssd1 vssd1 vccd1 vccd1 net867 sky130_fd_sc_hd__clkbuf_4
X_09866_ _03033_ _03081_ vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout1005_X net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout878 _01722_ vssd1 vssd1 vccd1 vccd1 net878 sky130_fd_sc_hd__clkbuf_8
Xhold1010 datapath.rf.registers\[31\]\[11\] vssd1 vssd1 vccd1 vccd1 net2358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1021 datapath.rf.registers\[14\]\[20\] vssd1 vssd1 vccd1 vccd1 net2369 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout889 _01713_ vssd1 vssd1 vccd1 vccd1 net889 sky130_fd_sc_hd__clkbuf_8
XFILLER_133_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08817_ net612 _03417_ _03644_ _03384_ vssd1 vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__a211oi_2
Xhold1032 datapath.rf.registers\[25\]\[17\] vssd1 vssd1 vccd1 vccd1 net2380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1043 datapath.rf.registers\[26\]\[10\] vssd1 vssd1 vccd1 vccd1 net2391 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07804__C net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09797_ _03642_ net347 _04251_ net650 vssd1 vssd1 vccd1 vccd1 _04633_ sky130_fd_sc_hd__o31a_1
XFILLER_100_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1054 datapath.rf.registers\[21\]\[2\] vssd1 vssd1 vccd1 vccd1 net2402 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1065 datapath.rf.registers\[27\]\[27\] vssd1 vssd1 vccd1 vccd1 net2413 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1076 datapath.rf.registers\[1\]\[26\] vssd1 vssd1 vccd1 vccd1 net2424 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1087 datapath.rf.registers\[29\]\[26\] vssd1 vssd1 vccd1 vccd1 net2435 sky130_fd_sc_hd__dlygate4sd3_1
X_08748_ _03507_ _03508_ _03582_ _03505_ vssd1 vssd1 vccd1 vccd1 _03584_ sky130_fd_sc_hd__a31o_1
Xhold1098 datapath.rf.registers\[25\]\[15\] vssd1 vssd1 vccd1 vccd1 net2446 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_54_773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08679_ _02523_ _02543_ vssd1 vssd1 vccd1 vccd1 _03515_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout632_X net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08486__A2 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12019__B1 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10710_ _02633_ _05368_ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i_n\[15\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__07694__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11690_ _04954_ _05885_ net148 net1443 vssd1 vssd1 vccd1 vccd1 _00575_ sky130_fd_sc_hd__a2bb2o_1
X_10641_ _05428_ _05444_ _05457_ _05460_ _05456_ vssd1 vssd1 vccd1 vccd1 _05461_ sky130_fd_sc_hd__o311a_1
XANTENNA__08238__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09435__A1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13360_ clknet_leaf_24_clk _00170_ net1157 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10572_ _02612_ _02660_ _02704_ _02750_ vssd1 vssd1 vccd1 vccd1 _05395_ sky130_fd_sc_hd__or4_1
X_12311_ net896 _04207_ net307 _06288_ vssd1 vssd1 vccd1 vccd1 _06289_ sky130_fd_sc_hd__o211a_1
XANTENNA__09747__B _04272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13291_ clknet_leaf_56_clk _00101_ net1171 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12242_ _06168_ _06236_ _06237_ vssd1 vssd1 vccd1 vccd1 _00776_ sky130_fd_sc_hd__nor3_1
XANTENNA__12742__A1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07267__B net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12173_ net1271 _06193_ _06194_ vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_75_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11124_ net242 net1690 net428 vssd1 vssd1 vccd1 vccd1 _00179_ sky130_fd_sc_hd__mux2_1
XFILLER_150_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11055_ net242 net1653 net432 vssd1 vssd1 vccd1 vccd1 _00115_ sky130_fd_sc_hd__mux2_1
XFILLER_67_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10006_ _04774_ _04791_ vssd1 vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11009__S net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12258__B1 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13858__RESET_B net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11957_ net1007 _05780_ vssd1 vssd1 vccd1 vccd1 _06003_ sky130_fd_sc_hd__nor2_1
XANTENNA__08477__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10908_ net1046 net652 _05651_ _05652_ vssd1 vssd1 vccd1 vccd1 _05653_ sky130_fd_sc_hd__o22a_2
XFILLER_60_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14676_ clknet_leaf_128_clk _01381_ net1210 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11888_ _02876_ net658 vssd1 vssd1 vccd1 vccd1 _05956_ sky130_fd_sc_hd__nand2_1
X_13627_ clknet_leaf_38_clk _00437_ net1145 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10839_ datapath.PC\[15\] datapath.PC\[16\] _05583_ vssd1 vssd1 vccd1 vccd1 _05593_
+ sky130_fd_sc_hd__and3_1
XFILLER_20_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08229__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13558_ clknet_leaf_140_clk _00368_ net1099 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_132_Right_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12509_ net169 net2613 net509 vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__mux2_1
XANTENNA__07988__B2 _02823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10441__C1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13489_ clknet_leaf_39_clk _00299_ net1141 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08561__B net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06660__B2 datapath.ru.latched_instruction\[29\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08937__A0 _01935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07981_ _02812_ _02814_ _02816_ vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__or3_1
X_09720_ _04549_ _04550_ _04555_ _03673_ vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__a2bb2o_1
X_06932_ net929 net920 vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_126_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09651_ _03008_ _03030_ _03721_ vssd1 vssd1 vccd1 vccd1 _04487_ sky130_fd_sc_hd__o21a_1
XFILLER_83_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06863_ _01662_ _01669_ _01680_ _01698_ vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__or4_1
X_08602_ _02881_ _03431_ _03435_ _02880_ vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__a31o_1
X_09582_ net460 _04345_ _04417_ vssd1 vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__a21oi_1
X_06794_ _01451_ net1002 net1018 net1027 datapath.ru.latched_instruction\[17\] vssd1
+ vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__a32o_4
X_08533_ datapath.rf.registers\[17\]\[0\] net852 _03365_ _03368_ vssd1 vssd1 vccd1
+ vccd1 _03369_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout160_A net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08468__A2 _01713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13134__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout258_A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08464_ datapath.rf.registers\[13\]\[1\] net988 net918 vssd1 vssd1 vccd1 vccd1 _03300_
+ sky130_fd_sc_hd__and3_1
X_07415_ datapath.rf.registers\[27\]\[22\] net807 net799 datapath.rf.registers\[15\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__a22o_1
XFILLER_11_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08395_ _03204_ _03228_ vssd1 vssd1 vccd1 vccd1 _03231_ sky130_fd_sc_hd__and2_1
XANTENNA__12973__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07346_ datapath.rf.registers\[9\]\[24\] net703 net661 datapath.rf.registers\[5\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__a22o_1
XFILLER_149_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07277_ datapath.rf.registers\[18\]\[25\] net791 _02096_ _02098_ _02110_ vssd1 vssd1
+ vccd1 vccd1 _02113_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_154_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09016_ _03682_ _03689_ net342 vssd1 vssd1 vccd1 vccd1 _03852_ sky130_fd_sc_hd__mux2_1
XFILLER_145_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout794_A net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold140 net103 vssd1 vssd1 vccd1 vccd1 net1488 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 net94 vssd1 vssd1 vccd1 vccd1 net1499 sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 datapath.ru.n_memwrite vssd1 vssd1 vccd1 vccd1 net1510 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold173 datapath.multiplication_module.multiplicand_i\[28\] vssd1 vssd1 vccd1 vccd1
+ net1521 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold184 mmio.memload_or_instruction\[23\] vssd1 vssd1 vccd1 vccd1 net1532 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07600__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold195 datapath.rf.registers\[4\]\[30\] vssd1 vssd1 vccd1 vccd1 net1543 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout620 net622 vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__buf_2
Xfanout631 net633 vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__clkbuf_4
XFILLER_120_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout642 _01622_ vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__buf_2
X_09918_ _01643_ net630 vssd1 vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__nor2_1
Xfanout653 net654 vssd1 vssd1 vccd1 vccd1 net653 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout664 net667 vssd1 vssd1 vccd1 vccd1 net664 sky130_fd_sc_hd__buf_4
Xfanout675 net678 vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout686 _01827_ vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09849_ net566 _01856_ vssd1 vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__nand2_1
Xfanout697 _01822_ vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__buf_4
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout847_X net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12860_ net172 net1985 net488 vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__mux2_1
XFILLER_85_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11811_ datapath.ru.latched_instruction\[17\] net333 net314 _01451_ vssd1 vssd1 vccd1
+ vccd1 _00677_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_1_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ net185 net2254 net495 vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__mux2_1
XFILLER_27_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09656__A1 _03604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13044__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14530_ clknet_leaf_151_clk _01235_ net1052 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11742_ net1425 net147 net142 _03292_ vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__a22o_1
XFILLER_30_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07131__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14461_ clknet_leaf_144_clk _01166_ net1085 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12883__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11673_ _05211_ net154 net150 net1421 vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__a22o_1
X_13412_ clknet_leaf_21_clk _00222_ net1164 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10624_ net122 net121 net123 net124 vssd1 vssd1 vccd1 vccd1 _05444_ sky130_fd_sc_hd__or4b_4
X_14392_ clknet_leaf_6_clk _01097_ net1068 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08662__A _02217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11499__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13343_ clknet_leaf_13_clk _00153_ net1078 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10555_ net37 net38 vssd1 vssd1 vccd1 vccd1 _05382_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_40_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08092__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07278__A net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13274_ clknet_leaf_14_clk _00084_ net1078 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10486_ screen.controlBus\[4\] screen.controlBus\[5\] vssd1 vssd1 vccd1 vccd1 _05316_
+ sky130_fd_sc_hd__or2_1
XFILLER_142_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12225_ screen.counter.currentCt\[11\] screen.counter.currentCt\[12\] _06223_ vssd1
+ vssd1 vccd1 vccd1 _06227_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_90_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07198__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12156_ _06160_ net567 _06179_ _06183_ vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__o211a_1
XANTENNA__06910__A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11107_ net207 net2502 net429 vssd1 vssd1 vccd1 vccd1 _00162_ sky130_fd_sc_hd__mux2_1
XFILLER_96_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12087_ screen.register.currentYbus\[22\] _05773_ net995 screen.register.currentXbus\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06126_ sky130_fd_sc_hd__a22o_1
XFILLER_1_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08147__A1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11038_ net209 net2594 net433 vssd1 vssd1 vccd1 vccd1 _00098_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_108_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09895__A1 _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08837__A _03669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12989_ net185 net1620 net479 vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_121_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14659_ clknet_leaf_119_clk _01364_ net1191 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12793__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07200_ datapath.rf.registers\[3\]\[27\] net770 net763 datapath.rf.registers\[1\]\[27\]
+ _02035_ vssd1 vssd1 vccd1 vccd1 _02036_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_41_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08180_ datapath.rf.registers\[12\]\[7\] net756 net681 datapath.rf.registers\[6\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03016_ sky130_fd_sc_hd__a22o_1
X_07131_ datapath.rf.registers\[28\]\[28\] net806 net800 datapath.rf.registers\[15\]\[28\]
+ _01966_ vssd1 vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__a221o_1
XFILLER_146_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10166__X _05002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_04_1306 vssd1 vssd1 vccd1 vccd1 team_04_1306/HI gpio_oeb[15] sky130_fd_sc_hd__conb_1
Xteam_04_1317 vssd1 vssd1 vccd1 vccd1 team_04_1317/HI gpio_out[21] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_136_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11202__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06633__A1 datapath.ru.latched_instruction\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xteam_04_1328 vssd1 vssd1 vccd1 vccd1 team_04_1328/HI gpio_out[32] sky130_fd_sc_hd__conb_1
X_07062_ datapath.rf.registers\[11\]\[30\] net712 _01897_ net788 vssd1 vssd1 vccd1
+ vccd1 _01898_ sky130_fd_sc_hd__a211o_1
XFILLER_145_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07830__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_04_1339 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] team_04_1339/LO sky130_fd_sc_hd__conb_1
XFILLER_145_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07189__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07475__X _02311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13129__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07964_ _02796_ _02797_ _02798_ _02799_ vssd1 vssd1 vccd1 vccd1 _02800_ sky130_fd_sc_hd__or4_1
XFILLER_101_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09703_ _03537_ _03567_ _03536_ vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__a21oi_1
X_06915_ _01742_ _01747_ _01750_ vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__or3_1
XFILLER_114_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11142__A0 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12968__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07895_ datapath.rf.registers\[7\]\[12\] net817 net816 datapath.rf.registers\[21\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02731_ sky130_fd_sc_hd__a22o_1
X_09634_ _03673_ net337 _04019_ _04467_ _04469_ vssd1 vssd1 vccd1 vccd1 _04470_ sky130_fd_sc_hd__a311o_1
XFILLER_95_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07897__B1 _01765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06846_ _01635_ _01636_ datapath.ru.latched_instruction\[22\] vssd1 vssd1 vccd1 vccd1
+ _01682_ sky130_fd_sc_hd__mux2_1
XFILLER_83_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09565_ _03149_ _03172_ net623 vssd1 vssd1 vccd1 vccd1 _04401_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout542_A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06777_ _01613_ vssd1 vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__inv_2
XANTENNA__09638__B2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08466__B net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08516_ datapath.rf.registers\[7\]\[1\] net970 _01820_ vssd1 vssd1 vccd1 vccd1 _03352_
+ sky130_fd_sc_hd__and3_1
XANTENNA__11604__C net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09496_ net324 _04113_ _04330_ _04331_ vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__o211a_1
XANTENNA__07113__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08447_ datapath.rf.registers\[21\]\[2\] net967 _01831_ net913 net914 vssd1 vssd1
+ vccd1 vccd1 _03283_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_156_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout807_A net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout428_X net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08378_ datapath.rf.registers\[22\]\[3\] net736 net685 datapath.rf.registers\[27\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03214_ sky130_fd_sc_hd__a22o_1
X_07329_ datapath.rf.registers\[7\]\[24\] net817 _02148_ _02152_ _02164_ vssd1 vssd1
+ vccd1 vccd1 _02165_ sky130_fd_sc_hd__a2111o_1
XFILLER_137_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10832__A2_N net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11112__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10340_ net223 _05175_ net1294 vssd1 vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__a21o_1
XFILLER_136_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout797_X net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10271_ _04517_ _04537_ vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__xor2_1
XANTENNA__10804__X _05564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12010_ screen.register.currentXbus\[17\] _05769_ _06019_ screen.register.currentYbus\[9\]
+ _06053_ vssd1 vssd1 vccd1 vccd1 _06054_ sky130_fd_sc_hd__a221o_1
XFILLER_151_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_72_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06730__A _01450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06927__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13039__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout450 net451 vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__clkbuf_4
XFILLER_94_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout461 net462 vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__buf_2
Xfanout472 net473 vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__buf_4
X_13961_ clknet_leaf_107_clk _00739_ net1220 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09877__A1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12878__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout483 _06554_ vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__clkbuf_4
XFILLER_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07264__C net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout494 _06550_ vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__clkbuf_8
X_12912_ net1790 net246 net482 vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__mux2_1
XFILLER_86_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13892_ clknet_leaf_49_clk keypad.decode.button_n\[3\] net1175 vssd1 vssd1 vccd1
+ vccd1 button\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08657__A _02126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12843_ net254 net1739 net487 vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_100_Left_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_87_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12774_ net271 net2625 net496 vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__mux2_1
XFILLER_42_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07104__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14513_ clknet_leaf_39_clk _01218_ net1141 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11725_ net11 net1035 net1025 mmio.memload_or_instruction\[18\] vssd1 vssd1 vccd1
+ vccd1 _00606_ sky130_fd_sc_hd__a22o_1
XFILLER_70_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14444_ clknet_leaf_14_clk _01149_ net1102 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11656_ net1449 _05875_ _05877_ vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__a21o_1
XANTENNA__09919__C net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10607_ screen.register.controlFill screen.register.xFill _05427_ vssd1 vssd1 vccd1
+ vccd1 screen.screenEdge.enableIn sky130_fd_sc_hd__and3_1
XFILLER_128_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14375_ clknet_leaf_140_clk _01080_ net1094 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11587_ _05805_ _05809_ _05810_ vssd1 vssd1 vccd1 vccd1 _05811_ sky130_fd_sc_hd__or3_1
XANTENNA__11022__S net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13326_ clknet_leaf_0_clk _00136_ net1055 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07812__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold909 datapath.rf.registers\[20\]\[1\] vssd1 vssd1 vccd1 vccd1 net2257 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_118_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10538_ _05074_ _05366_ vssd1 vssd1 vccd1 vccd1 mmio.ack_center.key_en sky130_fd_sc_hd__nor2_1
X_13257_ clknet_leaf_20_clk _00067_ net1165 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10469_ net1271 net1272 vssd1 vssd1 vccd1 vccd1 _05299_ sky130_fd_sc_hd__or2_1
XANTENNA__08368__A1 datapath.rf.registers\[0\]\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12208_ net2560 _06214_ net603 vssd1 vssd1 vccd1 vccd1 _06216_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09565__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13188_ datapath.rf.registers\[0\]\[25\] vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07455__B net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12139_ _05761_ net1012 net567 vssd1 vssd1 vccd1 vccd1 _06174_ sky130_fd_sc_hd__a21o_1
XFILLER_29_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07591__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12788__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06700_ _01519_ _01526_ _01531_ _01538_ vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__or4b_1
XFILLER_49_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07879__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07680_ datapath.rf.registers\[7\]\[17\] net818 _02492_ _02501_ _02502_ vssd1 vssd1
+ vccd1 vccd1 _02516_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07343__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06631_ net1287 net1282 mmio.memload_or_instruction\[19\] vssd1 vssd1 vccd1 vccd1
+ _01470_ sky130_fd_sc_hd__or3b_1
XFILLER_80_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09350_ net551 net547 _02612_ vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__a21o_1
XFILLER_52_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08301_ datapath.rf.registers\[17\]\[4\] net852 net833 datapath.rf.registers\[30\]\[4\]
+ net873 vssd1 vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_23_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09281_ net578 _04087_ _04116_ vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_138_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08232_ datapath.rf.registers\[20\]\[6\] net718 net687 datapath.rf.registers\[31\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03068_ sky130_fd_sc_hd__a22o_1
XFILLER_60_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08163_ datapath.rf.registers\[27\]\[7\] net809 _02985_ _02989_ _02990_ vssd1 vssd1
+ vccd1 vccd1 _02999_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10337__A net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09253__C1 _02419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07114_ datapath.rf.registers\[26\]\[29\] net779 net726 datapath.rf.registers\[25\]\[29\]
+ _01949_ vssd1 vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__a221o_1
XFILLER_146_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08094_ _02927_ _02929_ vssd1 vssd1 vccd1 vccd1 _02930_ sky130_fd_sc_hd__nor2_1
Xclkload60 clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 clkload60/Y sky130_fd_sc_hd__inv_6
Xclkload71 clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 clkload71/Y sky130_fd_sc_hd__inv_6
X_07045_ _01877_ _01878_ _01879_ _01880_ vssd1 vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__nor4_1
XFILLER_134_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload82 clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 clkload82/Y sky130_fd_sc_hd__inv_8
Xclkload93 clknet_leaf_114_clk vssd1 vssd1 vccd1 vccd1 clkload93/Y sky130_fd_sc_hd__inv_8
XANTENNA__09556__B1 _03604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout492_A _06551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07365__B net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08996_ _03593_ _03828_ net579 vssd1 vssd1 vccd1 vccd1 _03832_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_149_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07947_ datapath.rf.registers\[7\]\[11\] net941 net934 vssd1 vssd1 vccd1 vccd1 _02783_
+ sky130_fd_sc_hd__and3_1
XFILLER_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07878_ _02707_ _02709_ _02711_ _02713_ vssd1 vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__or4_1
XANTENNA__07334__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09617_ net578 _04451_ net605 vssd1 vssd1 vccd1 vccd1 _04453_ sky130_fd_sc_hd__a21oi_1
XFILLER_141_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06829_ _01505_ net1004 net1020 net1028 datapath.ru.latched_instruction\[21\] vssd1
+ vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__a32oi_4
XANTENNA_fanout924_A net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout545_X net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11107__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09548_ net364 _03763_ _03630_ net370 vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__o211a_1
XANTENNA__07098__B2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08295__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_144_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_144_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09479_ net325 _04107_ _04309_ _04313_ _03639_ vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout712_X net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11510_ net1368 _01426_ net1022 net1506 vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__a22o_1
XFILLER_12_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12490_ net262 net2262 net508 vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__mux2_1
XFILLER_133_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11441_ net168 net2383 net514 vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__mux2_1
XFILLER_137_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12394__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14160_ clknet_leaf_66_clk _00915_ net1240 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11372_ net183 net2562 net518 vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__mux2_1
XFILLER_125_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07259__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11777__S _05894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13111_ net244 net2495 net470 vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__mux2_1
X_10323_ datapath.PC\[15\] _03740_ vssd1 vssd1 vccd1 vccd1 _05159_ sky130_fd_sc_hd__nand2_1
XFILLER_4_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14091_ clknet_leaf_95_clk _00857_ net1227 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12146__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13042_ net254 net1623 net474 vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__mux2_1
XFILLER_79_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10254_ net1040 _05087_ _05089_ net635 vssd1 vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__a211oi_1
XFILLER_133_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1201 net1203 vssd1 vssd1 vccd1 vccd1 net1201 sky130_fd_sc_hd__clkbuf_4
Xfanout1212 net1213 vssd1 vssd1 vccd1 vccd1 net1212 sky130_fd_sc_hd__clkbuf_2
XFILLER_121_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10185_ net1043 _05020_ net635 vssd1 vssd1 vccd1 vccd1 _05021_ sky130_fd_sc_hd__a21oi_1
Xfanout1223 net1225 vssd1 vssd1 vccd1 vccd1 net1223 sky130_fd_sc_hd__clkbuf_4
Xfanout1234 net1251 vssd1 vssd1 vccd1 vccd1 net1234 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07573__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1245 net1249 vssd1 vssd1 vccd1 vccd1 net1245 sky130_fd_sc_hd__clkbuf_4
Xfanout1256 net1257 vssd1 vssd1 vccd1 vccd1 net1256 sky130_fd_sc_hd__buf_2
Xfanout1267 datapath.PC\[9\] vssd1 vssd1 vccd1 vccd1 net1267 sky130_fd_sc_hd__buf_2
Xfanout1278 screen.counter.ct\[7\] vssd1 vssd1 vccd1 vccd1 net1278 sky130_fd_sc_hd__buf_2
Xfanout280 _05554_ vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__clkbuf_2
Xfanout291 net293 vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__clkbuf_2
Xfanout1289 net1290 vssd1 vssd1 vccd1 vccd1 net1289 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13944_ clknet_leaf_110_clk _00722_ net1202 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10710__A _02633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07325__A2 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08522__A1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13875_ clknet_leaf_52_clk _00679_ net1184 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_85_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11017__S net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12826_ net1996 net184 net491 vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__mux2_1
XFILLER_61_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10856__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12757_ net1800 net195 net402 vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__mux2_1
XFILLER_43_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_135_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_135_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09483__C1 _03009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08834__B net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11708_ net13 net1035 net1025 net1529 vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__a22o_1
X_12688_ _06518_ _06519_ _06517_ vssd1 vssd1 vccd1 vccd1 _06521_ sky130_fd_sc_hd__o21ai_1
XFILLER_147_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14427_ clknet_leaf_45_clk _01132_ net1146 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_129_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08038__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11639_ _05820_ _05853_ _05862_ _05818_ _05819_ vssd1 vssd1 vccd1 vccd1 _05863_ sky130_fd_sc_hd__o221a_1
XFILLER_30_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14358_ clknet_leaf_140_clk _01063_ net1093 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_128_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06922__X _01758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08850__A _02264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_3_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold706 datapath.rf.registers\[8\]\[9\] vssd1 vssd1 vccd1 vccd1 net2054 sky130_fd_sc_hd__dlygate4sd3_1
Xhold717 datapath.rf.registers\[23\]\[13\] vssd1 vssd1 vccd1 vccd1 net2065 sky130_fd_sc_hd__dlygate4sd3_1
X_13309_ clknet_leaf_144_clk _00119_ net1085 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold728 datapath.rf.registers\[2\]\[27\] vssd1 vssd1 vccd1 vccd1 net2076 sky130_fd_sc_hd__dlygate4sd3_1
Xhold739 datapath.rf.registers\[5\]\[13\] vssd1 vssd1 vccd1 vccd1 net2087 sky130_fd_sc_hd__dlygate4sd3_1
X_14289_ clknet_leaf_66_clk _00994_ net1236 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_143_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08210__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08850_ _02264_ net444 vssd1 vssd1 vccd1 vccd1 _03686_ sky130_fd_sc_hd__nand2_1
XFILLER_69_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07801_ _02613_ _02635_ vssd1 vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__nor2_1
X_08781_ net566 _03615_ vssd1 vssd1 vccd1 vccd1 _03617_ sky130_fd_sc_hd__nor2_1
XANTENNA__11648__A1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07732_ datapath.rf.registers\[0\]\[16\] net866 _02557_ _02566_ vssd1 vssd1 vccd1
+ vccd1 _02568_ sky130_fd_sc_hd__o22ai_4
XANTENNA__12845__A0 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07663_ datapath.rf.registers\[13\]\[17\] net984 net917 vssd1 vssd1 vccd1 vccd1 _02499_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10320__A1 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09402_ _03673_ _04237_ _04236_ _04234_ vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__a211o_1
X_06614_ mmio.memload_or_instruction\[18\] net1048 vssd1 vssd1 vccd1 vccd1 _01453_
+ sky130_fd_sc_hd__and2_2
XANTENNA__10871__A2 _04084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07594_ datapath.rf.registers\[6\]\[19\] net681 net666 datapath.rf.registers\[15\]\[19\]
+ _02429_ vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__a221o_1
XFILLER_34_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09333_ net319 _03941_ _04168_ net322 vssd1 vssd1 vccd1 vccd1 _04169_ sky130_fd_sc_hd__a211o_1
XANTENNA__08277__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_126_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_126_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13142__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07485__D1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09264_ _02364_ net553 net549 vssd1 vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__or3_1
XANTENNA__11820__B2 _01503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08215_ _03048_ _03049_ _03050_ vssd1 vssd1 vccd1 vccd1 _03051_ sky130_fd_sc_hd__or3_1
XANTENNA__08463__C net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09195_ net367 _03955_ _04030_ vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__o21a_1
XANTENNA__12981__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1247_A net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08146_ net614 _02981_ vssd1 vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__or2_1
XFILLER_107_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08077_ datapath.rf.registers\[0\]\[9\] net869 _02911_ vssd1 vssd1 vccd1 vccd1 _02913_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_106_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1035_X net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07028_ datapath.rf.registers\[18\]\[30\] net791 _01861_ _01862_ _01863_ vssd1 vssd1
+ vccd1 vccd1 _01864_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout495_X net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout874_A _01723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold11 keypad.debounce.debounce\[6\] vssd1 vssd1 vccd1 vccd1 net1359 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 keypad.debounce.debounce\[11\] vssd1 vssd1 vccd1 vccd1 net1370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 screen.controlBus\[8\] vssd1 vssd1 vccd1 vccd1 net1381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 screen.controlBus\[28\] vssd1 vssd1 vccd1 vccd1 net1392 sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ net344 _03814_ vssd1 vssd1 vccd1 vccd1 _03815_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout662_X net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold55 net63 vssd1 vssd1 vccd1 vccd1 net1403 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold66 net55 vssd1 vssd1 vccd1 vccd1 net1414 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 net95 vssd1 vssd1 vccd1 vccd1 net1425 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 mmio.memload_or_instruction\[22\] vssd1 vssd1 vccd1 vccd1 net1436 sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ _05840_ _06032_ _06034_ net1001 vssd1 vssd1 vccd1 vccd1 _06035_ sky130_fd_sc_hd__o31a_1
XFILLER_91_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold99 screen.controlBus\[24\] vssd1 vssd1 vccd1 vccd1 net1447 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12300__A2 _06254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10941_ net902 _05680_ vssd1 vssd1 vccd1 vccd1 _05681_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_67_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout927_X net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13660_ clknet_leaf_10_clk _00470_ net1073 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10872_ datapath.mulitply_result\[20\] net615 net652 vssd1 vssd1 vccd1 vccd1 _05622_
+ sky130_fd_sc_hd__o21a_1
X_12611_ _06451_ _06455_ vssd1 vssd1 vccd1 vccd1 _06456_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_117_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_117_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13591_ clknet_leaf_130_clk _00401_ net1114 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_25_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13052__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08654__B _02091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10075__B1 _01702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12542_ _06396_ _06397_ _06395_ vssd1 vssd1 vccd1 vccd1 _06399_ sky130_fd_sc_hd__o21ai_1
XFILLER_12_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12473_ net164 _05994_ net126 screen.register.currentXbus\[29\] vssd1 vssd1 vccd1
+ vccd1 _00875_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12891__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14212_ clknet_leaf_48_clk datapath.multiplication_module.multiplicand_i_n\[23\]
+ net1177 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09766__A _04118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11424_ net252 net2359 net515 vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__mux2_1
XFILLER_6_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_8 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14143_ clknet_leaf_149_clk _00900_ net1059 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11355_ net263 net2486 net521 vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__mux2_1
XANTENNA__08440__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06902__B net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11300__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10306_ _04581_ _05141_ _05140_ net227 vssd1 vssd1 vccd1 vccd1 _05142_ sky130_fd_sc_hd__o211a_1
XANTENNA__07794__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14074_ clknet_leaf_122_clk _00841_ net1214 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_98_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11286_ net262 net2429 net525 vssd1 vssd1 vccd1 vccd1 _00334_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13025_ net1543 net175 net392 vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__mux2_1
X_10237_ _04919_ _05052_ _05061_ _05072_ vssd1 vssd1 vccd1 vccd1 _05073_ sky130_fd_sc_hd__or4b_4
XFILLER_121_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1020 net1021 vssd1 vssd1 vccd1 vccd1 net1020 sky130_fd_sc_hd__buf_4
XANTENNA__09753__B1_N net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1031 net1032 vssd1 vssd1 vccd1 vccd1 net1031 sky130_fd_sc_hd__buf_2
Xfanout1042 _03730_ vssd1 vssd1 vccd1 vccd1 net1042 sky130_fd_sc_hd__buf_2
XFILLER_121_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10168_ datapath.PC\[16\] _03741_ vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__and2_1
Xfanout1053 net1058 vssd1 vssd1 vccd1 vccd1 net1053 sky130_fd_sc_hd__buf_2
Xfanout1064 net1066 vssd1 vssd1 vccd1 vccd1 net1064 sky130_fd_sc_hd__clkbuf_4
Xfanout1075 net1121 vssd1 vssd1 vccd1 vccd1 net1075 sky130_fd_sc_hd__clkbuf_2
Xfanout1086 net1092 vssd1 vssd1 vccd1 vccd1 net1086 sky130_fd_sc_hd__clkbuf_4
Xfanout1097 net1101 vssd1 vssd1 vccd1 vccd1 net1097 sky130_fd_sc_hd__clkbuf_4
X_10099_ net468 _03830_ _03864_ _04934_ vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__a31o_1
XFILLER_81_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07452__C net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13927_ clknet_leaf_95_clk _00705_ net1226 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10302__A1 _01702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13858_ clknet_leaf_72_clk _00662_ net1243 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__06917__X _01753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08259__B1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12809_ net2300 net264 net493 vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_108_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_108_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13789_ clknet_leaf_73_clk _00598_ net1243 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08000_ datapath.rf.registers\[21\]\[10\] net947 net925 vssd1 vssd1 vccd1 vccd1 _02836_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12358__A2 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold503 datapath.multiplication_module.multiplicand_i\[4\] vssd1 vssd1 vccd1 vccd1
+ net1851 sky130_fd_sc_hd__dlygate4sd3_1
Xhold514 datapath.rf.registers\[31\]\[17\] vssd1 vssd1 vccd1 vccd1 net1862 sky130_fd_sc_hd__dlygate4sd3_1
Xhold525 datapath.rf.registers\[8\]\[28\] vssd1 vssd1 vccd1 vccd1 net1873 sky130_fd_sc_hd__dlygate4sd3_1
Xhold536 datapath.rf.registers\[26\]\[2\] vssd1 vssd1 vccd1 vccd1 net1884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold547 datapath.rf.registers\[31\]\[23\] vssd1 vssd1 vccd1 vccd1 net1895 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11210__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07785__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold558 datapath.rf.registers\[10\]\[28\] vssd1 vssd1 vccd1 vccd1 net1906 sky130_fd_sc_hd__dlygate4sd3_1
X_09951_ _04784_ _04785_ _04779_ vssd1 vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__a21bo_1
Xhold569 datapath.rf.registers\[21\]\[10\] vssd1 vssd1 vccd1 vccd1 net1917 sky130_fd_sc_hd__dlygate4sd3_1
X_08902_ datapath.PC\[11\] _03737_ vssd1 vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__or2_1
X_09882_ datapath.PC\[28\] net595 vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__or2_1
XANTENNA__07537__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08833_ _01611_ _01614_ _01618_ vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__or3b_2
Xhold1203 screen.register.currentXbus\[0\] vssd1 vssd1 vccd1 vccd1 net2551 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1214 datapath.rf.registers\[20\]\[29\] vssd1 vssd1 vccd1 vccd1 net2562 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1225 datapath.rf.registers\[31\]\[14\] vssd1 vssd1 vccd1 vccd1 net2573 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13137__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1236 datapath.mulitply_result\[20\] vssd1 vssd1 vccd1 vccd1 net2584 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1247 datapath.mulitply_result\[28\] vssd1 vssd1 vccd1 vccd1 net2595 sky130_fd_sc_hd__dlygate4sd3_1
X_08764_ _01601_ _01604_ vssd1 vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__nand2b_1
Xhold1258 datapath.rf.registers\[3\]\[14\] vssd1 vssd1 vccd1 vccd1 net2606 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1269 datapath.PC\[9\] vssd1 vssd1 vccd1 vccd1 net2617 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_54_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07715_ datapath.rf.registers\[22\]\[16\] net821 net819 datapath.rf.registers\[5\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__a22o_1
XANTENNA__12976__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07362__C net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08695_ _02805_ _02825_ vssd1 vssd1 vccd1 vccd1 _03531_ sky130_fd_sc_hd__nand2_2
XFILLER_38_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12829__X _06552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1197_A net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07646_ datapath.rf.registers\[28\]\[18\] net750 net668 datapath.rf.registers\[21\]\[18\]
+ _02481_ vssd1 vssd1 vccd1 vccd1 _02482_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_146_Right_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10844__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06827__X _01663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07577_ datapath.rf.registers\[20\]\[19\] net840 _02393_ _02394_ _02396_ vssd1 vssd1
+ vccd1 vccd1 _02413_ sky130_fd_sc_hd__a2111o_1
XFILLER_15_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09316_ _02523_ net561 net441 vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09247_ net608 _04058_ _04082_ net556 vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout410_X net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout508_X net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09178_ _03500_ net627 net624 _03501_ net644 vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout991_A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08129_ datapath.rf.registers\[26\]\[8\] net780 net677 datapath.rf.registers\[29\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__a22o_1
XANTENNA__08422__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11120__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07776__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08973__A1 _03204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11140_ _05517_ _05717_ vssd1 vssd1 vccd1 vccd1 _05718_ sky130_fd_sc_hd__nand2_1
Xoutput45 net45 vssd1 vssd1 vccd1 vccd1 ADR_O[14] sky130_fd_sc_hd__buf_2
XANTENNA_fanout877_X net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput56 net56 vssd1 vssd1 vccd1 vccd1 ADR_O[24] sky130_fd_sc_hd__buf_2
XFILLER_150_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput67 net67 vssd1 vssd1 vccd1 vccd1 ADR_O[5] sky130_fd_sc_hd__buf_2
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 DAT_O[14] sky130_fd_sc_hd__buf_2
X_11071_ _05690_ _05712_ vssd1 vssd1 vccd1 vccd1 _05713_ sky130_fd_sc_hd__or2_1
Xoutput89 net89 vssd1 vssd1 vccd1 vccd1 DAT_O[24] sky130_fd_sc_hd__buf_2
X_10022_ _04749_ _04750_ vssd1 vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__nor2_1
XFILLER_130_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13047__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07553__B net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input16_A DAT_I[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11973_ net1007 _05764_ vssd1 vssd1 vccd1 vccd1 _06018_ sky130_fd_sc_hd__nor2_2
XANTENNA__12886__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07272__C net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12285__B2 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09150__A1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13712_ clknet_leaf_22_clk _00522_ net1156 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10924_ datapath.PC\[27\] _05654_ datapath.PC\[28\] vssd1 vssd1 vccd1 vccd1 _05666_
+ sky130_fd_sc_hd__a21oi_1
X_14692_ clknet_leaf_23_clk _01397_ net1156 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07161__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Right_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07700__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10855_ _05606_ vssd1 vssd1 vccd1 vccd1 _05607_ sky130_fd_sc_hd__inv_2
X_13643_ clknet_leaf_54_clk _00453_ net1179 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13574_ clknet_leaf_29_clk _00384_ net1133 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10786_ datapath.PC\[8\] _05542_ vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__and2_1
XANTENNA__11796__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12525_ net2542 net504 net500 _06384_ vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_30_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12456_ net164 _05960_ net126 screen.register.currentXbus\[12\] vssd1 vssd1 vccd1
+ vccd1 _00858_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_97_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06913__A net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11407_ net2445 net174 net412 vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__mux2_1
X_12387_ _05944_ net159 vssd1 vssd1 vccd1 vccd1 _06341_ sky130_fd_sc_hd__nor2_1
XANTENNA__10435__A _05211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11030__S net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14126_ clknet_leaf_138_clk _00883_ net1100 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07767__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08964__A1 _02804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11338_ net2393 net181 net415 vssd1 vssd1 vccd1 vccd1 _00383_ sky130_fd_sc_hd__mux2_1
XFILLER_98_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10771__A1 _01441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14057_ clknet_leaf_95_clk _00824_ net1216 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11269_ net179 net1933 net421 vssd1 vssd1 vccd1 vccd1 _00318_ sky130_fd_sc_hd__mux2_1
XANTENNA__07519__A2 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13008_ net2053 net254 net390 vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08559__B net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09677__C1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07099__A2_N net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07500_ datapath.rf.registers\[9\]\[20\] net982 net943 vssd1 vssd1 vccd1 vccd1 _02336_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09141__A1 _03604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08480_ datapath.rf.registers\[12\]\[1\] net828 _01768_ datapath.rf.registers\[28\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03316_ sky130_fd_sc_hd__a22o_1
XFILLER_63_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_914 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07152__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09023__X _03859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07431_ datapath.rf.registers\[30\]\[22\] net758 net750 datapath.rf.registers\[28\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__a22o_1
XANTENNA__11205__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07362_ datapath.rf.registers\[6\]\[23\] net954 net932 vssd1 vssd1 vccd1 vccd1 _02198_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_44_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09101_ net344 _03792_ vssd1 vssd1 vccd1 vccd1 _03937_ sky130_fd_sc_hd__nor2_1
X_07293_ datapath.rf.registers\[12\]\[25\] net756 net696 datapath.rf.registers\[8\]\[25\]
+ _02128_ vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__a221o_1
X_09032_ net633 _03867_ vssd1 vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__nand2_1
Xhold300 datapath.rf.registers\[6\]\[30\] vssd1 vssd1 vccd1 vccd1 net1648 sky130_fd_sc_hd__dlygate4sd3_1
Xhold311 datapath.rf.registers\[5\]\[7\] vssd1 vssd1 vccd1 vccd1 net1659 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout203_A _05641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold322 datapath.rf.registers\[6\]\[2\] vssd1 vssd1 vccd1 vccd1 net1670 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09693__X _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08955__A1 _02523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold333 datapath.rf.registers\[14\]\[17\] vssd1 vssd1 vccd1 vccd1 net1681 sky130_fd_sc_hd__dlygate4sd3_1
Xhold344 datapath.rf.registers\[14\]\[11\] vssd1 vssd1 vccd1 vccd1 net1692 sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 datapath.rf.registers\[7\]\[24\] vssd1 vssd1 vccd1 vccd1 net1703 sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 datapath.rf.registers\[4\]\[29\] vssd1 vssd1 vccd1 vccd1 net1714 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07357__C net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10064__B net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold377 datapath.rf.registers\[4\]\[21\] vssd1 vssd1 vccd1 vccd1 net1725 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold388 datapath.rf.registers\[22\]\[2\] vssd1 vssd1 vccd1 vccd1 net1736 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout802 _01769_ vssd1 vssd1 vccd1 vccd1 net802 sky130_fd_sc_hd__buf_6
Xhold399 datapath.rf.registers\[5\]\[24\] vssd1 vssd1 vccd1 vccd1 net1747 sky130_fd_sc_hd__dlygate4sd3_1
X_09934_ net1268 _03077_ vssd1 vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__or2_1
Xfanout813 net814 vssd1 vssd1 vccd1 vccd1 net813 sky130_fd_sc_hd__buf_4
Xfanout824 net825 vssd1 vssd1 vccd1 vccd1 net824 sky130_fd_sc_hd__buf_4
Xfanout835 _01746_ vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout846 _01737_ vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07654__A _02467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input8_A DAT_I[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout857 net859 vssd1 vssd1 vccd1 vccd1 net857 sky130_fd_sc_hd__clkbuf_4
X_09865_ _03128_ _03426_ _03561_ _03563_ vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__a211o_1
Xhold1000 datapath.rf.registers\[20\]\[17\] vssd1 vssd1 vccd1 vccd1 net2348 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout868 net869 vssd1 vssd1 vccd1 vccd1 net868 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout572_A net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1011 datapath.rf.registers\[24\]\[14\] vssd1 vssd1 vccd1 vccd1 net2359 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout879 net881 vssd1 vssd1 vccd1 vccd1 net879 sky130_fd_sc_hd__clkbuf_8
XFILLER_86_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1022 datapath.rf.registers\[15\]\[21\] vssd1 vssd1 vccd1 vccd1 net2370 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08183__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08816_ _01666_ _03358_ _03643_ vssd1 vssd1 vccd1 vccd1 _03652_ sky130_fd_sc_hd__mux2_1
Xhold1033 datapath.rf.registers\[18\]\[2\] vssd1 vssd1 vccd1 vccd1 net2381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1044 datapath.rf.registers\[29\]\[25\] vssd1 vssd1 vccd1 vccd1 net2392 sky130_fd_sc_hd__dlygate4sd3_1
X_09796_ net380 _04256_ vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__nor2_1
XANTENNA__07391__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1055 screen.register.currentYbus\[23\] vssd1 vssd1 vccd1 vccd1 net2403 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1066 screen.counter.currentCt\[16\] vssd1 vssd1 vccd1 vccd1 net2414 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1077 mmio.memload_or_instruction\[17\] vssd1 vssd1 vccd1 vccd1 net2425 sky130_fd_sc_hd__dlygate4sd3_1
X_08747_ _03507_ _03508_ _03582_ vssd1 vssd1 vccd1 vccd1 _03583_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_90_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1088 datapath.rf.registers\[31\]\[20\] vssd1 vssd1 vccd1 vccd1 net2436 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1099 datapath.rf.registers\[17\]\[22\] vssd1 vssd1 vccd1 vccd1 net2447 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout837_A _01743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08678_ _02523_ _02543_ vssd1 vssd1 vccd1 vccd1 _03514_ sky130_fd_sc_hd__nand2_1
XANTENNA__10817__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08485__A net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14104__RESET_B net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07629_ _02464_ _02444_ net866 _02460_ vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__and4b_1
XANTENNA_fanout625_X net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11115__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10640_ _05431_ _05458_ keypad.alpha vssd1 vssd1 vccd1 vccd1 _05460_ sky130_fd_sc_hd__a21oi_1
XFILLER_42_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08772__X _03608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10571_ _02804_ _02856_ _02912_ _02960_ vssd1 vssd1 vccd1 vccd1 _05394_ sky130_fd_sc_hd__or4_1
XFILLER_155_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12310_ net228 _05589_ _06287_ net635 vssd1 vssd1 vccd1 vccd1 _06288_ sky130_fd_sc_hd__a211o_1
X_13290_ clknet_leaf_59_clk _00100_ net1168 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06733__A _01571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12241_ screen.counter.currentCt\[17\] screen.counter.currentCt\[18\] _06233_ vssd1
+ vssd1 vccd1 vccd1 _06237_ sky130_fd_sc_hd__and3_1
XFILLER_135_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07749__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12172_ _05802_ _06157_ _06170_ vssd1 vssd1 vccd1 vccd1 _06194_ sky130_fd_sc_hd__and3_1
XANTENNA__07267__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11123_ net245 net2217 net426 vssd1 vssd1 vccd1 vccd1 _00178_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_92_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_43_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11054_ net243 net2234 net430 vssd1 vssd1 vccd1 vccd1 _00114_ sky130_fd_sc_hd__mux2_1
XFILLER_107_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11702__B1 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09371__A1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08174__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10005_ _04840_ _04839_ vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__and2b_1
XANTENNA__09371__B2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07921__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_58_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10269__B1 net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_101_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11956_ _05784_ _05786_ net996 _05795_ vssd1 vssd1 vccd1 vccd1 _06002_ sky130_fd_sc_hd__or4b_1
XANTENNA__08395__A _03204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09674__A2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10907_ datapath.mulitply_result\[25\] net597 net617 vssd1 vssd1 vccd1 vccd1 _05652_
+ sky130_fd_sc_hd__a21o_1
X_11887_ net2635 net162 vssd1 vssd1 vccd1 vccd1 _05955_ sky130_fd_sc_hd__nand2_1
X_14675_ clknet_leaf_34_clk _01380_ net1127 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11025__S net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13626_ clknet_leaf_14_clk _00436_ net1078 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10838_ net247 net2028 net542 vssd1 vssd1 vccd1 vccd1 _00017_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_116_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13557_ clknet_leaf_19_clk _00367_ net1116 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10769_ net901 _04454_ _05533_ vssd1 vssd1 vccd1 vccd1 _05534_ sky130_fd_sc_hd__o21a_1
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07988__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12508_ net173 net1628 net507 vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__mux2_1
X_13488_ clknet_leaf_25_clk _00298_ net1158 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08561__C _01825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12439_ _05996_ net156 vssd1 vssd1 vccd1 vccd1 _06367_ sky130_fd_sc_hd__nor2_1
XANTENNA__07458__B net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08937__A1 _01981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14109_ clknet_leaf_111_clk _00875_ net1202 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_07980_ datapath.rf.registers\[19\]\[11\] net732 net685 datapath.rf.registers\[27\]\[11\]
+ _02815_ vssd1 vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__a221o_1
XFILLER_141_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06931_ datapath.rf.registers\[13\]\[31\] net810 net807 datapath.rf.registers\[27\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__a22o_1
XANTENNA__08165__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09650_ _03667_ _04480_ _04481_ _04485_ vssd1 vssd1 vccd1 vccd1 _04486_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_143_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06862_ datapath.ru.latched_instruction\[23\] net990 _01665_ datapath.ru.latched_instruction\[21\]
+ _01668_ vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__a221o_1
XFILLER_27_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08601_ _03431_ _03435_ vssd1 vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__nand2_1
XFILLER_67_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07912__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09581_ _04341_ _04342_ net457 vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__o21a_1
X_06793_ _01451_ net1003 net1019 net1026 datapath.ru.latched_instruction\[17\] vssd1
+ vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__a32oi_4
XFILLER_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08532_ datapath.rf.registers\[16\]\[0\] net862 _03366_ _03367_ vssd1 vssd1 vccd1
+ vccd1 _03368_ sky130_fd_sc_hd__a211o_1
XFILLER_24_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08873__A0 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08463_ datapath.rf.registers\[29\]\[1\] net979 net918 vssd1 vssd1 vccd1 vccd1 _03299_
+ sky130_fd_sc_hd__and3_1
XFILLER_50_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout153_A net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07414_ datapath.rf.registers\[24\]\[22\] net856 net790 datapath.rf.registers\[18\]\[22\]
+ _02244_ vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__a221o_1
X_08394_ _03204_ _03228_ vssd1 vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__or2_1
XANTENNA__10059__B net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07345_ datapath.rf.registers\[17\]\[24\] net746 net723 datapath.rf.registers\[18\]\[24\]
+ _02180_ vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__a221o_1
XANTENNA__13150__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout418_A _05722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_30_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07979__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07276_ datapath.rf.registers\[30\]\[25\] net834 _02100_ _02106_ _02109_ vssd1 vssd1
+ vccd1 vccd1 _02112_ sky130_fd_sc_hd__a2111o_1
XFILLER_12_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09015_ _03692_ _03703_ net342 vssd1 vssd1 vccd1 vccd1 _03851_ sky130_fd_sc_hd__mux2_1
XFILLER_152_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06703__D datapath.ru.latched_instruction\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold130 net81 vssd1 vssd1 vccd1 vccd1 net1478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 mmio.memload_or_instruction\[3\] vssd1 vssd1 vccd1 vccd1 net1489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 net82 vssd1 vssd1 vccd1 vccd1 net1500 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 screen.counter.currentCt\[17\] vssd1 vssd1 vccd1 vccd1 net1511 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout787_A net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold174 mmio.wishbone.curr_state\[2\] vssd1 vssd1 vccd1 vccd1 net1522 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold185 datapath.multiplication_module.multiplicand_i\[16\] vssd1 vssd1 vccd1 vccd1
+ net1533 sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 datapath.multiplication_module.multiplicand_i\[18\] vssd1 vssd1 vccd1 vccd1
+ net1544 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout610 _01782_ vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__clkbuf_4
Xfanout621 net622 vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09917_ net1266 _04751_ vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__xor2_1
Xfanout632 net633 vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout643 net646 vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__buf_2
Xfanout654 net655 vssd1 vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout575_X net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08199__B net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_97_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_97_clk sky130_fd_sc_hd__clkbuf_8
Xfanout665 net667 vssd1 vssd1 vccd1 vccd1 net665 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08156__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout676 net678 vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_13_Left_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout687 net690 vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09848_ _03477_ _03478_ _03611_ _04683_ vssd1 vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__a31o_1
Xfanout698 net701 vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07903__A2 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout742_X net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09779_ net575 _04613_ _04614_ _04612_ vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__a22o_1
X_11810_ _01523_ net1015 net313 net333 datapath.ru.latched_instruction\[16\] vssd1
+ vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_1_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ net194 net2242 net494 vssd1 vssd1 vccd1 vccd1 _01043_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07116__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06728__A net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11741_ net1428 net147 net142 _03357_ vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__a22o_1
XFILLER_53_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14460_ clknet_leaf_10_clk _01165_ net1081 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11672_ _05270_ net154 net150 net1408 vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__a22o_1
XFILLER_53_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10623_ net121 net123 net124 net122 vssd1 vssd1 vccd1 vccd1 _05443_ sky130_fd_sc_hd__or4b_4
X_13411_ clknet_leaf_120_clk _00221_ net1193 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_14391_ clknet_leaf_131_clk _01096_ net1205 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13060__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_21_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08662__B _02240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13342_ clknet_leaf_1_clk _00152_ net1063 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10554_ net37 _05380_ vssd1 vssd1 vccd1 vccd1 _05381_ sky130_fd_sc_hd__and2b_1
XFILLER_154_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13273_ clknet_leaf_30_clk _00083_ net1131 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10485_ _05307_ _05310_ _05313_ vssd1 vssd1 vccd1 vccd1 _05315_ sky130_fd_sc_hd__nand3_4
XFILLER_142_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11518__A3 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12224_ screen.counter.currentCt\[11\] _06223_ screen.counter.currentCt\[12\] vssd1
+ vssd1 vccd1 vccd1 _06226_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10726__A1 _02750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_90_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09592__A1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12155_ _06160_ net567 _06179_ vssd1 vssd1 vccd1 vccd1 _06184_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_9_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06910__B net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11106_ _05695_ _05715_ vssd1 vssd1 vccd1 vccd1 _05716_ sky130_fd_sc_hd__nand2_4
XFILLER_1_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12086_ screen.register.currentYbus\[14\] _05776_ net997 screen.register.currentXbus\[22\]
+ vssd1 vssd1 vccd1 vccd1 _06125_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_88_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_88_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08147__A2 _02980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11037_ _05695_ _05710_ vssd1 vssd1 vccd1 vccd1 _05711_ sky130_fd_sc_hd__nand2_1
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14026__RESET_B net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07581__X _02417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10859__S net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07107__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12988_ net192 net2435 net478 vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__mux2_1
XANTENNA__08855__A0 _02523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11939_ _02045_ screen.counter.ack vssd1 vssd1 vccd1 vccd1 _05990_ sky130_fd_sc_hd__or2_1
XFILLER_33_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14658_ clknet_leaf_151_clk _01363_ net1052 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13609_ clknet_leaf_21_clk _00419_ net1163 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14589_ clknet_leaf_147_clk _01294_ net1064 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_12_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08572__B net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07130_ datapath.rf.registers\[12\]\[28\] net828 net797 datapath.rf.registers\[29\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__a22o_1
Xteam_04_1307 vssd1 vssd1 vccd1 vccd1 team_04_1307/HI gpio_oeb[16] sky130_fd_sc_hd__conb_1
Xteam_04_1318 vssd1 vssd1 vccd1 vccd1 team_04_1318/HI gpio_out[22] sky130_fd_sc_hd__conb_1
Xteam_04_1329 vssd1 vssd1 vccd1 vccd1 team_04_1329/HI gpio_out[33] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_136_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07061_ datapath.rf.registers\[1\]\[30\] net764 net716 datapath.rf.registers\[4\]\[30\]
+ _01896_ vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__a221o_1
XANTENNA__06633__A2 _01466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13551__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08386__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11390__A1 _05582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07594__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07963_ datapath.rf.registers\[21\]\[11\] net816 _02781_ _02782_ _02783_ vssd1 vssd1
+ vccd1 vccd1 _02799_ sky130_fd_sc_hd__a2111o_1
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_79_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08138__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09702_ _04496_ _04516_ _04534_ _04536_ vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__and4_1
X_06914_ datapath.rf.registers\[14\]\[31\] net829 net827 datapath.rf.registers\[12\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__a22o_1
X_07894_ datapath.rf.registers\[25\]\[12\] net975 net943 vssd1 vssd1 vccd1 vccd1 _02730_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08587__X _03423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07346__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_52_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06845_ _01414_ net993 _01645_ _01670_ vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__a31o_1
X_09633_ _03541_ net628 _04468_ net645 vssd1 vssd1 vccd1 vccd1 _04469_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout270_A _05564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout368_A net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13145__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09564_ net606 _04399_ vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__or2_1
X_06776_ net1005 net1021 _01612_ net1030 datapath.ru.latched_instruction\[12\] vssd1
+ vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__a32o_2
XFILLER_130_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08466__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08515_ datapath.rf.registers\[14\]\[1\] net777 _03348_ _03349_ _03350_ vssd1 vssd1
+ vccd1 vccd1 _03351_ sky130_fd_sc_hd__a2111o_1
XFILLER_70_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13749__RESET_B net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12984__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09495_ _03544_ net626 net625 _03553_ net643 vssd1 vssd1 vccd1 vccd1 _04331_ sky130_fd_sc_hd__a221oi_1
XFILLER_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout535_A net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08310__A2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08446_ _03279_ _03280_ _03281_ vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_156_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08377_ datapath.rf.registers\[17\]\[3\] net748 net732 datapath.rf.registers\[19\]\[3\]
+ _03212_ vssd1 vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout702_A net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07328_ datapath.rf.registers\[22\]\[24\] net822 _02149_ _02150_ _02151_ vssd1 vssd1
+ vccd1 vccd1 _02164_ sky130_fd_sc_hd__a2111o_1
XFILLER_139_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07259_ datapath.rf.registers\[31\]\[25\] net978 net915 vssd1 vssd1 vccd1 vccd1 _02095_
+ sky130_fd_sc_hd__and3_1
X_10270_ _05097_ _05105_ datapath.PC\[13\] net1294 vssd1 vssd1 vccd1 vccd1 _05106_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_136_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10708__A1 _02725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout692_X net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14537__RESET_B net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08377__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07585__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout440 _03761_ vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout957_X net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14190__RESET_B net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08129__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout451 _03678_ vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__buf_2
Xfanout462 _03651_ vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__clkbuf_2
X_13960_ clknet_leaf_107_clk _00738_ net1221 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_59_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout473 _06561_ vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__buf_4
XANTENNA__07337__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout484 net485 vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09877__A2 _04710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout495 _06550_ vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__clkbuf_4
XFILLER_101_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12911_ net2312 net249 net483 vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__mux2_1
XFILLER_74_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13891_ clknet_leaf_43_clk keypad.decode.button_n\[2\] net1152 vssd1 vssd1 vccd1
+ vccd1 button\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13055__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12842_ net264 net2525 net489 vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12894__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12773_ net274 net2320 net496 vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__mux2_1
XFILLER_54_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08301__A2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14512_ clknet_leaf_25_clk _01217_ net1159 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11724_ net10 net1035 net1025 net2425 vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__a22o_1
XANTENNA__09769__A _03978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08673__A _02419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11655_ button\[1\] _05874_ vssd1 vssd1 vccd1 vccd1 _05877_ sky130_fd_sc_hd__and2_1
X_14443_ clknet_leaf_56_clk _01148_ net1160 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11303__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06905__B net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10606_ screen.register.currentYbus\[18\] _05422_ _05423_ _05426_ vssd1 vssd1 vccd1
+ vccd1 _05427_ sky130_fd_sc_hd__or4_1
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11586_ net1273 net1270 screen.counter.ct\[16\] net1274 vssd1 vssd1 vccd1 vccd1 _05810_
+ sky130_fd_sc_hd__or4b_1
XANTENNA__08960__X _03796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14374_ clknet_leaf_23_clk _01079_ net1154 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_13325_ clknet_leaf_126_clk _00135_ net1205 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10537_ net180 net189 _05271_ _05365_ vssd1 vssd1 vccd1 vccd1 _05366_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_118_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10468_ screen.counter.ct\[11\] net1275 net1273 net1274 vssd1 vssd1 vccd1 vccd1 _05298_
+ sky130_fd_sc_hd__or4_1
X_13256_ clknet_leaf_66_clk _00066_ net1236 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09565__A1 _03149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12207_ screen.counter.currentCt\[6\] _06214_ vssd1 vssd1 vccd1 vccd1 _06215_ sky130_fd_sc_hd__and2_1
X_13187_ net2624 vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__clkbuf_1
X_10399_ _01605_ net642 _03603_ vssd1 vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10175__A2 _01701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12138_ screen.counter.ct\[1\] net567 _06173_ net601 vssd1 vssd1 vccd1 vccd1 _00736_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10162__B _04177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07455__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09317__A1 _02418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12069_ screen.register.currentYbus\[5\] _05778_ _05786_ screen.register.currentYbus\[29\]
+ vssd1 vssd1 vccd1 vccd1 _06109_ sky130_fd_sc_hd__a22o_1
XFILLER_84_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_1_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06630_ mmio.memload_or_instruction\[19\] net1048 vssd1 vssd1 vccd1 vccd1 _01469_
+ sky130_fd_sc_hd__and2_1
XANTENNA__08540__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08828__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08300_ datapath.rf.registers\[21\]\[4\] net815 _03129_ _03135_ vssd1 vssd1 vccd1
+ vccd1 _03136_ sky130_fd_sc_hd__a211o_1
X_09280_ net317 _04113_ _04115_ _04110_ _04112_ vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_138_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08231_ datapath.rf.registers\[28\]\[6\] net750 net675 datapath.rf.registers\[29\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03067_ sky130_fd_sc_hd__a22o_1
XANTENNA__06854__A2 _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11213__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08162_ datapath.rf.registers\[2\]\[7\] net889 net818 datapath.rf.registers\[7\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02998_ sky130_fd_sc_hd__a22o_1
XANTENNA__09253__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07113_ datapath.rf.registers\[7\]\[29\] net671 _01948_ net787 vssd1 vssd1 vccd1
+ vccd1 _01949_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_151_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06606__A2 _01441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08093_ datapath.rf.registers\[8\]\[9\] net696 net666 datapath.rf.registers\[15\]\[9\]
+ _02928_ vssd1 vssd1 vccd1 vccd1 _02929_ sky130_fd_sc_hd__a221o_1
XFILLER_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload50 clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 clkload50/Y sky130_fd_sc_hd__inv_6
X_07044_ datapath.rf.registers\[10\]\[30\] net881 net812 datapath.rf.registers\[13\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__a22o_1
XANTENNA__09005__B1 _01934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload61 clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 clkload61/Y sky130_fd_sc_hd__clkinv_4
Xclkload72 clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 clkload72/Y sky130_fd_sc_hd__inv_12
XFILLER_115_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload83 clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 clkload83/Y sky130_fd_sc_hd__clkinv_2
XFILLER_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload94 clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 clkload94/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__08359__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07365__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12979__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08995_ _03593_ _03828_ vssd1 vssd1 vccd1 vccd1 _03831_ sky130_fd_sc_hd__nand2_1
XFILLER_141_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout485_A _06554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07946_ datapath.rf.registers\[5\]\[11\] net947 net934 vssd1 vssd1 vccd1 vccd1 _02782_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07319__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07877_ datapath.rf.registers\[3\]\[13\] net771 net703 datapath.rf.registers\[9\]\[13\]
+ _02712_ vssd1 vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__a221o_1
XFILLER_29_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08531__A2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09616_ net607 _04430_ vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__or2_1
X_06828_ _01663_ vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__inv_2
XFILLER_141_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06759_ _01503_ net1005 net1021 net1031 datapath.ru.latched_instruction\[26\] vssd1
+ vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout440_X net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09547_ net377 _04374_ _04382_ net330 vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__o211ai_1
XANTENNA_fanout538_X net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout917_A _01764_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08764__Y _03600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11912__A _02487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09478_ net326 _04107_ _04309_ _04313_ vssd1 vssd1 vccd1 vccd1 _04314_ sky130_fd_sc_hd__o22a_1
X_08429_ _01637_ _01783_ _03264_ _01704_ vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__10528__A _05315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout705_X net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11123__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload0 clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clkload0/X sky130_fd_sc_hd__clkbuf_8
X_11440_ net175 net2183 net516 vssd1 vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__mux2_1
XFILLER_137_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11371_ net176 net1667 net518 vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__mux2_1
XFILLER_4_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10322_ datapath.PC\[15\] _04207_ net467 vssd1 vssd1 vccd1 vccd1 _05158_ sky130_fd_sc_hd__mux2_1
X_13110_ net250 net2280 net470 vssd1 vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__mux2_1
X_14090_ clknet_leaf_96_clk _00856_ net1226 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06741__A _01579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13041_ net262 net2314 net475 vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__mux2_1
X_10253_ _03738_ _05088_ net1040 vssd1 vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__a21oi_1
XFILLER_152_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10263__A net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07556__B net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14300__RESET_B net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10184_ datapath.PC\[17\] _03742_ vssd1 vssd1 vccd1 vccd1 _05020_ sky130_fd_sc_hd__xnor2_1
Xfanout1202 net1203 vssd1 vssd1 vccd1 vccd1 net1202 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12889__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1213 net1262 vssd1 vssd1 vccd1 vccd1 net1213 sky130_fd_sc_hd__buf_2
XFILLER_132_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1224 net1225 vssd1 vssd1 vccd1 vccd1 net1224 sky130_fd_sc_hd__buf_2
Xfanout1235 net1238 vssd1 vssd1 vccd1 vccd1 net1235 sky130_fd_sc_hd__clkbuf_4
Xfanout1246 net1248 vssd1 vssd1 vccd1 vccd1 net1246 sky130_fd_sc_hd__clkbuf_4
Xfanout1257 net1261 vssd1 vssd1 vccd1 vccd1 net1257 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_89_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08668__A _02312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout270 _05564_ vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__clkbuf_2
Xfanout1268 datapath.PC\[6\] vssd1 vssd1 vccd1 vccd1 net1268 sky130_fd_sc_hd__buf_2
Xfanout1279 screen.counter.ct\[6\] vssd1 vssd1 vccd1 vccd1 net1279 sky130_fd_sc_hd__clkbuf_2
Xfanout281 _05554_ vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__buf_1
Xfanout292 net293 vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11699__A2_N _05885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13943_ clknet_leaf_122_clk _00721_ net1216 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08020__X _02856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10710__B _05368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08522__A2 _03357_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10865__B1 _05614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13874_ clknet_leaf_51_clk _00678_ net1182 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_35_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14178__Q datapath.mulitply_result\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12825_ net2278 net179 net493 vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__mux2_1
XFILLER_15_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07089__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12756_ net2338 net198 net404 vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__mux2_1
XANTENNA__09483__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11707_ net2 net1033 net1023 net1457 vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__o22a_1
X_12687_ _06517_ _06518_ _06519_ vssd1 vssd1 vccd1 vccd1 _06520_ sky130_fd_sc_hd__or3_1
XANTENNA__06635__B net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11033__S net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14426_ clknet_leaf_146_clk _01131_ net1088 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_11638_ _05785_ _05812_ _05859_ _05783_ _05852_ vssd1 vssd1 vccd1 vccd1 _05862_ sky130_fd_sc_hd__o221a_1
XFILLER_128_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14357_ clknet_leaf_129_clk _01062_ net1117 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_144_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11569_ _05294_ net1008 vssd1 vssd1 vccd1 vccd1 _05793_ sky130_fd_sc_hd__nor2_1
Xhold707 screen.controlBus\[2\] vssd1 vssd1 vccd1 vccd1 net2055 sky130_fd_sc_hd__dlygate4sd3_1
X_13308_ clknet_leaf_8_clk _00118_ net1072 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold718 datapath.rf.registers\[13\]\[8\] vssd1 vssd1 vccd1 vccd1 net2066 sky130_fd_sc_hd__dlygate4sd3_1
Xhold729 datapath.rf.registers\[22\]\[5\] vssd1 vssd1 vccd1 vccd1 net2077 sky130_fd_sc_hd__dlygate4sd3_1
X_14288_ clknet_leaf_58_clk _00993_ net1160 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_131_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13239_ clknet_leaf_130_clk _00049_ net1114 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07549__B1 _02384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07013__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12799__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07800_ _02613_ _02635_ vssd1 vssd1 vccd1 vccd1 _02636_ sky130_fd_sc_hd__nand2_1
XFILLER_112_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08780_ net647 net606 _03614_ vssd1 vssd1 vccd1 vccd1 _03616_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_127_Right_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07731_ datapath.rf.registers\[0\]\[16\] net866 _02557_ _02566_ vssd1 vssd1 vccd1
+ vccd1 _02567_ sky130_fd_sc_hd__o22a_4
XANTENNA__10856__A0 _04600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11208__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07662_ datapath.rf.registers\[4\]\[17\] net959 net935 vssd1 vssd1 vccd1 vccd1 _02498_
+ sky130_fd_sc_hd__and3_1
XFILLER_53_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06613_ net1290 net1281 mmio.memload_or_instruction\[17\] vssd1 vssd1 vccd1 vccd1
+ _01452_ sky130_fd_sc_hd__or3b_1
X_09401_ _04011_ _04019_ net320 vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__mux2_1
X_07593_ datapath.rf.registers\[14\]\[19\] net776 net693 datapath.rf.registers\[13\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__a22o_1
XFILLER_52_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09332_ net320 _03936_ vssd1 vssd1 vccd1 vccd1 _04168_ sky130_fd_sc_hd__nor2_1
X_09263_ net350 _03842_ _03845_ _03846_ net356 vssd1 vssd1 vccd1 vccd1 _04099_ sky130_fd_sc_hd__o311ai_1
X_08214_ datapath.rf.registers\[21\]\[6\] net815 _03037_ _03038_ _03040_ vssd1 vssd1
+ vccd1 vccd1 _03050_ sky130_fd_sc_hd__a2111o_1
X_09194_ net563 net440 _04029_ net364 vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__a211o_1
X_08145_ _01600_ _01784_ vssd1 vssd1 vccd1 vccd1 _02981_ sky130_fd_sc_hd__nor2_1
XFILLER_146_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10782__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout400_A net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07788__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07252__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08076_ datapath.rf.registers\[0\]\[9\] net869 _02911_ vssd1 vssd1 vccd1 vccd1 _02912_
+ sky130_fd_sc_hd__o21a_2
XFILLER_150_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07027_ datapath.rf.registers\[4\]\[30\] net959 net935 vssd1 vssd1 vccd1 vccd1 _01863_
+ sky130_fd_sc_hd__and3_1
XFILLER_103_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07004__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout390_X net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout867_A _01724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout488_X net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold12 keypad.debounce.debounce\[2\] vssd1 vssd1 vccd1 vccd1 net1360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 screen.counter.ack2 vssd1 vssd1 vccd1 vccd1 net1371 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12502__S net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold34 screen.controlBus\[10\] vssd1 vssd1 vccd1 vccd1 net1382 sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ net448 _03813_ vssd1 vssd1 vccd1 vccd1 _03814_ sky130_fd_sc_hd__or2_1
XANTENNA__08488__A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06763__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold45 net116 vssd1 vssd1 vccd1 vccd1 net1393 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 net57 vssd1 vssd1 vccd1 vccd1 net1404 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07960__B1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold67 screen.controlBus\[14\] vssd1 vssd1 vccd1 vccd1 net1415 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold78 net46 vssd1 vssd1 vccd1 vccd1 net1426 sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ datapath.rf.registers\[17\]\[12\] net748 net678 datapath.rf.registers\[29\]\[12\]
+ _02762_ vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__a221o_1
Xhold89 net48 vssd1 vssd1 vccd1 vccd1 net1437 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout655_X net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08504__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11118__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10940_ _05678_ _05679_ vssd1 vssd1 vccd1 vccd1 _05680_ sky130_fd_sc_hd__nand2_1
XANTENNA__08000__B net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10871_ net898 _04084_ _05620_ net600 vssd1 vssd1 vccd1 vccd1 _05621_ sky130_fd_sc_hd__a211o_2
XANTENNA_fanout822_X net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12610_ net499 _06454_ _06455_ net503 net1878 vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__a32o_1
X_13590_ clknet_leaf_139_clk _00400_ net1099 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_12541_ _06395_ _06396_ _06397_ vssd1 vssd1 vccd1 vccd1 _06398_ sky130_fd_sc_hd__or3_1
XANTENNA__11811__A2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12472_ net165 _05992_ net127 screen.register.currentXbus\[28\] vssd1 vssd1 vccd1
+ vccd1 _00874_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07491__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14211_ clknet_leaf_44_clk datapath.multiplication_module.multiplicand_i_n\[22\]
+ net1177 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11423_ net255 net1871 net515 vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__mux2_1
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07779__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_9 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14142_ clknet_leaf_144_clk _00899_ net1085 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11354_ net267 net2482 net520 vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__mux2_1
XANTENNA__07243__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10305_ _04564_ _04580_ net890 vssd1 vssd1 vccd1 vccd1 _05141_ sky130_fd_sc_hd__a21o_1
XFILLER_140_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14073_ clknet_leaf_122_clk _00840_ net1214 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11285_ net266 net2614 net524 vssd1 vssd1 vccd1 vccd1 _00333_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13024_ net1714 net183 net390 vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_5_Left_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10236_ datapath.PC\[28\] net1258 _05068_ _05071_ vssd1 vssd1 vccd1 vccd1 _05072_
+ sky130_fd_sc_hd__a2bb2o_1
Xfanout1010 net1011 vssd1 vssd1 vccd1 vccd1 net1010 sky130_fd_sc_hd__buf_2
Xfanout1021 _01566_ vssd1 vssd1 vccd1 vccd1 net1021 sky130_fd_sc_hd__buf_2
XFILLER_67_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10167_ datapath.PC\[16\] _04178_ net467 vssd1 vssd1 vccd1 vccd1 _05003_ sky130_fd_sc_hd__mux2_1
Xfanout1032 _01565_ vssd1 vssd1 vccd1 vccd1 net1032 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10280__X _05116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1043 net1044 vssd1 vssd1 vccd1 vccd1 net1043 sky130_fd_sc_hd__clkbuf_4
Xfanout1054 net1058 vssd1 vssd1 vccd1 vccd1 net1054 sky130_fd_sc_hd__clkbuf_4
XFILLER_121_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1065 net1066 vssd1 vssd1 vccd1 vccd1 net1065 sky130_fd_sc_hd__buf_2
XANTENNA__12288__C1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1076 net1084 vssd1 vssd1 vccd1 vccd1 net1076 sky130_fd_sc_hd__clkbuf_4
X_10098_ datapath.PC\[27\] net468 net1038 vssd1 vssd1 vccd1 vccd1 _04934_ sky130_fd_sc_hd__o21ai_1
Xfanout1087 net1092 vssd1 vssd1 vccd1 vccd1 net1087 sky130_fd_sc_hd__clkbuf_2
Xfanout1098 net1101 vssd1 vssd1 vccd1 vccd1 net1098 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11028__S net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13926_ clknet_leaf_96_clk _00704_ net1226 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10302__A2 _04580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07703__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13857_ clknet_leaf_71_clk _00661_ net1244 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12648__A datapath.mulitply_result\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12808_ net2261 net266 net492 vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__mux2_1
XANTENNA__12055__A2 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13788_ clknet_leaf_73_clk _00597_ net1243 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12739_ net1876 net281 net405 vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07482__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06933__X _01769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11015__A0 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14293__RESET_B net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14409_ clknet_leaf_20_clk _01114_ net1165 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_156_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14222__RESET_B net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold504 datapath.rf.registers\[12\]\[19\] vssd1 vssd1 vccd1 vccd1 net1852 sky130_fd_sc_hd__dlygate4sd3_1
Xhold515 datapath.rf.registers\[5\]\[20\] vssd1 vssd1 vccd1 vccd1 net1863 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold526 datapath.rf.registers\[26\]\[21\] vssd1 vssd1 vccd1 vccd1 net1874 sky130_fd_sc_hd__dlygate4sd3_1
Xhold537 datapath.rf.registers\[20\]\[25\] vssd1 vssd1 vccd1 vccd1 net1885 sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 datapath.rf.registers\[5\]\[1\] vssd1 vssd1 vccd1 vccd1 net1896 sky130_fd_sc_hd__dlygate4sd3_1
Xhold559 datapath.rf.registers\[5\]\[8\] vssd1 vssd1 vccd1 vccd1 net1907 sky130_fd_sc_hd__dlygate4sd3_1
X_09950_ _04779_ _04785_ vssd1 vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__nand2_1
X_08901_ net1267 datapath.PC\[10\] _03736_ vssd1 vssd1 vccd1 vccd1 _03737_ sky130_fd_sc_hd__or3_1
XANTENNA_clkbuf_4_9_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09881_ datapath.PC\[28\] net595 vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__and2_1
XFILLER_97_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08832_ _03661_ net347 net575 vssd1 vssd1 vccd1 vccd1 _03668_ sky130_fd_sc_hd__o21a_1
XFILLER_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1204 datapath.rf.registers\[16\]\[14\] vssd1 vssd1 vccd1 vccd1 net2552 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1215 datapath.rf.registers\[30\]\[0\] vssd1 vssd1 vccd1 vccd1 net2563 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1226 datapath.rf.registers\[16\]\[27\] vssd1 vssd1 vccd1 vccd1 net2574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1237 screen.register.currentXbus\[1\] vssd1 vssd1 vccd1 vccd1 net2585 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1248 screen.register.currentYbus\[22\] vssd1 vssd1 vccd1 vccd1 net2596 sky130_fd_sc_hd__dlygate4sd3_1
X_08763_ _03481_ _03598_ _01859_ vssd1 vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08101__A _02913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1259 mmio.memload_or_instruction\[15\] vssd1 vssd1 vccd1 vccd1 net2607 sky130_fd_sc_hd__dlygate4sd3_1
X_07714_ datapath.rf.registers\[23\]\[16\] net940 net922 vssd1 vssd1 vccd1 vccd1 _02550_
+ sky130_fd_sc_hd__and3_1
XFILLER_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12294__A2 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08694_ _03529_ vssd1 vssd1 vccd1 vccd1 _03530_ sky130_fd_sc_hd__inv_2
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07645_ datapath.rf.registers\[24\]\[18\] net766 net706 datapath.rf.registers\[10\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02481_ sky130_fd_sc_hd__a22o_1
XFILLER_25_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1092_A net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13153__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07576_ datapath.rf.registers\[5\]\[19\] net820 _02395_ _02398_ _02399_ vssd1 vssd1
+ vccd1 vccd1 _02412_ sky130_fd_sc_hd__a2111o_1
XFILLER_34_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09315_ net557 net576 net546 _02466_ vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__o211a_1
XFILLER_139_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12992__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout615_A net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09246_ _04075_ _04077_ _04081_ vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_32_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07473__A2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08771__A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09177_ net338 _04007_ _04012_ net322 vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout403_X net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08490__B net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11401__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08128_ datapath.rf.registers\[30\]\[8\] net761 net696 datapath.rf.registers\[8\]\[8\]
+ _02963_ vssd1 vssd1 vccd1 vccd1 _02964_ sky130_fd_sc_hd__a221o_1
XFILLER_147_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07225__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout984_A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08059_ datapath.rf.registers\[18\]\[9\] net977 net951 vssd1 vssd1 vccd1 vccd1 _02895_
+ sky130_fd_sc_hd__and3_1
Xoutput46 net46 vssd1 vssd1 vccd1 vccd1 ADR_O[15] sky130_fd_sc_hd__buf_2
Xoutput57 net57 vssd1 vssd1 vccd1 vccd1 ADR_O[25] sky130_fd_sc_hd__buf_2
X_11070_ _01643_ _01663_ vssd1 vssd1 vccd1 vccd1 _05712_ sky130_fd_sc_hd__nand2_1
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 ADR_O[6] sky130_fd_sc_hd__buf_2
XFILLER_131_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 DAT_O[15] sky130_fd_sc_hd__buf_2
XANTENNA_fanout772_X net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08186__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10021_ _04856_ _04855_ vssd1 vssd1 vccd1 vccd1 _04857_ sky130_fd_sc_hd__and2b_1
XFILLER_103_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07933__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06736__B2 _01441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07553__C net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11972_ _05332_ _05795_ _05843_ _05849_ _06016_ vssd1 vssd1 vccd1 vccd1 _06017_ sky130_fd_sc_hd__a311o_4
XANTENNA__12285__A2 _06254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_2_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13711_ clknet_leaf_26_clk _00521_ net1137 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10923_ datapath.PC\[27\] datapath.PC\[28\] _05654_ vssd1 vssd1 vccd1 vccd1 _05665_
+ sky130_fd_sc_hd__and3_1
X_14691_ clknet_leaf_138_clk _01396_ net1100 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13063__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08665__B _02284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13642_ clknet_leaf_59_clk _00452_ net1168 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10854_ datapath.PC\[18\] _05600_ vssd1 vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__xnor2_1
XFILLER_71_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13573_ clknet_leaf_116_clk _00383_ net1188 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10785_ net284 net2272 net544 vssd1 vssd1 vccd1 vccd1 _00009_ sky130_fd_sc_hd__mux2_1
XANTENNA__08110__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11796__B2 _01443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09777__A net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12524_ _06382_ _06383_ vssd1 vssd1 vccd1 vccd1 _06384_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07464__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12455_ net166 _05958_ net128 screen.register.currentXbus\[11\] vssd1 vssd1 vccd1
+ vccd1 _00857_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_97_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06913__B net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11311__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11406_ net1707 net183 net411 vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__mux2_1
XFILLER_125_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07216__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12386_ net2260 net133 _06340_ vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10435__B _05240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06632__C datapath.ru.latched_instruction\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14125_ clknet_leaf_16_clk _00882_ net1106 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11337_ net1687 net178 net416 vssd1 vssd1 vccd1 vccd1 _00382_ sky130_fd_sc_hd__mux2_1
XFILLER_126_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10771__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14056_ clknet_leaf_95_clk _00823_ net1216 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_98_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11268_ net186 net2388 net419 vssd1 vssd1 vccd1 vccd1 _00317_ sky130_fd_sc_hd__mux2_1
XANTENNA__08177__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13007_ net2170 net262 net391 vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__mux2_1
X_10219_ _04626_ _04645_ vssd1 vssd1 vccd1 vccd1 _05055_ sky130_fd_sc_hd__xnor2_1
X_11199_ net198 net1776 net424 vssd1 vssd1 vccd1 vccd1 _00251_ sky130_fd_sc_hd__mux2_1
XANTENNA__07924__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06928__X _01764_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13909_ clknet_leaf_43_clk net1355 net1149 vssd1 vssd1 vccd1 vccd1 keypad.debounce.debounce\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_59_Left_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07430_ datapath.rf.registers\[17\]\[22\] net746 net687 datapath.rf.registers\[31\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__a22o_1
XFILLER_63_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_926 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07361_ datapath.rf.registers\[21\]\[23\] net945 net921 vssd1 vssd1 vccd1 vccd1 _02197_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_44_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09100_ _03797_ _03802_ net341 vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__mux2_1
X_07292_ datapath.rf.registers\[3\]\[25\] net772 net685 datapath.rf.registers\[27\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__a22o_1
XANTENNA__06663__X _01502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09031_ _03467_ _03866_ vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11221__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_68_Left_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold301 datapath.rf.registers\[12\]\[10\] vssd1 vssd1 vccd1 vccd1 net1649 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold312 datapath.rf.registers\[15\]\[2\] vssd1 vssd1 vccd1 vccd1 net1660 sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 datapath.rf.registers\[7\]\[4\] vssd1 vssd1 vccd1 vccd1 net1671 sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 datapath.multiplication_module.multiplicand_i\[11\] vssd1 vssd1 vccd1 vccd1
+ net1682 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10913__X _05657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold345 datapath.rf.registers\[1\]\[3\] vssd1 vssd1 vccd1 vccd1 net1693 sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 datapath.rf.registers\[15\]\[27\] vssd1 vssd1 vccd1 vccd1 net1704 sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 datapath.rf.registers\[5\]\[27\] vssd1 vssd1 vccd1 vccd1 net1715 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10762__A2 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold378 datapath.rf.registers\[4\]\[27\] vssd1 vssd1 vccd1 vccd1 net1726 sky130_fd_sc_hd__dlygate4sd3_1
Xhold389 datapath.rf.registers\[6\]\[10\] vssd1 vssd1 vccd1 vccd1 net1737 sky130_fd_sc_hd__dlygate4sd3_1
X_09933_ net1268 _03077_ vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__and2_1
XFILLER_132_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout803 _01769_ vssd1 vssd1 vccd1 vccd1 net803 sky130_fd_sc_hd__buf_2
Xfanout814 _01760_ vssd1 vssd1 vccd1 vccd1 net814 sky130_fd_sc_hd__clkbuf_8
XFILLER_113_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout825 _01753_ vssd1 vssd1 vccd1 vccd1 net825 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08168__B1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13148__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout398_A net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout836 _01743_ vssd1 vssd1 vccd1 vccd1 net836 sky130_fd_sc_hd__buf_4
X_09864_ _02637_ _02683_ _04698_ _04699_ _02636_ vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__o2111a_1
Xfanout847 _01737_ vssd1 vssd1 vccd1 vccd1 net847 sky130_fd_sc_hd__clkbuf_8
Xfanout858 net859 vssd1 vssd1 vccd1 vccd1 net858 sky130_fd_sc_hd__clkbuf_8
XFILLER_133_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1001 datapath.rf.registers\[2\]\[6\] vssd1 vssd1 vccd1 vccd1 net2349 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1105_A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout869 net871 vssd1 vssd1 vccd1 vccd1 net869 sky130_fd_sc_hd__buf_4
Xhold1012 mmio.memload_or_instruction\[14\] vssd1 vssd1 vccd1 vccd1 net2360 sky130_fd_sc_hd__dlygate4sd3_1
X_08815_ net972 _03359_ _03643_ vssd1 vssd1 vccd1 vccd1 _03651_ sky130_fd_sc_hd__mux2_1
Xhold1023 datapath.rf.registers\[11\]\[20\] vssd1 vssd1 vccd1 vccd1 net2371 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_86_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12987__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09795_ _03596_ _04628_ _04630_ net579 vssd1 vssd1 vccd1 vccd1 _04631_ sky130_fd_sc_hd__o211a_1
Xhold1034 datapath.rf.registers\[4\]\[11\] vssd1 vssd1 vccd1 vccd1 net2382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1045 datapath.rf.registers\[12\]\[29\] vssd1 vssd1 vccd1 vccd1 net2393 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout565_A _01786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1056 datapath.rf.registers\[0\]\[5\] vssd1 vssd1 vccd1 vccd1 net2404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1067 datapath.rf.registers\[28\]\[22\] vssd1 vssd1 vccd1 vccd1 net2415 sky130_fd_sc_hd__dlygate4sd3_1
X_08746_ _03513_ _03514_ _03579_ _03511_ _03509_ vssd1 vssd1 vccd1 vccd1 _03582_ sky130_fd_sc_hd__a311o_1
XPHY_EDGE_ROW_77_Left_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1078 datapath.rf.registers\[20\]\[10\] vssd1 vssd1 vccd1 vccd1 net2426 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1089 datapath.rf.registers\[26\]\[5\] vssd1 vssd1 vccd1 vccd1 net2437 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08766__A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout732_A _01811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08677_ _02489_ _02490_ vssd1 vssd1 vccd1 vccd1 _03513_ sky130_fd_sc_hd__or2_2
XFILLER_26_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07628_ _02447_ _02461_ _02462_ _02463_ vssd1 vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__or4_1
XANTENNA__12019__A2 _05778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10300__S net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07694__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout520_X net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07559_ datapath.rf.registers\[21\]\[19\] net947 net924 vssd1 vssd1 vccd1 vccd1 _02395_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1262_X net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10570_ _05388_ _05391_ _05393_ vssd1 vssd1 vccd1 vccd1 screen.register.xFill sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09229_ net372 _03921_ vssd1 vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__nor2_1
XFILLER_154_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_86_Left_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10536__A _05085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11131__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12240_ screen.counter.currentCt\[17\] _06233_ screen.counter.currentCt\[18\] vssd1
+ vssd1 vccd1 vccd1 _06236_ sky130_fd_sc_hd__a21oi_1
XFILLER_5_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout987_X net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10202__A1 _03978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12171_ net1272 _06192_ _06193_ vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__o21a_1
XFILLER_123_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11122_ net248 net2225 net427 vssd1 vssd1 vccd1 vccd1 _00177_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_92_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold890 datapath.rf.registers\[29\]\[10\] vssd1 vssd1 vccd1 vccd1 net2238 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08159__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13058__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11053_ net249 net2428 net431 vssd1 vssd1 vccd1 vccd1 _00113_ sky130_fd_sc_hd__mux2_1
XANTENNA__07906__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11702__A1 _04909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10004_ _04788_ _04790_ vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__xnor2_1
XFILLER_49_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12897__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_95_Left_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09108__C1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08676__A _02466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11955_ screen.counter.ct\[5\] _06000_ vssd1 vssd1 vccd1 vccd1 _06001_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_106_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12198__A _06168_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08331__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08395__B _03228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10906_ _03916_ _05650_ net902 vssd1 vssd1 vccd1 vccd1 _05651_ sky130_fd_sc_hd__mux2_2
X_14674_ clknet_leaf_32_clk _01379_ net1126 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11886_ net137 _05954_ _05953_ vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06893__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13625_ clknet_leaf_31_clk _00435_ net1124 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10837_ _01510_ net653 _05590_ _05591_ vssd1 vssd1 vccd1 vccd1 _05592_ sky130_fd_sc_hd__o22a_2
XFILLER_32_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11769__B2 _01954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07437__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13556_ clknet_leaf_93_clk _00366_ net1212 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06924__A net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10768_ net901 _05532_ vssd1 vssd1 vccd1 vccd1 _05533_ sky130_fd_sc_hd__nand2_1
X_12507_ net181 net2334 net509 vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__mux2_1
XANTENNA__10441__A1 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13487_ clknet_leaf_25_clk _00297_ net1137 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10699_ net1471 _03170_ net570 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i_n\[4\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA__11041__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12438_ net1390 net132 _06366_ vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__a21o_1
XFILLER_8_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07458__C net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10880__S net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12369_ datapath.PC\[31\] net309 _06330_ _03756_ vssd1 vssd1 vccd1 vccd1 _00810_
+ sky130_fd_sc_hd__a22o_1
XFILLER_113_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14108_ clknet_leaf_110_clk _00874_ net1202 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07070__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06930_ net974 net939 vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__and2_1
XFILLER_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14039_ clknet_leaf_85_clk _00808_ net1258 vssd1 vssd1 vccd1 vccd1 datapath.PC\[29\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_68_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_143_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06861_ datapath.ru.latched_instruction\[25\] _01604_ _01693_ _01694_ _01696_ vssd1
+ vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__a2111o_1
XFILLER_83_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08570__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08600_ _03430_ _03434_ _02984_ vssd1 vssd1 vccd1 vccd1 _03436_ sky130_fd_sc_hd__a21oi_1
X_06792_ _01576_ _01584_ _01585_ _01624_ vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__or4_1
X_09580_ net360 _04415_ vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__nor2_1
XFILLER_55_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08531_ datapath.rf.registers\[14\]\[0\] net831 net812 datapath.rf.registers\[13\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03367_ sky130_fd_sc_hd__a22o_1
XANTENNA__08322__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11216__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08462_ _03262_ _03293_ _03294_ vssd1 vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__and3_1
XANTENNA__07676__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08873__A1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07413_ datapath.rf.registers\[8\]\[22\] net876 net832 datapath.rf.registers\[30\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__a22o_1
XFILLER_149_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08393_ _03228_ vssd1 vssd1 vccd1 vccd1 _03229_ sky130_fd_sc_hd__inv_2
XANTENNA__10908__X _05653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout146_A net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07344_ datapath.rf.registers\[13\]\[24\] net692 net684 datapath.rf.registers\[27\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__a22o_1
XFILLER_148_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07428__A2 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07275_ datapath.rf.registers\[16\]\[25\] net862 net802 datapath.rf.registers\[3\]\[25\]
+ _02095_ vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_154_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1055_A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09014_ _03667_ _03848_ _03849_ _03839_ vssd1 vssd1 vccd1 vccd1 _03850_ sky130_fd_sc_hd__o22a_1
XANTENNA__11739__X _05891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold120 datapath.multiplication_module.multiplier_i\[8\] vssd1 vssd1 vccd1 vccd1
+ net1468 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10790__S net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold131 net119 vssd1 vssd1 vccd1 vccd1 net1479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 mmio.memload_or_instruction\[9\] vssd1 vssd1 vccd1 vccd1 net1490 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1222_A net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold153 net93 vssd1 vssd1 vccd1 vccd1 net1501 sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 datapath.rf.registers\[0\]\[13\] vssd1 vssd1 vccd1 vccd1 net1512 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07061__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold175 screen.counter.currentCt\[4\] vssd1 vssd1 vccd1 vccd1 net1523 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07600__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold186 datapath.multiplication_module.multiplicand_i\[29\] vssd1 vssd1 vccd1 vccd1
+ net1534 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout682_A _01828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout600 datapath.MUL_EN vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__clkbuf_4
Xhold197 datapath.rf.registers\[7\]\[2\] vssd1 vssd1 vccd1 vccd1 net1545 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout611 _01782_ vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__buf_2
X_09916_ net1266 _04751_ vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__and2_1
Xfanout622 MemRead vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout633 _01705_ vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__clkbuf_4
XFILLER_132_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout644 net646 vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__clkbuf_4
Xfanout655 _01592_ vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08199__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout666 net667 vssd1 vssd1 vccd1 vccd1 net666 sky130_fd_sc_hd__buf_4
XANTENNA__11696__B1 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09847_ _04682_ vssd1 vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__inv_2
Xfanout677 net678 vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__buf_4
XANTENNA_fanout470_X net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout688 net690 vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__buf_2
XFILLER_59_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_70_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout699 net701 vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout947_A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11915__A _02438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09778_ net649 _04613_ net439 vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__a21o_1
X_08729_ _02984_ _03433_ vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__or2_2
XFILLER_26_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout735_X net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11126__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06728__B net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11740_ net1515 net143 net138 _03417_ vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__a22o_1
XFILLER_53_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10120__B1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11671_ _05240_ net154 net150 net1411 vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout902_X net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13410_ clknet_leaf_1_clk _00220_ net1056 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10622_ net121 net123 net124 net122 vssd1 vssd1 vccd1 vccd1 _05442_ sky130_fd_sc_hd__nor4b_1
X_14390_ clknet_leaf_141_clk _01095_ net1096 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13341_ clknet_leaf_147_clk _00151_ net1064 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10553_ net35 net36 vssd1 vssd1 vccd1 vccd1 _05380_ sky130_fd_sc_hd__nor2_1
XANTENNA__07559__B net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10266__A net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08092__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13272_ clknet_leaf_4_clk _00082_ net1069 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10484_ _05307_ _05310_ _05313_ vssd1 vssd1 vccd1 vccd1 _05314_ sky130_fd_sc_hd__and3_1
X_12223_ net1513 _06223_ _06225_ vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__a21oi_1
XFILLER_154_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07052__B1 _01887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12154_ net1278 net1279 _06180_ net1277 vssd1 vssd1 vccd1 vccd1 _06183_ sky130_fd_sc_hd__a31o_1
XFILLER_2_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11105_ _05514_ _05707_ vssd1 vssd1 vccd1 vccd1 _05715_ sky130_fd_sc_hd__nor2_2
XFILLER_151_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12085_ _05324_ _05767_ _05847_ _06024_ _06073_ vssd1 vssd1 vccd1 vccd1 _06124_ sky130_fd_sc_hd__a2111o_1
XFILLER_1_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11036_ _05692_ _05707_ vssd1 vssd1 vccd1 vccd1 _05710_ sky130_fd_sc_hd__nor2_1
XFILLER_103_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06919__A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12987_ net198 net2392 net480 vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__mux2_1
XANTENNA__08304__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09501__C1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11938_ net2630 net162 vssd1 vssd1 vccd1 vccd1 _05989_ sky130_fd_sc_hd__nand2_1
XFILLER_73_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08855__A1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14657_ clknet_leaf_25_clk _01362_ net1159 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11869_ screen.register.currentYbus\[4\] net161 vssd1 vssd1 vccd1 vccd1 _05943_ sky130_fd_sc_hd__nand2_1
X_13608_ clknet_leaf_91_clk _00418_ net1233 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14588_ clknet_leaf_7_clk _01293_ net1071 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_119_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08572__C _01823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13539_ clknet_leaf_120_clk _00349_ net1199 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_145_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xteam_04_1308 vssd1 vssd1 vccd1 vccd1 team_04_1308/HI gpio_oeb[17] sky130_fd_sc_hd__conb_1
X_07060_ datapath.rf.registers\[3\]\[30\] net772 net708 datapath.rf.registers\[10\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_136_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xteam_04_1319 vssd1 vssd1 vccd1 vccd1 team_04_1319/HI gpio_out[23] sky130_fd_sc_hd__conb_1
XANTENNA__07291__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07830__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07043__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07962_ datapath.rf.registers\[20\]\[11\] net840 _02784_ _02785_ _02786_ vssd1 vssd1
+ vccd1 vccd1 _02798_ sky130_fd_sc_hd__a2111o_1
X_09701_ _04534_ _04536_ vssd1 vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__and2_1
X_06913_ net955 net920 vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__and2_1
XFILLER_68_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11678__B1 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07893_ datapath.rf.registers\[29\]\[12\] net975 net917 vssd1 vssd1 vccd1 vccd1 _02729_
+ sky130_fd_sc_hd__and3_1
XFILLER_110_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08543__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09632_ net905 _03561_ net624 _03560_ vssd1 vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__a22o_1
XANTENNA__12330__S net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06844_ _01412_ net993 _01642_ _01674_ vssd1 vssd1 vccd1 vccd1 _01680_ sky130_fd_sc_hd__a31o_1
XANTENNA__07897__A2 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09563_ net609 _04397_ _04398_ net580 vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__a22o_1
X_06775_ datapath.ru.latched_instruction\[12\] _01480_ net1017 vssd1 vssd1 vccd1 vccd1
+ _01612_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout263_A _05575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08514_ datapath.rf.registers\[31\]\[1\] net963 _01825_ vssd1 vssd1 vccd1 vccd1 _03350_
+ sky130_fd_sc_hd__and3_1
X_09494_ net904 _03554_ vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__or2_1
X_08445_ datapath.rf.registers\[26\]\[2\] net781 net769 datapath.rf.registers\[24\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout430_A net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10785__S net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_42_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1172_A net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout149_X net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13161__S net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout528_A _05721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13789__RESET_B net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08376_ datapath.rf.registers\[25\]\[3\] net729 net682 datapath.rf.registers\[6\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03212_ sky130_fd_sc_hd__a22o_1
XFILLER_149_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07327_ datapath.rf.registers\[12\]\[24\] net827 net790 datapath.rf.registers\[18\]\[24\]
+ _02162_ vssd1 vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__a221o_1
XANTENNA__10086__A net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1058_X net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09875__A net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07258_ _02069_ _02091_ vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_57_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07821__A2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout897_A _01626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12505__S net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07189_ datapath.rf.registers\[0\]\[27\] net871 _02012_ _02024_ vssd1 vssd1 vccd1
+ vccd1 _02025_ sky130_fd_sc_hd__o22a_4
XANTENNA_clkbuf_leaf_100_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1225_X net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07034__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout685_X net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08782__A0 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout430 net433 vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08003__B net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout441 net443 vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__clkbuf_4
XFILLER_120_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout452 _03658_ vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_115_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout463 _03149_ vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__buf_4
XANTENNA_fanout852_X net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout474 net475 vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__buf_4
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08534__B1 _01743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout485 _06554_ vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__buf_4
X_12910_ net2552 net252 net482 vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__mux2_1
Xfanout496 _06550_ vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__clkbuf_8
XFILLER_47_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13890_ clknet_leaf_44_clk keypad.decode.button_n\[1\] net1152 vssd1 vssd1 vccd1
+ vccd1 button\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_73_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13738__SET_B net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12841_ net268 net1904 net488 vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772_ net278 net2200 net497 vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__mux2_1
X_14511_ clknet_leaf_27_clk _01216_ net1132 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11723_ net9 net1033 net1023 net1554 vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__o22a_1
XANTENNA__11651__Y _05874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13071__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14442_ clknet_leaf_58_clk _01147_ net1167 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11654_ net1475 _05875_ _05876_ vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__a21o_1
XFILLER_156_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06905__C net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10605_ _05419_ _05421_ _05425_ vssd1 vssd1 vccd1 vccd1 _05426_ sky130_fd_sc_hd__or3_1
X_14373_ clknet_leaf_117_clk _01078_ net1190 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11585_ net1276 net1277 screen.counter.ct\[11\] screen.counter.ct\[10\] vssd1 vssd1
+ vccd1 vccd1 _05809_ sky130_fd_sc_hd__nand4_1
XANTENNA__12763__X _06550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13324_ clknet_leaf_133_clk _00134_ net1104 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10536_ _05085_ _05281_ vssd1 vssd1 vccd1 vccd1 _05365_ sky130_fd_sc_hd__nor2_1
XANTENNA__07812__A2 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13255_ clknet_leaf_137_clk _00065_ net1097 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09014__A1 _03667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_108_Right_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10467_ net1270 screen.counter.ct\[16\] _05295_ _05296_ vssd1 vssd1 vccd1 vccd1 _05297_
+ sky130_fd_sc_hd__or4_1
X_12206_ _06168_ _06213_ _06214_ vssd1 vssd1 vccd1 vccd1 _00763_ sky130_fd_sc_hd__nor3_1
X_13186_ net1807 vssd1 vssd1 vccd1 vccd1 _01008_ sky130_fd_sc_hd__clkbuf_1
X_10398_ net631 _04666_ vssd1 vssd1 vccd1 vccd1 _05234_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_131_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12137_ _05753_ _05774_ vssd1 vssd1 vccd1 vccd1 _06173_ sky130_fd_sc_hd__nand2_1
XFILLER_151_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09317__A2 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12068_ screen.register.currentXbus\[29\] net996 net995 screen.register.currentXbus\[5\]
+ _06107_ vssd1 vssd1 vccd1 vccd1 _06108_ sky130_fd_sc_hd__a221o_1
XFILLER_38_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14247__RESET_B net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11019_ net249 net2002 net539 vssd1 vssd1 vccd1 vccd1 _00081_ sky130_fd_sc_hd__mux2_1
XFILLER_93_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07879__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08567__C _01825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_32_Left_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06936__X _01772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08230_ datapath.rf.registers\[17\]\[6\] net746 net738 datapath.rf.registers\[16\]\[6\]
+ _03065_ vssd1 vssd1 vccd1 vccd1 _03066_ sky130_fd_sc_hd__a221o_1
XANTENNA__09031__Y _03867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08161_ datapath.rf.registers\[6\]\[7\] net825 net797 datapath.rf.registers\[29\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02997_ sky130_fd_sc_hd__a22o_1
XFILLER_118_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07112_ datapath.rf.registers\[17\]\[29\] net747 net692 datapath.rf.registers\[13\]\[29\]
+ _01937_ vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_151_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08092_ datapath.rf.registers\[18\]\[9\] net724 net704 datapath.rf.registers\[9\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02928_ sky130_fd_sc_hd__a22o_1
XFILLER_9_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload40 clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 clkload40/Y sky130_fd_sc_hd__clkinv_2
X_07043_ datapath.rf.registers\[7\]\[30\] net818 net874 vssd1 vssd1 vccd1 vccd1 _01879_
+ sky130_fd_sc_hd__a21o_1
Xclkload51 clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 clkload51/Y sky130_fd_sc_hd__inv_6
XANTENNA__12325__S net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_41_Left_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload62 clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 clkload62/Y sky130_fd_sc_hd__clkinv_4
Xclkload73 clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 clkload73/Y sky130_fd_sc_hd__inv_6
XFILLER_133_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06831__B net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload84 clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 clkload84/Y sky130_fd_sc_hd__inv_8
Xclkload95 clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 clkload95/Y sky130_fd_sc_hd__bufinv_16
XFILLER_115_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10921__X _05664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08994_ net632 _03829_ vssd1 vssd1 vccd1 vccd1 _03830_ sky130_fd_sc_hd__nand2_1
X_07945_ datapath.rf.registers\[22\]\[11\] net952 net924 vssd1 vssd1 vccd1 vccd1 _02781_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_149_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout478_A _06556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13156__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07662__B net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07876_ datapath.rf.registers\[23\]\[13\] net699 net676 datapath.rf.registers\[29\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__a22o_1
XFILLER_83_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09615_ _03557_ _03558_ vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__xnor2_1
X_06827_ _01467_ _01568_ net1029 datapath.ru.latched_instruction\[8\] vssd1 vssd1
+ vccd1 vccd1 _01663_ sky130_fd_sc_hd__a2bb2o_2
XANTENNA__12995__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09546_ net371 _04379_ _04380_ _04381_ net329 vssd1 vssd1 vccd1 vccd1 _04382_ sky130_fd_sc_hd__a221o_1
XFILLER_83_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06758_ datapath.ru.latched_instruction\[26\] net1032 _01568_ _01504_ vssd1 vssd1
+ vccd1 vccd1 _01595_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__11912__B net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout812_A _01765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08295__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09477_ net359 _04311_ _04312_ net345 vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__a31o_1
X_06689_ _01414_ _01527_ vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout433_X net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11404__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08428_ datapath.ru.latched_instruction\[9\] net1029 _01659_ vssd1 vssd1 vccd1 vccd1
+ _03264_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_82_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload1 clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clkload1/X sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout600_X net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08359_ datapath.rf.registers\[1\]\[3\] net848 _03184_ _03186_ _03189_ vssd1 vssd1
+ vccd1 vccd1 _03195_ sky130_fd_sc_hd__a2111o_1
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07255__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11370_ net185 net2306 net518 vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__mux2_1
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10321_ net1268 net1259 _05153_ _05156_ vssd1 vssd1 vccd1 vccd1 _05157_ sky130_fd_sc_hd__o22a_1
XFILLER_153_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07007__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13040_ net266 net2397 net476 vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__mux2_1
X_10252_ datapath.PC\[11\] _03737_ vssd1 vssd1 vccd1 vccd1 _05088_ sky130_fd_sc_hd__nand2_1
XFILLER_1_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07556__C net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10263__B _04272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10183_ net1264 net1260 _05015_ _05018_ vssd1 vssd1 vccd1 vccd1 _05019_ sky130_fd_sc_hd__o22a_1
Xfanout1203 net1204 vssd1 vssd1 vccd1 vccd1 net1203 sky130_fd_sc_hd__clkbuf_2
Xfanout1214 net1216 vssd1 vssd1 vccd1 vccd1 net1214 sky130_fd_sc_hd__clkbuf_4
Xfanout1225 net1231 vssd1 vssd1 vccd1 vccd1 net1225 sky130_fd_sc_hd__clkbuf_4
Xfanout1236 net1238 vssd1 vssd1 vccd1 vccd1 net1236 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input39_A nrst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1247 net1248 vssd1 vssd1 vccd1 vccd1 net1247 sky130_fd_sc_hd__clkbuf_4
Xfanout1258 net1259 vssd1 vssd1 vccd1 vccd1 net1258 sky130_fd_sc_hd__buf_2
Xfanout260 net261 vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_89_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13066__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout271 _05564_ vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__buf_1
Xfanout1269 datapath.PC\[2\] vssd1 vssd1 vccd1 vccd1 net1269 sky130_fd_sc_hd__buf_2
XANTENNA__12303__B2 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout282 net285 vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__clkbuf_2
X_13942_ clknet_leaf_96_clk _00720_ net1226 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[26\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout293 _05541_ vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09180__A0 _03805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13873_ clknet_leaf_53_clk _00677_ net1182 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[17\]
+ sky130_fd_sc_hd__dfrtp_4
X_12824_ net2113 net186 net491 vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__mux2_1
XANTENNA__12067__B1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12755_ net1771 net201 net403 vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__mux2_1
XANTENNA__11314__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11706_ net1291 net1035 mmio.wishbone.prev_BUSY_O vssd1 vssd1 vccd1 vccd1 _05890_
+ sky130_fd_sc_hd__or3b_1
X_12686_ datapath.mulitply_result\[29\] datapath.multiplication_module.multiplicand_i\[29\]
+ vssd1 vssd1 vccd1 vccd1 _06519_ sky130_fd_sc_hd__nor2_1
XANTENNA__10438__B _01702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14425_ clknet_leaf_31_clk _01130_ net1124 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_11637_ _05358_ _05860_ vssd1 vssd1 vccd1 vccd1 _05861_ sky130_fd_sc_hd__and2_1
XANTENNA__08038__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07246__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14356_ clknet_leaf_93_clk _01061_ net1211 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_155_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11568_ net1008 _05758_ vssd1 vssd1 vccd1 vccd1 _05792_ sky130_fd_sc_hd__nor2_1
XANTENNA__06932__A net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold708 datapath.rf.registers\[16\]\[13\] vssd1 vssd1 vccd1 vccd1 net2056 sky130_fd_sc_hd__dlygate4sd3_1
X_13307_ clknet_leaf_36_clk _00117_ net1135 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10519_ _05335_ _05343_ vssd1 vssd1 vccd1 vccd1 _05349_ sky130_fd_sc_hd__nor2_1
Xhold719 datapath.rf.registers\[18\]\[13\] vssd1 vssd1 vccd1 vccd1 net2067 sky130_fd_sc_hd__dlygate4sd3_1
X_14287_ clknet_leaf_26_clk _00992_ net1155 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_11499_ net214 net2041 net510 vssd1 vssd1 vccd1 vccd1 _00535_ sky130_fd_sc_hd__mux2_1
X_13238_ clknet_leaf_137_clk _00048_ net1097 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10173__B _04987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08210__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13169_ net2241 vssd1 vssd1 vccd1 vccd1 _00991_ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14081__RESET_B net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08578__B net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07730_ _02559_ _02561_ _02563_ _02565_ vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__or4_2
X_07661_ datapath.rf.registers\[9\]\[17\] net982 net944 vssd1 vssd1 vccd1 vccd1 _02497_
+ sky130_fd_sc_hd__and3_1
XFILLER_93_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09400_ _03522_ net626 _04235_ net643 vssd1 vssd1 vccd1 vccd1 _04236_ sky130_fd_sc_hd__a211o_1
X_06612_ mmio.memload_or_instruction\[17\] net1048 vssd1 vssd1 vccd1 vccd1 _01451_
+ sky130_fd_sc_hd__and2_2
XANTENNA__06666__X _01505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07592_ datapath.rf.registers\[9\]\[19\] net704 _02426_ _02427_ net788 vssd1 vssd1
+ vccd1 vccd1 _02428_ sky130_fd_sc_hd__a2111oi_2
XFILLER_53_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09331_ net574 _04165_ _04166_ _04157_ vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__a22o_1
XANTENNA__08277__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09474__A1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11224__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_5_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09262_ net379 _04097_ net312 vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__o21bai_1
X_08213_ datapath.rf.registers\[22\]\[6\] net821 net818 datapath.rf.registers\[7\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03049_ sky130_fd_sc_hd__a22o_1
X_09193_ net557 net577 net546 _02311_ vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__o211a_1
XANTENNA__08029__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07237__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08144_ _02971_ _02976_ _02979_ net782 datapath.rf.registers\[0\]\[8\] vssd1 vssd1
+ vccd1 vccd1 _02980_ sky130_fd_sc_hd__o32a_4
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload140 clknet_leaf_87_clk vssd1 vssd1 vccd1 vccd1 clkload140/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__07657__B net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08075_ _02901_ _02906_ _02910_ vssd1 vssd1 vccd1 vccd1 _02911_ sky130_fd_sc_hd__or3_4
XFILLER_136_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1135_A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10792__B1 _05552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07026_ datapath.rf.registers\[2\]\[30\] net981 net950 vssd1 vssd1 vccd1 vccd1 _01862_
+ sky130_fd_sc_hd__and3_1
Xmax_cap950 net951 vssd1 vssd1 vccd1 vccd1 net950 sky130_fd_sc_hd__clkbuf_2
Xmax_cap972 _01665_ vssd1 vssd1 vccd1 vccd1 net972 sky130_fd_sc_hd__buf_2
XFILLER_0_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout595_A net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14169__RESET_B net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold13 keypad.debounce.debounce\[4\] vssd1 vssd1 vccd1 vccd1 net1361 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold24 screen.register.cFill2 vssd1 vssd1 vccd1 vccd1 net1372 sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ net558 net446 vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__or2_1
Xhold35 screen.controlBus\[9\] vssd1 vssd1 vccd1 vccd1 net1383 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout762_A net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout383_X net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold46 screen.controlBus\[23\] vssd1 vssd1 vccd1 vccd1 net1394 sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ datapath.rf.registers\[2\]\[12\] net745 net686 datapath.rf.registers\[27\]\[12\]
+ _02763_ vssd1 vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__a221o_1
Xhold57 net64 vssd1 vssd1 vccd1 vccd1 net1405 sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 net67 vssd1 vssd1 vccd1 vccd1 net1416 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 net54 vssd1 vssd1 vccd1 vccd1 net1427 sky130_fd_sc_hd__dlygate4sd3_1
X_07859_ datapath.rf.registers\[20\]\[13\] net840 net822 datapath.rf.registers\[22\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1292_X net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08000__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10870_ net898 _05619_ vssd1 vssd1 vccd1 vccd1 _05620_ sky130_fd_sc_hd__nor2_1
XFILLER_44_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09529_ net340 net319 _04017_ vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout815_X net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11134__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12540_ datapath.mulitply_result\[5\] datapath.multiplication_module.multiplicand_i\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06397_ sky130_fd_sc_hd__and2_1
XFILLER_40_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12471_ net166 _05990_ net128 screen.register.currentXbus\[27\] vssd1 vssd1 vccd1
+ vccd1 _00873_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10973__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14210_ clknet_leaf_47_clk datapath.multiplication_module.multiplicand_i_n\[21\]
+ net1172 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07228__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11422_ net265 net2637 net517 vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__mux2_1
XANTENNA__09766__C _04600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14141_ clknet_leaf_8_clk _00898_ net1072 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_115_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10232__C1 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11353_ net271 net2426 net520 vssd1 vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__mux2_1
XANTENNA__08440__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10304_ net1043 _05139_ _05138_ net635 vssd1 vssd1 vccd1 vccd1 _05140_ sky130_fd_sc_hd__a211o_1
XFILLER_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14072_ clknet_leaf_122_clk _00839_ net1216 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11284_ net272 net2218 net524 vssd1 vssd1 vccd1 vccd1 _00332_ sky130_fd_sc_hd__mux2_1
X_13023_ net1919 net178 net393 vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__mux2_1
XFILLER_112_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10235_ net224 _05070_ net1293 vssd1 vssd1 vccd1 vccd1 _05071_ sky130_fd_sc_hd__a21oi_1
XFILLER_152_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08679__A _02523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1011 _05742_ vssd1 vssd1 vccd1 vccd1 net1011 sky130_fd_sc_hd__clkbuf_2
Xfanout1022 _01435_ vssd1 vssd1 vccd1 vccd1 net1022 sky130_fd_sc_hd__buf_2
XANTENNA__11376__Y _05730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1033 _05888_ vssd1 vssd1 vccd1 vccd1 net1033 sky130_fd_sc_hd__buf_2
X_10166_ net899 _04711_ vssd1 vssd1 vccd1 vccd1 _05002_ sky130_fd_sc_hd__or2_4
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1044 _03729_ vssd1 vssd1 vccd1 vccd1 net1044 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08398__B net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1055 net1058 vssd1 vssd1 vccd1 vccd1 net1055 sky130_fd_sc_hd__buf_2
XANTENNA__11309__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1066 net1121 vssd1 vssd1 vccd1 vccd1 net1066 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1077 net1084 vssd1 vssd1 vccd1 vccd1 net1077 sky130_fd_sc_hd__buf_2
X_10097_ datapath.PC\[27\] net1259 vssd1 vssd1 vccd1 vccd1 _04933_ sky130_fd_sc_hd__or2_1
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1088 net1091 vssd1 vssd1 vccd1 vccd1 net1088 sky130_fd_sc_hd__clkbuf_4
Xfanout1099 net1101 vssd1 vssd1 vccd1 vccd1 net1099 sky130_fd_sc_hd__clkbuf_4
X_13925_ clknet_leaf_97_clk _00703_ net1227 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload4_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13856_ clknet_leaf_54_clk _00660_ net1180 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_90_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12807_ net2187 net273 net492 vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__mux2_1
XFILLER_90_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13787_ clknet_leaf_73_clk _00596_ net1243 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08259__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10999_ net2265 net172 net434 vssd1 vssd1 vccd1 vccd1 _00064_ sky130_fd_sc_hd__mux2_1
XANTENNA__11044__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12738_ net1780 net283 net404 vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_106_Left_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12669_ _06502_ _06503_ _06504_ _06498_ vssd1 vssd1 vccd1 vccd1 _06505_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_13_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07219__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14408_ clknet_leaf_59_clk _01113_ net1169 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12383__B net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08967__A0 _02960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14339_ clknet_leaf_139_clk _01044_ net1100 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold505 datapath.rf.registers\[4\]\[31\] vssd1 vssd1 vccd1 vccd1 net1853 sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 datapath.rf.registers\[0\]\[22\] vssd1 vssd1 vccd1 vccd1 net1864 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10774__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold527 datapath.rf.registers\[7\]\[8\] vssd1 vssd1 vccd1 vccd1 net1875 sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 datapath.rf.registers\[6\]\[25\] vssd1 vssd1 vccd1 vccd1 net1886 sky130_fd_sc_hd__dlygate4sd3_1
Xhold549 datapath.rf.registers\[2\]\[28\] vssd1 vssd1 vccd1 vccd1 net1897 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_98_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08900_ datapath.PC\[8\] _03735_ vssd1 vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_115_Left_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09880_ _03755_ _04665_ net224 _04715_ vssd1 vssd1 vccd1 vccd1 _04716_ sky130_fd_sc_hd__or4_1
XANTENNA__09392__A0 _02613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08831_ _03636_ _03638_ vssd1 vssd1 vccd1 vccd1 _03667_ sky130_fd_sc_hd__or2_4
Xhold1205 datapath.rf.registers\[24\]\[9\] vssd1 vssd1 vccd1 vccd1 net2553 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1216 screen.register.currentYbus\[26\] vssd1 vssd1 vccd1 vccd1 net2564 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11219__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1227 datapath.rf.registers\[21\]\[6\] vssd1 vssd1 vccd1 vccd1 net2575 sky130_fd_sc_hd__dlygate4sd3_1
X_08762_ _03482_ _03484_ _03597_ vssd1 vssd1 vccd1 vccd1 _03598_ sky130_fd_sc_hd__and3_1
Xhold1238 datapath.rf.registers\[0\]\[12\] vssd1 vssd1 vccd1 vccd1 net2586 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1249 datapath.rf.registers\[28\]\[6\] vssd1 vssd1 vccd1 vccd1 net2597 sky130_fd_sc_hd__dlygate4sd3_1
X_07713_ datapath.rf.registers\[7\]\[16\] net940 net932 vssd1 vssd1 vccd1 vccd1 _02549_
+ sky130_fd_sc_hd__and3_1
XFILLER_26_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08693_ _02773_ _03442_ vssd1 vssd1 vccd1 vccd1 _03529_ sky130_fd_sc_hd__nor2_1
XFILLER_26_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout176_A _05670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07644_ datapath.rf.registers\[6\]\[18\] net679 _02479_ net786 vssd1 vssd1 vccd1
+ vccd1 _02480_ sky130_fd_sc_hd__a211o_1
XANTENNA__07940__B net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_124_Left_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07575_ datapath.rf.registers\[11\]\[19\] net883 net858 datapath.rf.registers\[24\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__a22o_1
XFILLER_41_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10359__A net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1085_A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09314_ _03577_ _04149_ net580 vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12451__B1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09245_ _01620_ _03506_ net317 _04080_ _04079_ vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_32_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout510_A _05735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10793__S net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout608_A _03608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08771__B net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1252_A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09176_ net338 _04011_ vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__nor2_1
XANTENNA__06572__A datapath.ru.latched_instruction\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11698__A2_N _05885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08958__A0 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08490__C _01800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08127_ datapath.rf.registers\[11\]\[8\] net712 net709 datapath.rf.registers\[10\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1040_X net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08422__A2 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_133_Left_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08058_ datapath.rf.registers\[25\]\[9\] net977 net944 vssd1 vssd1 vccd1 vccd1 _02894_
+ sky130_fd_sc_hd__and3_1
XFILLER_123_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout977_A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput47 net47 vssd1 vssd1 vccd1 vccd1 ADR_O[16] sky130_fd_sc_hd__buf_2
XFILLER_134_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07009_ datapath.rf.registers\[22\]\[31\] net734 net726 datapath.rf.registers\[25\]\[31\]
+ _01842_ vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__a221o_1
XANTENNA__11918__A _02385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput58 net58 vssd1 vssd1 vccd1 vccd1 ADR_O[26] sky130_fd_sc_hd__buf_2
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 ADR_O[7] sky130_fd_sc_hd__buf_2
X_10020_ _04753_ _04802_ vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__xnor2_1
XFILLER_49_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout765_X net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11129__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11971_ _05835_ _06015_ vssd1 vssd1 vccd1 vccd1 _06016_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout932_X net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10968__S net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13710_ clknet_leaf_5_clk _00520_ net1069 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10922_ net186 net2422 net545 vssd1 vssd1 vccd1 vccd1 _00029_ sky130_fd_sc_hd__mux2_1
XANTENNA__07850__B net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14690_ clknet_leaf_152_clk _01395_ net1054 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07697__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06747__A _01585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07161__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13641_ clknet_leaf_61_clk _00451_ net1166 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10853_ net242 net1971 net543 vssd1 vssd1 vccd1 vccd1 _00019_ sky130_fd_sc_hd__mux2_1
X_13572_ clknet_leaf_22_clk _00382_ net1154 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10784_ _01438_ net655 _05545_ _05546_ vssd1 vssd1 vccd1 vccd1 _05547_ sky130_fd_sc_hd__o22a_1
XANTENNA__11796__A2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12523_ datapath.mulitply_result\[1\] datapath.multiplication_module.multiplicand_i\[1\]
+ _06377_ vssd1 vssd1 vccd1 vccd1 _06383_ sky130_fd_sc_hd__a21oi_1
XFILLER_9_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12454_ net166 _05956_ net128 net2656 vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_97_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11405_ net1848 net177 net413 vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__mux2_1
X_12385_ _05942_ net159 vssd1 vssd1 vccd1 vccd1 _06340_ sky130_fd_sc_hd__nor2_1
XANTENNA__09610__A1 _03667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08413__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10435__C _05270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14124_ clknet_leaf_56_clk _00881_ net1159 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11336_ net2069 net186 net415 vssd1 vssd1 vccd1 vccd1 _00381_ sky130_fd_sc_hd__mux2_1
X_14055_ clknet_leaf_95_clk _00822_ net1216 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_140_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11267_ net194 net2127 net418 vssd1 vssd1 vccd1 vccd1 _00316_ sky130_fd_sc_hd__mux2_1
XFILLER_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13006_ net2382 net266 net392 vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__mux2_1
X_10218_ datapath.PC\[29\] _03750_ _05053_ vssd1 vssd1 vccd1 vccd1 _05054_ sky130_fd_sc_hd__a21o_1
X_11198_ net199 net2570 net423 vssd1 vssd1 vccd1 vccd1 _00250_ sky130_fd_sc_hd__mux2_1
XANTENNA__11039__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10149_ _04889_ _04984_ vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_128_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09126__B1 _02217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09677__A1 _03604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13908_ clknet_leaf_43_clk net1362 net1149 vssd1 vssd1 vccd1 vccd1 keypad.debounce.debounce\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07688__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07152__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13839_ clknet_leaf_113_clk _00648_ net1189 vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__dfrtp_1
XFILLER_51_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10039__A2 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07360_ datapath.rf.registers\[5\]\[23\] net945 net932 vssd1 vssd1 vccd1 vccd1 _02196_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_44_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07291_ datapath.rf.registers\[30\]\[25\] net760 net752 datapath.rf.registers\[28\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02127_ sky130_fd_sc_hd__a22o_1
XANTENNA__11502__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09030_ _02147_ _03463_ vssd1 vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__and2b_2
XANTENNA__07860__B1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold302 datapath.rf.registers\[27\]\[3\] vssd1 vssd1 vccd1 vccd1 net1650 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold313 datapath.rf.registers\[14\]\[8\] vssd1 vssd1 vccd1 vccd1 net1661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 datapath.rf.registers\[25\]\[25\] vssd1 vssd1 vccd1 vccd1 net1672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 datapath.rf.registers\[13\]\[18\] vssd1 vssd1 vccd1 vccd1 net1683 sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 datapath.rf.registers\[7\]\[14\] vssd1 vssd1 vccd1 vccd1 net1694 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold357 datapath.rf.registers\[7\]\[3\] vssd1 vssd1 vccd1 vccd1 net1705 sky130_fd_sc_hd__dlygate4sd3_1
Xhold368 datapath.rf.registers\[19\]\[19\] vssd1 vssd1 vccd1 vccd1 net1716 sky130_fd_sc_hd__dlygate4sd3_1
X_09932_ _04766_ _04767_ vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__and2b_1
Xhold379 datapath.rf.registers\[21\]\[23\] vssd1 vssd1 vccd1 vccd1 net1727 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout804 net806 vssd1 vssd1 vccd1 vccd1 net804 sky130_fd_sc_hd__clkbuf_8
Xfanout815 net816 vssd1 vssd1 vccd1 vccd1 net815 sky130_fd_sc_hd__buf_4
XANTENNA__09208__A net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout826 net828 vssd1 vssd1 vccd1 vccd1 net826 sky130_fd_sc_hd__buf_4
XFILLER_131_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout837 _01743_ vssd1 vssd1 vccd1 vccd1 net837 sky130_fd_sc_hd__buf_2
X_09863_ _03443_ _03524_ _04179_ vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__or3b_1
Xfanout848 _01737_ vssd1 vssd1 vccd1 vccd1 net848 sky130_fd_sc_hd__buf_2
XANTENNA_fanout293_A _05541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout859 _01730_ vssd1 vssd1 vccd1 vccd1 net859 sky130_fd_sc_hd__buf_4
XANTENNA__11711__A2 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1002 datapath.rf.registers\[2\]\[26\] vssd1 vssd1 vccd1 vccd1 net2350 sky130_fd_sc_hd__dlygate4sd3_1
X_08814_ _03295_ _03644_ _03648_ vssd1 vssd1 vccd1 vccd1 _03650_ sky130_fd_sc_hd__o21a_1
XFILLER_133_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1013 datapath.rf.registers\[11\]\[2\] vssd1 vssd1 vccd1 vccd1 net2361 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1024 datapath.rf.registers\[28\]\[7\] vssd1 vssd1 vccd1 vccd1 net2372 sky130_fd_sc_hd__dlygate4sd3_1
X_09794_ _03487_ _03489_ _03594_ _04627_ _03485_ vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__a311o_1
Xhold1035 datapath.rf.registers\[24\]\[31\] vssd1 vssd1 vccd1 vccd1 net2383 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07391__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1046 datapath.rf.registers\[1\]\[9\] vssd1 vssd1 vccd1 vccd1 net2394 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1057 datapath.rf.registers\[10\]\[12\] vssd1 vssd1 vccd1 vccd1 net2405 sky130_fd_sc_hd__dlygate4sd3_1
X_08745_ _03513_ _03514_ _03579_ _03511_ vssd1 vssd1 vccd1 vccd1 _03581_ sky130_fd_sc_hd__a31o_1
Xhold1068 datapath.rf.registers\[9\]\[7\] vssd1 vssd1 vccd1 vccd1 net2416 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1079 datapath.rf.registers\[6\]\[11\] vssd1 vssd1 vccd1 vccd1 net2427 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout558_A _03383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08766__B _03601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07679__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07670__B net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08676_ _02466_ _02488_ vssd1 vssd1 vccd1 vccd1 _03512_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_37_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07627_ datapath.rf.registers\[24\]\[18\] net856 net849 datapath.rf.registers\[17\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__a22o_1
XFILLER_53_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07558_ datapath.rf.registers\[7\]\[19\] net941 net934 vssd1 vssd1 vccd1 vccd1 _02394_
+ sky130_fd_sc_hd__and3_1
XFILLER_139_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07489_ datapath.rf.registers\[8\]\[21\] net694 net664 datapath.rf.registers\[15\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__a22o_1
XANTENNA__12508__S net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout513_X net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11412__S net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09228_ net363 _04063_ _04062_ vssd1 vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__o21a_1
XFILLER_108_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10536__B _05281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09159_ net552 net548 net563 vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__a21o_1
XFILLER_5_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08006__B net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07685__X _02521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12170_ net1272 _06192_ _06178_ vssd1 vssd1 vccd1 vccd1 _06193_ sky130_fd_sc_hd__a21oi_1
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout882_X net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11121_ net251 net2500 net427 vssd1 vssd1 vccd1 vccd1 _00176_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_92_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold880 datapath.rf.registers\[1\]\[17\] vssd1 vssd1 vccd1 vccd1 net2228 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold891 datapath.rf.registers\[24\]\[11\] vssd1 vssd1 vccd1 vccd1 net2239 sky130_fd_sc_hd__dlygate4sd3_1
X_11052_ net252 net2363 net431 vssd1 vssd1 vccd1 vccd1 _00112_ sky130_fd_sc_hd__mux2_1
XANTENNA__07564__C net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10003_ _04837_ _04838_ vssd1 vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__nor2_1
XFILLER_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09108__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input21_A DAT_I[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14258__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09659__B2 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13074__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_13_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11954_ _01422_ _05780_ vssd1 vssd1 vccd1 vccd1 _06000_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_123_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10905_ _05649_ vssd1 vssd1 vccd1 vccd1 _05650_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_123_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14673_ clknet_leaf_40_clk _01378_ net1143 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11885_ _02934_ net658 vssd1 vssd1 vccd1 vccd1 _05954_ sky130_fd_sc_hd__nand2_1
XANTENNA__11670__X _05886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13624_ clknet_leaf_7_clk _00434_ net1068 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10836_ datapath.mulitply_result\[15\] net597 net617 vssd1 vssd1 vccd1 vccd1 _05591_
+ sky130_fd_sc_hd__a21o_1
XFILLER_60_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08692__A _02751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10426__C1 _03614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13555_ clknet_leaf_36_clk _00365_ net1129 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08095__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10767_ _05530_ _05531_ vssd1 vssd1 vccd1 vccd1 _05532_ sky130_fd_sc_hd__or2_1
XFILLER_9_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06924__B net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11322__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12506_ net179 net2233 net508 vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__mux2_1
XANTENNA__07842__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13486_ clknet_leaf_1_clk _00296_ net1056 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10698_ net1509 _03227_ net570 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i_n\[3\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA__10446__B _05281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12437_ _05994_ net157 vssd1 vssd1 vccd1 vccd1 _06366_ sky130_fd_sc_hd__nor2_1
X_12368_ net309 _06329_ vssd1 vssd1 vccd1 vccd1 _06330_ sky130_fd_sc_hd__nor2_1
XANTENNA__06940__A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_895 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14107_ clknet_leaf_122_clk _00873_ net1216 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11319_ net1649 net270 net416 vssd1 vssd1 vccd1 vccd1 _00364_ sky130_fd_sc_hd__mux2_1
XANTENNA__07755__B net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12299_ net635 _04856_ vssd1 vssd1 vccd1 vccd1 _06280_ sky130_fd_sc_hd__nor2_1
XFILLER_141_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14038_ clknet_leaf_86_clk _00807_ net1259 vssd1 vssd1 vccd1 vccd1 datapath.PC\[28\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_68_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06860_ datapath.ru.latched_instruction\[14\] _01610_ _01640_ datapath.ru.latched_instruction\[11\]
+ _01695_ vssd1 vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_143_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07373__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06791_ _01585_ net897 vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__nor2_1
XFILLER_55_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08530_ datapath.rf.registers\[19\]\[0\] net855 net803 datapath.rf.registers\[3\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03366_ sky130_fd_sc_hd__a22o_1
XANTENNA__11457__A1 _05582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08461_ _03293_ _03294_ _03262_ vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__a21o_1
X_07412_ datapath.rf.registers\[4\]\[22\] net957 net931 vssd1 vssd1 vccd1 vccd1 _02248_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09698__A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06674__X _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08392_ _03207_ _03226_ net614 vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__mux2_4
X_07343_ datapath.rf.registers\[30\]\[24\] net758 net675 datapath.rf.registers\[29\]\[24\]
+ _02178_ vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__a221o_1
XANTENNA__08086__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11232__S net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout139_A net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07833__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07274_ datapath.rf.registers\[28\]\[25\] net929 net920 vssd1 vssd1 vccd1 vccd1 _02110_
+ sky130_fd_sc_hd__and3_1
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09013_ net647 _03848_ _03770_ vssd1 vssd1 vccd1 vccd1 _03849_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_154_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout306_A net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold110 datapath.multiplication_module.multiplier_i\[14\] vssd1 vssd1 vccd1 vccd1
+ net1458 sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 net98 vssd1 vssd1 vccd1 vccd1 net1469 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold132 net99 vssd1 vssd1 vccd1 vccd1 net1480 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_1_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold143 net85 vssd1 vssd1 vccd1 vccd1 net1491 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13159__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold154 net96 vssd1 vssd1 vccd1 vccd1 net1502 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold165 screen.counter.currentCt\[11\] vssd1 vssd1 vccd1 vccd1 net1513 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07665__B net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold176 net74 vssd1 vssd1 vccd1 vccd1 net1524 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout601 _06170_ vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__buf_2
Xhold187 datapath.rf.registers\[15\]\[17\] vssd1 vssd1 vccd1 vccd1 net1535 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout612 net613 vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__buf_4
XFILLER_104_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold198 datapath.multiplication_module.multiplicand_i\[15\] vssd1 vssd1 vccd1 vccd1
+ net1546 sky130_fd_sc_hd__dlygate4sd3_1
X_09915_ _01613_ _03670_ net604 vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__a21o_1
XANTENNA__13577__RESET_B net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout623 _03722_ vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12998__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout634 net636 vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout675_A net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout645 net646 vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout656 net657 vssd1 vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__buf_2
X_09846_ _04301_ _04677_ _04680_ _04681_ vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__or4_2
Xfanout667 _01834_ vssd1 vssd1 vccd1 vccd1 net667 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08777__A _03601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout678 _01829_ vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout689 net690 vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__clkbuf_8
XFILLER_100_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11915__B screen.counter.ack vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09777_ net347 _04541_ vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__or2_1
XANTENNA__12299__A net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout842_A net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout463_X net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06989_ net991 _01637_ _01647_ _01666_ vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__and4_2
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11407__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08728_ _03562_ _03563_ _03540_ vssd1 vssd1 vccd1 vccd1 _03564_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_1_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07116__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08659_ _02169_ _02190_ vssd1 vssd1 vccd1 vccd1 _03495_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout630_X net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10120__A1 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout728_X net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11670_ _01405_ _05291_ _05883_ _05290_ vssd1 vssd1 vccd1 vccd1 _05886_ sky130_fd_sc_hd__a22o_2
X_10621_ _05430_ _05438_ _05428_ vssd1 vssd1 vccd1 vccd1 _05441_ sky130_fd_sc_hd__a21oi_1
XFILLER_139_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08077__B1 _02911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11142__S net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13340_ clknet_leaf_7_clk _00150_ net1071 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10552_ _05376_ _05377_ _05378_ vssd1 vssd1 vccd1 vccd1 _05379_ sky130_fd_sc_hd__and3_1
XANTENNA__07559__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13271_ clknet_leaf_124_clk _00081_ net1208 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10981__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10483_ _05311_ _05312_ vssd1 vssd1 vccd1 vccd1 _05313_ sky130_fd_sc_hd__nor2_1
X_12222_ screen.counter.currentCt\[11\] _06223_ net602 vssd1 vssd1 vccd1 vccd1 _06225_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__12258__A2_N _05002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07052__A1 datapath.rf.registers\[0\]\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13069__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12153_ net1278 _06181_ _06182_ _06170_ vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__a22o_1
X_11104_ net170 net2033 net534 vssd1 vssd1 vccd1 vccd1 _00161_ sky130_fd_sc_hd__mux2_1
X_12084_ screen.register.currentYbus\[30\] _05757_ _06019_ screen.register.currentYbus\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06123_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_9_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11035_ net170 net1945 net538 vssd1 vssd1 vccd1 vccd1 _00097_ sky130_fd_sc_hd__mux2_1
XFILLER_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08687__A _02660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06919__B net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11317__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12986_ net202 net2009 net478 vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__mux2_1
XANTENNA__07107__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11937_ net136 _05988_ _05987_ vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__o21ai_1
XFILLER_60_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14656_ clknet_leaf_134_clk _01361_ net1104 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_11868_ net137 _05942_ _05941_ vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06935__A _01630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10819_ net1266 datapath.PC\[13\] _05565_ vssd1 vssd1 vccd1 vccd1 _05576_ sky130_fd_sc_hd__and3_1
X_13607_ clknet_leaf_137_clk _00417_ net1089 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11799_ datapath.ru.latched_instruction\[5\] net336 net316 _01441_ vssd1 vssd1 vccd1
+ vccd1 _00665_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_41_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08607__A2 _02750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09804__A1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14587_ clknet_leaf_39_clk _01292_ net1145 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11052__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13538_ clknet_leaf_151_clk _00348_ net1052 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
Xteam_04_1309 vssd1 vssd1 vccd1 vccd1 team_04_1309/HI gpio_oeb[18] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_136_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13469_ clknet_leaf_146_clk _00279_ net1088 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12391__B net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08240__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07594__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07961_ datapath.rf.registers\[24\]\[11\] net858 net812 datapath.rf.registers\[13\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__a22o_1
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09700_ _04519_ _04520_ _04535_ net605 vssd1 vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__a211o_1
X_06912_ net981 net919 vssd1 vssd1 vccd1 vccd1 _01748_ sky130_fd_sc_hd__and2_1
X_07892_ datapath.rf.registers\[28\]\[12\] net930 _01744_ vssd1 vssd1 vccd1 vccd1
+ _02728_ sky130_fd_sc_hd__and3_1
XANTENNA__08597__A _02960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07346__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09631_ net575 _04460_ _04461_ _04466_ vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__o2bb2a_1
X_06843_ _01413_ _01678_ vssd1 vssd1 vccd1 vccd1 _01679_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_52_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11227__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09562_ _03555_ _03556_ vssd1 vssd1 vccd1 vccd1 _04398_ sky130_fd_sc_hd__xnor2_1
X_06774_ _01513_ _01568_ net1030 datapath.ru.latched_instruction\[14\] vssd1 vssd1
+ vccd1 vccd1 _01611_ sky130_fd_sc_hd__a2bb2o_2
X_08513_ datapath.rf.registers\[24\]\[1\] net963 net911 net908 vssd1 vssd1 vccd1 vccd1
+ _03349_ sky130_fd_sc_hd__and4_1
X_09493_ _01603_ _04328_ _04315_ _03611_ _03600_ vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10919__X _05662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08444_ datapath.rf.registers\[14\]\[2\] net777 _03267_ _03268_ _03270_ vssd1 vssd1
+ vccd1 vccd1 _03280_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_156_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08375_ datapath.rf.registers\[7\]\[3\] net673 net662 datapath.rf.registers\[5\]\[3\]
+ _03210_ vssd1 vssd1 vccd1 vccd1 _03211_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout423_A net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07326_ datapath.rf.registers\[25\]\[24\] net842 net802 datapath.rf.registers\[3\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__a22o_1
XANTENNA__10405__A2 _03384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07806__B1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09875__B _04710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07257_ _02092_ vssd1 vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_59_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout309_X net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13758__RESET_B net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07188_ _02014_ _02016_ _02019_ _02023_ vssd1 vssd1 vccd1 vccd1 _02024_ sky130_fd_sc_hd__or4_1
XANTENNA__08124__X _02960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08231__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1120_X net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07585__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout580_X net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout420 _05722_ vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_6_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout431 net433 vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__buf_4
XANTENNA__08778__Y _03614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout678_X net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08003__C net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout442 net443 vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__clkbuf_4
Xfanout453 _03658_ vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__clkbuf_2
Xfanout464 _03104_ vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07337__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout475 net477 vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__clkbuf_8
Xfanout486 _06552_ vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__buf_6
XFILLER_101_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10877__C1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09731__B1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09829_ _03756_ _04626_ _04645_ _04664_ vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__nor4_1
Xfanout497 _06550_ vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout845_X net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11137__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12840_ net270 net2387 net488 vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__mux2_1
XFILLER_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ net283 net1928 net496 vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_147_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_147_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09495__C1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10976__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ net8 net1033 net1023 net2607 vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__o22a_1
XANTENNA__06848__A1 datapath.ru.latched_instruction\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14510_ clknet_leaf_5_clk _01215_ net1069 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11653_ button\[0\] _05874_ vssd1 vssd1 vccd1 vccd1 _05876_ sky130_fd_sc_hd__and2_1
X_14441_ clknet_leaf_91_clk _01146_ net1241 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_42_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09247__C1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10604_ screen.register.currentYbus\[17\] screen.register.currentYbus\[16\] screen.register.currentYbus\[19\]
+ _05424_ vssd1 vssd1 vccd1 vccd1 _05425_ sky130_fd_sc_hd__or4_1
X_14372_ clknet_leaf_22_clk _01077_ net1157 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11584_ net1272 screen.counter.ct\[19\] screen.counter.ct\[18\] net1271 vssd1 vssd1
+ vccd1 vccd1 _05808_ sky130_fd_sc_hd__or4bb_1
X_13323_ clknet_leaf_55_clk _00133_ net1173 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10535_ net656 vssd1 vssd1 vccd1 vccd1 screen.counter.ack sky130_fd_sc_hd__inv_2
XANTENNA__08470__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06761__Y _01598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13254_ clknet_leaf_17_clk _00064_ net1107 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10466_ screen.counter.ct\[18\] screen.counter.ct\[19\] vssd1 vssd1 vccd1 vccd1 _05296_
+ sky130_fd_sc_hd__or2_1
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12205_ screen.counter.currentCt\[5\] screen.counter.currentCt\[4\] _06210_ vssd1
+ vssd1 vccd1 vccd1 _06214_ sky130_fd_sc_hd__and3_1
XFILLER_142_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08222__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13185_ net1864 vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08969__X _03805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10397_ net326 _05230_ _05232_ vssd1 vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__a21oi_1
XFILLER_124_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07576__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12136_ net1012 net567 screen.counter.ct\[0\] vssd1 vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__mux2_1
XANTENNA__07592__Y _02428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12067_ screen.register.currentYbus\[13\] _05776_ net999 screen.register.currentXbus\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06107_ sky130_fd_sc_hd__a22o_1
XFILLER_111_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07328__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12321__A2 _06254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11018_ net251 net2461 net539 vssd1 vssd1 vccd1 vccd1 _00080_ sky130_fd_sc_hd__mux2_1
XANTENNA__10332__A1 _04239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11047__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08289__A0 _03123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_138_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_138_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09486__C1 _03204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08828__A2 _03661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12969_ net282 net2085 net480 vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__mux2_1
XFILLER_33_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06839__B2 datapath.ru.latched_instruction\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14639_ clknet_leaf_26_clk _01344_ net1137 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10187__A _04146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12388__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08160_ datapath.rf.registers\[16\]\[7\] net862 net838 datapath.rf.registers\[26\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02996_ sky130_fd_sc_hd__a22o_1
XFILLER_119_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08880__A _01614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07111_ _01942_ _01944_ _01946_ vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__or3_1
XANTENNA__08461__B1 _03262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08091_ datapath.rf.registers\[4\]\[9\] net716 net681 datapath.rf.registers\[6\]\[9\]
+ _02926_ vssd1 vssd1 vccd1 vccd1 _02927_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_151_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload30 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 clkload30/Y sky130_fd_sc_hd__clkinv_4
Xclkload41 clknet_leaf_143_clk vssd1 vssd1 vccd1 vccd1 clkload41/Y sky130_fd_sc_hd__inv_8
X_07042_ datapath.rf.registers\[6\]\[30\] net825 net823 datapath.rf.registers\[22\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__a22o_1
XANTENNA__13851__RESET_B net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload52 clknet_leaf_133_clk vssd1 vssd1 vccd1 vccd1 clkload52/X sky130_fd_sc_hd__clkbuf_8
Xclkload63 clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 clkload63/Y sky130_fd_sc_hd__bufinv_16
Xclkload74 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 clkload74/Y sky130_fd_sc_hd__bufinv_16
Xclkload85 clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 clkload85/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__08213__B1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload96 clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 clkload96/Y sky130_fd_sc_hd__inv_8
XFILLER_115_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_1_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08993_ _03469_ _03828_ vssd1 vssd1 vccd1 vccd1 _03829_ sky130_fd_sc_hd__xor2_1
XANTENNA__07943__B net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07944_ datapath.rf.registers\[3\]\[11\] net985 net927 vssd1 vssd1 vccd1 vccd1 _02780_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_149_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07319__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12312__A2 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07875_ datapath.rf.registers\[1\]\[13\] net763 net691 datapath.rf.registers\[13\]\[13\]
+ _02710_ vssd1 vssd1 vccd1 vccd1 _02711_ sky130_fd_sc_hd__a221o_1
XANTENNA__07662__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09614_ net644 _04448_ _04449_ _04446_ vssd1 vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__or4b_1
X_06826_ _01652_ _01653_ _01658_ _01661_ vssd1 vssd1 vccd1 vccd1 _01662_ sky130_fd_sc_hd__or4_1
XANTENNA__12076__A1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09545_ net366 _04376_ net373 vssd1 vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_129_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_129_clk
+ sky130_fd_sc_hd__clkbuf_8
X_06757_ _01497_ net1017 net994 net1030 datapath.ru.latched_instruction\[29\] vssd1
+ vssd1 vccd1 vccd1 _01594_ sky130_fd_sc_hd__a32oi_4
XANTENNA_fanout161_X net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout540_A net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout638_A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09476_ net459 _04307_ _04308_ net354 vssd1 vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__a211o_1
X_06688_ net1286 net1281 mmio.memload_or_instruction\[23\] vssd1 vssd1 vccd1 vccd1
+ _01527_ sky130_fd_sc_hd__nor3b_2
XANTENNA__11823__B2 datapath.ru.latched_instruction\[29\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_51_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07023__X _01859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08427_ datapath.rf.registers\[0\]\[2\] net868 _03261_ vssd1 vssd1 vccd1 vccd1 _03263_
+ sky130_fd_sc_hd__o21ai_4
XANTENNA_fanout426_X net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout805_A net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08358_ datapath.rf.registers\[11\]\[3\] net884 _03176_ _03180_ _03187_ vssd1 vssd1
+ vccd1 vccd1 _03194_ sky130_fd_sc_hd__a2111o_1
Xclkload2 clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clkload2/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__13939__RESET_B net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07309_ datapath.rf.registers\[0\]\[25\] net783 _02139_ _02144_ vssd1 vssd1 vccd1
+ vccd1 _02145_ sky130_fd_sc_hd__o22a_4
XANTENNA__08452__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08289_ _03123_ _03124_ net611 vssd1 vssd1 vccd1 vccd1 _03125_ sky130_fd_sc_hd__mux2_1
XFILLER_153_916 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11420__S net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10320_ net224 _05155_ net1293 vssd1 vssd1 vccd1 vccd1 _05156_ sky130_fd_sc_hd__a21o_1
XFILLER_4_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout795_X net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10251_ datapath.PC\[11\] _04300_ net467 vssd1 vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__mux2_1
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10182_ net226 _05017_ net1295 vssd1 vssd1 vccd1 vccd1 _05018_ sky130_fd_sc_hd__a21o_1
XFILLER_133_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1204 net1262 vssd1 vssd1 vccd1 vccd1 net1204 sky130_fd_sc_hd__clkbuf_4
Xfanout1215 net1216 vssd1 vssd1 vccd1 vccd1 net1215 sky130_fd_sc_hd__buf_2
Xfanout1226 net1227 vssd1 vssd1 vccd1 vccd1 net1226 sky130_fd_sc_hd__clkbuf_4
Xfanout1237 net1238 vssd1 vssd1 vccd1 vccd1 net1237 sky130_fd_sc_hd__clkbuf_2
Xfanout250 _05592_ vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__clkbuf_2
Xfanout1248 net1249 vssd1 vssd1 vccd1 vccd1 net1248 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_89_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12303__A2 _06254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1259 net1260 vssd1 vssd1 vccd1 vccd1 net1259 sky130_fd_sc_hd__buf_2
Xfanout261 _05703_ vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_89_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09704__B1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout272 _05564_ vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__clkbuf_2
X_13941_ clknet_leaf_95_clk _00719_ net1226 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[25\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout283 net285 vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout294 net297 vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__clkbuf_2
X_13872_ clknet_leaf_51_clk _00676_ net1182 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[16\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07191__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12823_ net2424 net192 net490 vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__mux2_1
XANTENNA__06756__Y _01593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13082__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10078__B1 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_141_Right_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12754_ net1941 net203 net402 vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__mux2_1
XFILLER_91_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09483__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11705_ net1291 mmio.wishbone.prev_BUSY_O net1034 vssd1 vssd1 vccd1 vccd1 _05889_
+ sky130_fd_sc_hd__and3b_1
X_12685_ datapath.mulitply_result\[29\] datapath.multiplication_module.multiplicand_i\[29\]
+ vssd1 vssd1 vccd1 vccd1 _06518_ sky130_fd_sc_hd__and2_1
XANTENNA__07868__X _02704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11636_ _05820_ _05852_ _05859_ _05758_ _05858_ vssd1 vssd1 vccd1 vccd1 _05860_ sky130_fd_sc_hd__o221a_1
X_14424_ clknet_leaf_3_clk _01129_ net1076 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06772__X _01609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11567_ net1008 _05775_ vssd1 vssd1 vccd1 vccd1 _05791_ sky130_fd_sc_hd__or2_1
X_14355_ clknet_leaf_34_clk _01060_ net1128 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08443__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11330__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06932__B net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10518_ _05335_ _05342_ _05346_ _05347_ _05341_ vssd1 vssd1 vccd1 vccd1 _05348_ sky130_fd_sc_hd__o2111a_1
X_13306_ clknet_leaf_14_clk _00116_ net1102 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold709 datapath.mulitply_result\[29\] vssd1 vssd1 vccd1 vccd1 net2057 sky130_fd_sc_hd__dlygate4sd3_1
X_14286_ clknet_leaf_2_clk _00991_ net1063 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_144_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11498_ net232 net2006 net512 vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__mux2_1
X_13237_ clknet_leaf_129_clk _00047_ net1117 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10449_ _05204_ _05284_ vssd1 vssd1 vccd1 vccd1 _05285_ sky130_fd_sc_hd__or2_2
XANTENNA__07549__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13168_ net2404 vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_41_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12119_ net1276 net1274 _06155_ vssd1 vssd1 vccd1 vccd1 _06156_ sky130_fd_sc_hd__and3_1
XFILLER_2_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13099_ net300 net2150 net472 vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__mux2_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08578__C _01816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07660_ datapath.rf.registers\[14\]\[17\] net982 net919 vssd1 vssd1 vccd1 vccd1 _02496_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07182__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_56_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06611_ mmio.key_data\[4\] net1048 _01448_ vssd1 vssd1 vccd1 vccd1 _01450_ sky130_fd_sc_hd__o21a_1
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07591_ datapath.rf.registers\[3\]\[19\] net772 net716 datapath.rf.registers\[4\]\[19\]
+ _02420_ vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__a221o_1
XANTENNA__11505__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09330_ net648 _04165_ net438 vssd1 vssd1 vccd1 vccd1 _04166_ sky130_fd_sc_hd__a21o_1
XFILLER_34_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09261_ _04095_ _04096_ vssd1 vssd1 vccd1 vccd1 _04097_ sky130_fd_sc_hd__nor2_1
X_08212_ datapath.rf.registers\[20\]\[6\] net839 net813 datapath.rf.registers\[23\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03048_ sky130_fd_sc_hd__a22o_1
XFILLER_138_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09192_ net375 _03873_ _03627_ vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_114_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08143_ _02962_ _02967_ _02977_ _02978_ vssd1 vssd1 vccd1 vccd1 _02979_ sky130_fd_sc_hd__or4_1
XANTENNA__07938__B net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07788__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload130 clknet_leaf_92_clk vssd1 vssd1 vccd1 vccd1 clkload130/Y sky130_fd_sc_hd__clkinv_8
X_08074_ _02907_ _02908_ _02909_ vssd1 vssd1 vccd1 vccd1 _02910_ sky130_fd_sc_hd__or3_1
Xclkload141 clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 clkload141/Y sky130_fd_sc_hd__inv_6
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10364__B _05116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07657__C net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07025_ datapath.rf.registers\[25\]\[30\] net973 net944 vssd1 vssd1 vccd1 vccd1 _01861_
+ sky130_fd_sc_hd__and3_1
XFILLER_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_129_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1030_A net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout490_A _06551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11741__B1 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold14 keypad.debounce.debounce\[9\] vssd1 vssd1 vccd1 vccd1 net1362 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08976_ net448 _03809_ vssd1 vssd1 vccd1 vccd1 _03812_ sky130_fd_sc_hd__or2_1
XFILLER_152_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold25 screen.register.xFill2 vssd1 vssd1 vccd1 vccd1 net1373 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 screen.controlBus\[15\] vssd1 vssd1 vccd1 vccd1 net1384 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold47 datapath.multiplication_module.multiplier_i\[6\] vssd1 vssd1 vccd1 vccd1 net1395
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07960__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold58 screen.controlBus\[12\] vssd1 vssd1 vccd1 vccd1 net1406 sky130_fd_sc_hd__dlygate4sd3_1
X_07927_ datapath.rf.registers\[30\]\[12\] net761 net753 datapath.rf.registers\[28\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02763_ sky130_fd_sc_hd__a22o_1
Xhold69 net71 vssd1 vssd1 vccd1 vccd1 net1417 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout755_A net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07858_ datapath.rf.registers\[6\]\[13\] net825 net820 datapath.rf.registers\[5\]\[13\]
+ _02686_ vssd1 vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__a221o_1
XFILLER_84_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07173__B1 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06809_ datapath.ru.latched_instruction\[23\] _01527_ net1015 vssd1 vssd1 vccd1 vccd1
+ _01645_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_67_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07789_ _02623_ _02624_ vssd1 vssd1 vccd1 vccd1 _02625_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout922_A net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout543_X net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11415__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09528_ net345 _04362_ _04363_ _04357_ _01607_ vssd1 vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__a311o_1
XFILLER_40_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10539__B net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout710_X net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09459_ _03531_ net625 _03718_ _03532_ vssd1 vssd1 vccd1 vccd1 _04295_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout808_X net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12470_ net166 _05988_ net128 screen.register.currentXbus\[26\] vssd1 vssd1 vccd1
+ vccd1 _00872_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_131_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11421_ net268 net2239 net516 vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__mux2_1
XFILLER_138_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07848__B net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11150__S net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07779__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14140_ clknet_leaf_36_clk _00897_ net1136 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11352_ net276 net2632 net520 vssd1 vssd1 vccd1 vccd1 _00395_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_115_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07567__C net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10303_ net1266 _03738_ vssd1 vssd1 vccd1 vccd1 _05139_ sky130_fd_sc_hd__xnor2_1
X_14071_ clknet_leaf_122_clk _00838_ net1214 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_152_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11283_ net274 net2323 net524 vssd1 vssd1 vccd1 vccd1 _00331_ sky130_fd_sc_hd__mux2_1
X_13022_ net1726 net188 net390 vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__mux2_1
X_10234_ _04893_ _05069_ vssd1 vssd1 vccd1 vccd1 _05070_ sky130_fd_sc_hd__or2_1
XFILLER_10_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1001 _05332_ vssd1 vssd1 vccd1 vccd1 net1001 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13077__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10165_ _04864_ _04865_ vssd1 vssd1 vccd1 vccd1 _05001_ sky130_fd_sc_hd__xnor2_1
Xfanout1023 _05890_ vssd1 vssd1 vccd1 vccd1 net1023 sky130_fd_sc_hd__buf_2
XFILLER_86_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1034 _05888_ vssd1 vssd1 vccd1 vccd1 net1034 sky130_fd_sc_hd__buf_2
Xfanout1056 net1058 vssd1 vssd1 vccd1 vccd1 net1056 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08398__C net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12288__A1 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10096_ net1258 _04929_ _04931_ _04920_ vssd1 vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__a31o_1
Xfanout1067 net1068 vssd1 vssd1 vccd1 vccd1 net1067 sky130_fd_sc_hd__clkbuf_4
Xfanout1078 net1084 vssd1 vssd1 vccd1 vccd1 net1078 sky130_fd_sc_hd__clkbuf_4
Xfanout1089 net1091 vssd1 vssd1 vccd1 vccd1 net1089 sky130_fd_sc_hd__clkbuf_4
X_13924_ clknet_leaf_96_clk _00702_ net1227 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_63_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08695__A _02805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07703__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13855_ clknet_leaf_50_clk net2433 net1176 vssd1 vssd1 vccd1 vccd1 keypad.apps.app_c\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06911__B1 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11325__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12806_ net2394 net274 net492 vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__mux2_1
X_13786_ clknet_leaf_73_clk _00595_ net1243 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10998_ net2421 net183 net434 vssd1 vssd1 vccd1 vccd1 _00063_ sky130_fd_sc_hd__mux2_1
XFILLER_43_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12737_ net1811 net292 net402 vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__mux2_1
XFILLER_43_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12668_ _06497_ _06499_ vssd1 vssd1 vccd1 vccd1 _06504_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_13_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14407_ clknet_leaf_142_clk _01112_ net1093 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06690__A2 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11619_ _05752_ _05842_ vssd1 vssd1 vccd1 vccd1 _05843_ sky130_fd_sc_hd__and2_1
XANTENNA__07758__B net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08416__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06662__B _01500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11060__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12599_ datapath.mulitply_result\[15\] datapath.multiplication_module.multiplicand_i\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06446_ sky130_fd_sc_hd__and2_1
XFILLER_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08967__A1 _03008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14338_ clknet_leaf_152_clk _01043_ net1054 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold506 datapath.rf.registers\[16\]\[25\] vssd1 vssd1 vccd1 vccd1 net1854 sky130_fd_sc_hd__dlygate4sd3_1
Xhold517 datapath.rf.registers\[22\]\[21\] vssd1 vssd1 vccd1 vccd1 net1865 sky130_fd_sc_hd__dlygate4sd3_1
Xhold528 datapath.rf.registers\[15\]\[8\] vssd1 vssd1 vccd1 vccd1 net1876 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold539 datapath.rf.registers\[6\]\[21\] vssd1 vssd1 vccd1 vccd1 net1887 sky130_fd_sc_hd__dlygate4sd3_1
X_14269_ clknet_leaf_143_clk _00974_ net1085 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_143_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09392__A1 _02661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08830_ _03636_ _03638_ vssd1 vssd1 vccd1 vccd1 _03666_ sky130_fd_sc_hd__nor2_1
Xhold1206 datapath.rf.registers\[11\]\[12\] vssd1 vssd1 vccd1 vccd1 net2554 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1217 datapath.rf.registers\[2\]\[7\] vssd1 vssd1 vccd1 vccd1 net2565 sky130_fd_sc_hd__dlygate4sd3_1
X_08761_ _03487_ _03489_ _03594_ _03485_ _03483_ vssd1 vssd1 vccd1 vccd1 _03597_ sky130_fd_sc_hd__a311o_1
Xhold1228 datapath.rf.registers\[17\]\[29\] vssd1 vssd1 vccd1 vccd1 net2576 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1239 screen.register.currentYbus\[9\] vssd1 vssd1 vccd1 vccd1 net2587 sky130_fd_sc_hd__dlygate4sd3_1
X_07712_ datapath.rf.registers\[6\]\[16\] net954 net931 vssd1 vssd1 vccd1 vccd1 _02548_
+ sky130_fd_sc_hd__and3_1
XFILLER_66_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08692_ _02751_ _02772_ vssd1 vssd1 vccd1 vccd1 _03528_ sky130_fd_sc_hd__nand2_1
XANTENNA__07155__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09695__A2 _03718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07643_ datapath.rf.registers\[14\]\[18\] net774 net694 datapath.rf.registers\[8\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__a22o_1
XFILLER_54_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07940__C _01712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11235__S net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07574_ net874 _02407_ _02408_ _02409_ vssd1 vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__or4_1
XFILLER_22_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09313_ _03521_ _03576_ _03518_ vssd1 vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_60_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1078_A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09244_ net337 _03816_ vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_62_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_888 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08771__C _03601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09175_ _04008_ _04010_ net341 vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__mux2_1
XANTENNA__07668__B net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout503_A net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1245_A net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08958__A1 _02613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08126_ datapath.rf.registers\[25\]\[8\] net728 net689 datapath.rf.registers\[31\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__a22o_1
XFILLER_119_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08057_ datapath.rf.registers\[24\]\[9\] _01712_ net929 vssd1 vssd1 vccd1 vccd1 _02893_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07630__B2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1033_X net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07008_ datapath.rf.registers\[16\]\[31\] net738 net730 datapath.rf.registers\[19\]\[31\]
+ _01843_ vssd1 vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__a221o_1
XANTENNA__11477__Y _05735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput48 net48 vssd1 vssd1 vccd1 vccd1 ADR_O[17] sky130_fd_sc_hd__buf_2
Xoutput59 net59 vssd1 vssd1 vccd1 vccd1 ADR_O[27] sky130_fd_sc_hd__buf_2
XANTENNA_fanout872_A _01723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout493_X net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08499__B net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08186__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_866 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07394__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07933__A2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout660_X net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08959_ _03794_ vssd1 vssd1 vccd1 vccd1 _03795_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout758_X net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11970_ _05861_ _05868_ _05819_ vssd1 vssd1 vccd1 vccd1 _06015_ sky130_fd_sc_hd__o21ai_1
XFILLER_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07146__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11653__B _05874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10921_ _01479_ net622 _05662_ _05663_ vssd1 vssd1 vccd1 vccd1 _05664_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_29_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07850__C net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout925_X net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11145__S net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10852_ _01451_ _05604_ net653 vssd1 vssd1 vccd1 vccd1 _05605_ sky130_fd_sc_hd__mux2_2
X_13640_ clknet_leaf_91_clk _00450_ net1233 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13571_ clknet_leaf_121_clk _00381_ net1192 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10984__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10783_ datapath.mulitply_result\[7\] net598 net620 vssd1 vssd1 vccd1 vccd1 _05546_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__10837__X _05592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_51_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08110__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12522_ _06380_ _06381_ vssd1 vssd1 vccd1 vccd1 _06382_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_10_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12453_ net167 _05954_ net129 screen.register.currentXbus\[9\] vssd1 vssd1 vccd1
+ vccd1 _00855_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_97_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11404_ net2304 net186 net411 vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12384_ net2055 net133 _06339_ vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__a21o_1
X_11335_ net1745 net193 net414 vssd1 vssd1 vccd1 vccd1 _00380_ sky130_fd_sc_hd__mux2_1
XFILLER_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14123_ clknet_leaf_59_clk _00880_ net1170 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_126_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14054_ clknet_4_11_0_clk _00821_ net1222 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_11266_ net198 net2108 net420 vssd1 vssd1 vccd1 vccd1 _00315_ sky130_fd_sc_hd__mux2_1
XFILLER_140_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08177__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13005_ net2441 net270 net392 vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__mux2_1
X_10217_ net1044 _03751_ vssd1 vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__nand2_1
X_11197_ net206 net2468 net422 vssd1 vssd1 vccd1 vccd1 _00249_ sky130_fd_sc_hd__mux2_1
XANTENNA__08202__B net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07385__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07924__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10148_ _04885_ _04888_ vssd1 vssd1 vccd1 vccd1 _04984_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_128_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10079_ _04911_ _04912_ _04914_ net637 vssd1 vssd1 vccd1 vccd1 _04915_ sky130_fd_sc_hd__a211oi_1
XFILLER_36_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13907_ clknet_leaf_43_clk net1357 net1149 vssd1 vssd1 vccd1 vccd1 keypad.debounce.debounce\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11055__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13838_ clknet_leaf_115_clk _00647_ net1195 vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__dfrtp_1
X_13769_ clknet_leaf_81_clk _00578_ net1255 vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_42_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_43_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10444__B1 net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07290_ datapath.rf.registers\[0\]\[25\] net868 _02124_ vssd1 vssd1 vccd1 vccd1 _02126_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06960__X _01796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold303 datapath.rf.registers\[20\]\[22\] vssd1 vssd1 vccd1 vccd1 net1651 sky130_fd_sc_hd__dlygate4sd3_1
Xhold314 datapath.rf.registers\[19\]\[17\] vssd1 vssd1 vccd1 vccd1 net1662 sky130_fd_sc_hd__dlygate4sd3_1
Xhold325 datapath.rf.registers\[1\]\[16\] vssd1 vssd1 vccd1 vccd1 net1673 sky130_fd_sc_hd__dlygate4sd3_1
Xhold336 datapath.rf.registers\[6\]\[12\] vssd1 vssd1 vccd1 vccd1 net1684 sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 datapath.rf.registers\[22\]\[28\] vssd1 vssd1 vccd1 vccd1 net1695 sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 datapath.rf.registers\[31\]\[10\] vssd1 vssd1 vccd1 vccd1 net1706 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold369 datapath.rf.registers\[30\]\[7\] vssd1 vssd1 vccd1 vccd1 net1717 sky130_fd_sc_hd__dlygate4sd3_1
X_09931_ datapath.PC\[7\] _03029_ vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__or2_1
Xfanout805 net806 vssd1 vssd1 vccd1 vccd1 net805 sky130_fd_sc_hd__clkbuf_4
Xfanout816 _01759_ vssd1 vssd1 vccd1 vccd1 net816 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08168__A2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout827 net828 vssd1 vssd1 vccd1 vccd1 net827 sky130_fd_sc_hd__clkbuf_4
X_09862_ _02826_ _04697_ _04673_ vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__a21o_1
Xfanout838 _01743_ vssd1 vssd1 vccd1 vccd1 net838 sky130_fd_sc_hd__buf_4
XFILLER_140_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07376__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout849 _01735_ vssd1 vssd1 vccd1 vccd1 net849 sky130_fd_sc_hd__buf_4
Xhold1003 datapath.rf.registers\[9\]\[27\] vssd1 vssd1 vccd1 vccd1 net2351 sky130_fd_sc_hd__dlygate4sd3_1
X_08813_ _03295_ _03644_ _03648_ vssd1 vssd1 vccd1 vccd1 _03649_ sky130_fd_sc_hd__o21ai_1
XFILLER_133_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1014 datapath.rf.registers\[14\]\[31\] vssd1 vssd1 vccd1 vccd1 net2362 sky130_fd_sc_hd__dlygate4sd3_1
X_09793_ _03474_ _04627_ vssd1 vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__xnor2_2
Xhold1025 mmio.memload_or_instruction\[10\] vssd1 vssd1 vccd1 vccd1 net2373 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_86_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1036 datapath.rf.registers\[19\]\[16\] vssd1 vssd1 vccd1 vccd1 net2384 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1047 datapath.rf.registers\[8\]\[13\] vssd1 vssd1 vccd1 vccd1 net2395 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1058 datapath.rf.registers\[27\]\[30\] vssd1 vssd1 vccd1 vccd1 net2406 sky130_fd_sc_hd__dlygate4sd3_1
X_08744_ _03514_ _03579_ vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__nand2_1
Xhold1069 datapath.rf.registers\[11\]\[23\] vssd1 vssd1 vccd1 vccd1 net2417 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07670__C net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08675_ _03510_ vssd1 vssd1 vccd1 vccd1 _03511_ sky130_fd_sc_hd__inv_2
XANTENNA__08876__A0 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10132__C1 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07626_ datapath.rf.registers\[19\]\[18\] net853 net793 datapath.rf.registers\[31\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__a22o_1
XFILLER_81_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07557_ datapath.rf.registers\[4\]\[19\] net959 net935 vssd1 vssd1 vccd1 vccd1 _02393_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout718_A net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_33_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_8
X_07488_ datapath.rf.registers\[4\]\[21\] net714 net679 datapath.rf.registers\[6\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02324_ sky130_fd_sc_hd__a22o_1
XANTENNA__07300__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09227_ _02312_ _02365_ net443 vssd1 vssd1 vccd1 vccd1 _04063_ sky130_fd_sc_hd__mux2_1
XFILLER_10_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout506_X net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1248_X net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09158_ _02217_ net553 net549 vssd1 vssd1 vccd1 vccd1 _03994_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_79_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08006__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08109_ datapath.rf.registers\[1\]\[8\] net848 net831 datapath.rf.registers\[14\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__a22o_1
X_09089_ net330 _03924_ net311 vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__a21oi_1
XFILLER_107_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11120_ net257 net2458 net427 vssd1 vssd1 vccd1 vccd1 _00175_ sky130_fd_sc_hd__mux2_1
Xhold870 datapath.rf.registers\[25\]\[10\] vssd1 vssd1 vccd1 vccd1 net2218 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout875_X net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold881 datapath.rf.registers\[30\]\[17\] vssd1 vssd1 vccd1 vccd1 net2229 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08159__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14153__RESET_B net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold892 datapath.rf.registers\[21\]\[29\] vssd1 vssd1 vccd1 vccd1 net2240 sky130_fd_sc_hd__dlygate4sd3_1
X_11051_ net254 net2395 net431 vssd1 vssd1 vccd1 vccd1 _00111_ sky130_fd_sc_hd__mux2_1
XANTENNA__07367__B1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07906__A2 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10002_ _04778_ _04787_ vssd1 vssd1 vccd1 vccd1 _04838_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10979__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10371__C1 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07119__B1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input14_A DAT_I[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11953_ _05349_ net996 vssd1 vssd1 vccd1 vccd1 _05999_ sky130_fd_sc_hd__nor2_1
XFILLER_91_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08331__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10904_ _05647_ _05648_ vssd1 vssd1 vccd1 vccd1 _05649_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_123_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14672_ clknet_leaf_23_clk _01377_ net1155 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_123_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11884_ net2587 net163 vssd1 vssd1 vccd1 vccd1 _05953_ sky130_fd_sc_hd__nand2_1
X_13623_ clknet_leaf_129_clk _00433_ net1114 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10835_ _04207_ _05589_ net899 vssd1 vssd1 vccd1 vccd1 _05590_ sky130_fd_sc_hd__mux2_1
XANTENNA__06893__A2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13090__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_24_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_8
X_13554_ clknet_leaf_33_clk _00364_ net1125 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09292__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10766_ datapath.PC\[5\] _05524_ vssd1 vssd1 vccd1 vccd1 _05531_ sky130_fd_sc_hd__nor2_1
X_12505_ net188 net1825 net506 vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__mux2_1
XFILLER_12_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13485_ clknet_leaf_131_clk _00295_ net1113 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10697_ net1477 _03292_ net570 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i_n\[2\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_145_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12436_ net1392 net130 _06365_ vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__a21o_1
XANTENNA__10729__A1 _02612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12367_ net229 _04906_ _05002_ _05685_ net893 vssd1 vssd1 vccd1 vccd1 _06329_ sky130_fd_sc_hd__o221a_1
XANTENNA__06940__B net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14106_ clknet_leaf_95_clk _00872_ net1226 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07070__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11318_ net2498 net275 net416 vssd1 vssd1 vccd1 vccd1 _00363_ sky130_fd_sc_hd__mux2_1
X_12298_ net890 _04580_ vssd1 vssd1 vccd1 vccd1 _06279_ sky130_fd_sc_hd__nor2_1
XANTENNA__07755__C net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14037_ clknet_leaf_85_clk _00806_ net1259 vssd1 vssd1 vccd1 vccd1 datapath.PC\[27\]
+ sky130_fd_sc_hd__dfrtp_4
X_11249_ net280 net2544 net420 vssd1 vssd1 vccd1 vccd1 _00298_ sky130_fd_sc_hd__mux2_1
XANTENNA__07358__B1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08570__A2 _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06790_ _01576_ _01584_ _01624_ vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__or3_2
XANTENNA__12103__B1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12389__B net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08858__A0 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10114__C1 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08322__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08460_ _03293_ _03294_ vssd1 vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__and2_2
XFILLER_91_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08883__A net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07530__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07411_ datapath.rf.registers\[7\]\[22\] net940 net931 vssd1 vssd1 vccd1 vccd1 _02247_
+ sky130_fd_sc_hd__and3_1
X_08391_ _03226_ vssd1 vssd1 vccd1 vccd1 _03227_ sky130_fd_sc_hd__inv_2
XANTENNA__09807__C1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_15_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_149_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07342_ datapath.rf.registers\[16\]\[24\] net739 _02177_ net787 vssd1 vssd1 vccd1
+ vccd1 _02178_ sky130_fd_sc_hd__a211o_1
XFILLER_31_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07273_ datapath.rf.registers\[14\]\[25\] net986 net919 vssd1 vssd1 vccd1 vccd1 _02109_
+ sky130_fd_sc_hd__and3_1
X_09012_ net346 _03847_ vssd1 vssd1 vccd1 vccd1 _03848_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_154_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold100 mmio.memload_or_instruction\[2\] vssd1 vssd1 vccd1 vccd1 net1448 sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 net59 vssd1 vssd1 vccd1 vccd1 net1459 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12344__S net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07946__B net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold122 net89 vssd1 vssd1 vccd1 vccd1 net1470 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold133 net77 vssd1 vssd1 vccd1 vccd1 net1481 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07597__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold144 net100 vssd1 vssd1 vccd1 vccd1 net1492 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold155 net86 vssd1 vssd1 vccd1 vccd1 net1503 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07061__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold166 datapath.multiplication_module.multiplicand_i\[24\] vssd1 vssd1 vccd1 vccd1
+ net1514 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07665__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_57_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold177 datapath.rf.registers\[7\]\[0\] vssd1 vssd1 vccd1 vccd1 net1525 sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 datapath.rf.registers\[15\]\[13\] vssd1 vssd1 vccd1 vccd1 net1536 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09914_ net604 _04747_ datapath.PC\[13\] vssd1 vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__o21a_1
Xfanout602 _06169_ vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__buf_2
Xhold199 datapath.rf.registers\[12\]\[0\] vssd1 vssd1 vccd1 vccd1 net1547 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout613 net614 vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1110_A net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout624 net625 vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__clkbuf_4
Xfanout635 net636 vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12342__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1208_A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout646 _01621_ vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input6_A DAT_I[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout657 _05364_ vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__buf_2
XFILLER_86_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09845_ _04670_ _04671_ _04672_ _04679_ vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__or4_1
XANTENNA__11696__A2 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout668 _01832_ vssd1 vssd1 vccd1 vccd1 net668 sky130_fd_sc_hd__buf_4
XANTENNA__09880__C net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout679 _01828_ vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__buf_4
XANTENNA_fanout668_A _01832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09776_ net332 _04545_ net311 vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__a21o_1
XFILLER_100_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06988_ net969 _01823_ vssd1 vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__and2_2
XFILLER_27_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08849__A0 _01935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08727_ _03031_ _03033_ vssd1 vssd1 vccd1 vccd1 _03563_ sky130_fd_sc_hd__or2_2
XFILLER_66_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08313__A2 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06865__X _01701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08658_ _02126_ _02146_ vssd1 vssd1 vccd1 vccd1 _03494_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_105_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07609_ datapath.rf.registers\[13\]\[18\] net981 net917 vssd1 vssd1 vccd1 vccd1 _02445_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10387__X _05223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout623_X net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08589_ _03173_ _03424_ _03174_ vssd1 vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__o21ba_1
XANTENNA__11423__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10620_ net38 _05381_ _05434_ vssd1 vssd1 vccd1 vccd1 _05440_ sky130_fd_sc_hd__and3_1
X_10551_ keypad.debounce.debounce\[9\] keypad.debounce.debounce\[8\] keypad.debounce.debounce\[11\]
+ keypad.debounce.debounce\[10\] vssd1 vssd1 vccd1 vccd1 _05378_ sky130_fd_sc_hd__and4_1
XFILLER_139_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13270_ clknet_leaf_142_clk _00080_ net1094 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10482_ screen.controlBus\[17\] screen.controlBus\[16\] screen.controlBus\[19\] screen.controlBus\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05312_ sky130_fd_sc_hd__or4_1
XFILLER_136_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout992_X net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12221_ _06223_ _06224_ vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__nor2_1
XFILLER_5_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07588__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12152_ _05800_ _06154_ vssd1 vssd1 vccd1 vccd1 _06182_ sky130_fd_sc_hd__and2b_1
XFILLER_150_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11103_ net172 net2141 net535 vssd1 vssd1 vccd1 vccd1 _00160_ sky130_fd_sc_hd__mux2_1
XANTENNA__10850__X _05603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12083_ screen.register.currentXbus\[6\] net1000 _05769_ screen.register.currentXbus\[22\]
+ vssd1 vssd1 vccd1 vccd1 _06122_ sky130_fd_sc_hd__a22o_1
XFILLER_150_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08968__A net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08537__C1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11034_ net172 net2406 net538 vssd1 vssd1 vccd1 vccd1 _00096_ sky130_fd_sc_hd__mux2_1
XANTENNA__13085__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08552__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07760__B1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12985_ net203 net2165 net478 vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__mux2_1
XFILLER_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08304__A2 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09501__A1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09501__B2 _03604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11936_ _02090_ net658 vssd1 vssd1 vccd1 vccd1 _05988_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_28_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14655_ clknet_leaf_11_clk _01360_ net1082 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_11867_ _03226_ screen.counter.ack vssd1 vssd1 vccd1 vccd1 _05942_ sky130_fd_sc_hd__or2_1
XFILLER_14_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06935__B _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11333__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13606_ clknet_leaf_17_clk _00416_ net1106 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_151_Left_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10818_ net262 net2131 net544 vssd1 vssd1 vccd1 vccd1 _00014_ sky130_fd_sc_hd__mux2_1
X_14586_ clknet_leaf_146_clk _01291_ net1065 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09265__B1 _02418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11798_ datapath.ru.latched_instruction\[4\] net333 net313 _01569_ vssd1 vssd1 vccd1
+ vccd1 _00664_ sky130_fd_sc_hd__a22o_1
XANTENNA__08208__A net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13537_ clknet_leaf_56_clk _00347_ net1171 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10749_ _01606_ _01783_ vssd1 vssd1 vccd1 vccd1 _05516_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_136_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13468_ clknet_leaf_10_clk _00278_ net1080 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07291__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06951__A net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09568__A1 _02805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12419_ _05976_ net156 vssd1 vssd1 vccd1 vccd1 _06357_ sky130_fd_sc_hd__nor2_1
XFILLER_127_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13399_ clknet_leaf_127_clk _00209_ net1208 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07043__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11856__X _05934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09981__B net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07960_ datapath.rf.registers\[14\]\[11\] net830 net828 datapath.rf.registers\[12\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__a22o_1
XANTENNA__12324__A0 _04118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_4_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_8
X_06911_ datapath.rf.registers\[26\]\[31\] net836 net832 datapath.rf.registers\[30\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__a22o_1
XANTENNA__10335__C1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07891_ _02704_ _02726_ vssd1 vssd1 vccd1 vccd1 _02727_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_155_Right_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11508__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10886__B1 _05632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09630_ net380 _04464_ _04465_ _03613_ vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__o211a_1
XANTENNA__08543__A2 _01740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06842_ net1003 net1019 _01677_ net1027 datapath.ru.latched_instruction\[15\] vssd1
+ vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__a32o_2
XTAP_TAPCELL_ROW_52_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07751__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06773_ datapath.ru.latched_instruction\[14\] net1030 _01568_ _01513_ vssd1 vssd1
+ vccd1 vccd1 _01610_ sky130_fd_sc_hd__o2bb2a_2
X_09561_ _03424_ _03556_ vssd1 vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__xnor2_2
X_08512_ datapath.rf.registers\[21\]\[1\] net963 _01831_ vssd1 vssd1 vccd1 vccd1 _03348_
+ sky130_fd_sc_hd__and3_1
XFILLER_130_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09492_ net331 _04095_ _04096_ _04316_ _04327_ vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__o32a_2
XFILLER_63_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06857__A2 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08443_ datapath.rf.registers\[8\]\[2\] net697 net666 datapath.rf.registers\[15\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__a22o_1
XANTENNA__12339__S net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout151_A _05886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout249_A net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11243__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08374_ datapath.rf.registers\[16\]\[3\] net740 net690 datapath.rf.registers\[31\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03210_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_156_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07325_ datapath.rf.registers\[10\]\[24\] net880 net855 datapath.rf.registers\[19\]\[24\]
+ _02160_ vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__a221o_1
XFILLER_139_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10935__X _05676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout416_A net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1158_A net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07256_ _02069_ _02091_ vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__nand2_1
XANTENNA__09008__B1 _02025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07282__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07187_ datapath.rf.registers\[12\]\[27\] net827 _02020_ _02021_ _02022_ vssd1 vssd1
+ vccd1 vccd1 _02023_ sky130_fd_sc_hd__a2111o_1
XFILLER_3_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07034__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14005__D screen.counter.ack vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12802__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13798__RESET_B net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout410 _05730_ vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08788__A _01637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout421 _05722_ vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout432 net433 vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_6_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout443 _03760_ vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__clkbuf_4
Xfanout454 net456 vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__buf_2
XANTENNA_fanout573_X net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout952_A net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11418__S net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08534__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout476 net477 vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__clkbuf_8
Xfanout487 _06552_ vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__clkbuf_4
X_09828_ _04649_ _04663_ _04647_ vssd1 vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__a21o_2
XPHY_EDGE_ROW_122_Right_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout498 net499 vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__buf_2
XFILLER_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07742__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09759_ net337 _04593_ _04594_ net322 vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout740_X net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout838_X net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11942__A _02001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ net290 net2475 net494 vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__mux2_1
XANTENNA__09495__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ net7 net1036 _05889_ net2360 vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__a22o_1
XANTENNA__11661__B _05874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06848__A2 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10558__A _05315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11153__S net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14440_ clknet_leaf_90_clk _01145_ net1233 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11652_ _04711_ _05874_ vssd1 vssd1 vccd1 vccd1 _05875_ sky130_fd_sc_hd__nor2_2
XANTENNA__12458__A1_N net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10603_ screen.register.currentYbus\[21\] screen.register.currentYbus\[20\] screen.register.currentYbus\[23\]
+ screen.register.currentYbus\[22\] vssd1 vssd1 vccd1 vccd1 _05424_ sky130_fd_sc_hd__or4_1
XANTENNA__09798__A1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14371_ clknet_leaf_120_clk _01076_ net1192 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10992__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10845__X _05599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11583_ _01422_ screen.counter.ct\[5\] net1278 net1279 vssd1 vssd1 vccd1 vccd1 _05807_
+ sky130_fd_sc_hd__or4_1
XFILLER_156_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13322_ clknet_leaf_21_clk _00132_ net1164 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10534_ _05333_ _05348_ _05363_ _05321_ _05304_ vssd1 vssd1 vccd1 vccd1 _05364_ sky130_fd_sc_hd__a32oi_2
XFILLER_6_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06771__A _01575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13253_ clknet_leaf_139_clk _00063_ net1099 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10465_ screen.counter.ct\[21\] screen.counter.ct\[20\] screen.counter.ct\[22\] vssd1
+ vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__or3_1
XFILLER_6_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12204_ screen.counter.currentCt\[4\] _06210_ screen.counter.currentCt\[5\] vssd1
+ vssd1 vccd1 vccd1 _06213_ sky130_fd_sc_hd__a21oi_1
X_13184_ net2021 vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__clkbuf_1
X_10396_ net346 _04164_ _05231_ _03644_ vssd1 vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__a22o_1
XFILLER_135_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12135_ _06168_ net601 vssd1 vssd1 vccd1 vccd1 _06172_ sky130_fd_sc_hd__or2_2
XFILLER_96_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08698__A _02857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12066_ _05330_ _05795_ _05842_ _06074_ vssd1 vssd1 vccd1 vccd1 _06106_ sky130_fd_sc_hd__a31o_1
XANTENNA__11328__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11017_ net256 net1918 net539 vssd1 vssd1 vccd1 vccd1 _00079_ sky130_fd_sc_hd__mux2_1
XANTENNA__07733__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12968_ net291 net1859 net478 vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__mux2_1
XANTENNA__09486__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08828__A3 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_0_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11919_ net134 _05976_ _05975_ vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11063__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12899_ net1685 net302 net484 vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__mux2_1
XFILLER_21_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14638_ clknet_leaf_0_clk _01343_ net1055 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_138_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09238__B1 _03770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14569_ clknet_leaf_20_clk _01274_ net1165 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_147_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08880__B _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07110_ datapath.rf.registers\[12\]\[29\] net755 net730 datapath.rf.registers\[19\]\[29\]
+ _01945_ vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__a221o_1
XANTENNA__10399__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07777__A _02612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08090_ datapath.rf.registers\[14\]\[9\] net776 net712 datapath.rf.registers\[11\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_151_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload20 clknet_leaf_148_clk vssd1 vssd1 vccd1 vccd1 clkload20/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_151_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07041_ datapath.rf.registers\[5\]\[30\] net820 net816 datapath.rf.registers\[21\]\[30\]
+ _01876_ vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__a221o_1
Xclkload31 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 clkload31/X sky130_fd_sc_hd__clkbuf_8
Xclkload42 clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 clkload42/Y sky130_fd_sc_hd__inv_6
Xclkload53 clknet_leaf_134_clk vssd1 vssd1 vccd1 vccd1 clkload53/Y sky130_fd_sc_hd__inv_8
Xclkload64 clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 clkload64/Y sky130_fd_sc_hd__bufinv_16
Xclkload75 clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 clkload75/Y sky130_fd_sc_hd__bufinv_16
Xclkload86 clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 clkload86/Y sky130_fd_sc_hd__inv_6
XANTENNA__09410__B1 _02704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload97 clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 clkload97/Y sky130_fd_sc_hd__inv_8
XFILLER_142_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08992_ _02048_ _02049_ vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__and2b_1
XFILLER_142_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09056__X _03892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07972__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07943_ datapath.rf.registers\[27\]\[11\] net976 net938 vssd1 vssd1 vccd1 vccd1 _02779_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07943__C net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11238__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09713__B2 _03614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07874_ datapath.rf.registers\[11\]\[13\] net710 net683 datapath.rf.registers\[27\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__a22o_1
XFILLER_29_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07724__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09613_ net323 _04053_ vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__nor2_1
X_06825_ _01659_ _01660_ datapath.ru.latched_instruction\[9\] vssd1 vssd1 vccd1 vccd1
+ _01661_ sky130_fd_sc_hd__mux2_1
XFILLER_141_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout366_A net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09544_ net363 _04375_ vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__or2_1
X_06756_ _01477_ net1016 net994 net1029 datapath.ru.latched_instruction\[31\] vssd1
+ vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__a32oi_4
XANTENNA__09477__B1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11823__A2 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06687_ _01520_ _01521_ _01522_ _01525_ vssd1 vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__or4_1
X_09475_ net457 _04303_ _04310_ net350 vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__a211o_1
XANTENNA__10378__A _01859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08426_ datapath.rf.registers\[0\]\[2\] net868 _03261_ vssd1 vssd1 vccd1 vccd1 _03262_
+ sky130_fd_sc_hd__o21a_2
XTAP_TAPCELL_ROW_22_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10097__B net1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout700_A net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08357_ datapath.rf.registers\[17\]\[3\] net851 net797 datapath.rf.registers\[29\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03193_ sky130_fd_sc_hd__a22o_1
XFILLER_20_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout419_X net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload3 clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clkload3/X sky130_fd_sc_hd__clkbuf_8
XFILLER_50_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07308_ _02127_ _02133_ _02135_ _02143_ vssd1 vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__or4_4
XANTENNA__07255__A2 _02090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08288_ _01604_ _01784_ vssd1 vssd1 vccd1 vccd1 _03124_ sky130_fd_sc_hd__nor2_1
XFILLER_137_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07239_ datapath.rf.registers\[18\]\[26\] net722 net698 datapath.rf.registers\[23\]\[26\]
+ _02072_ vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__a221o_1
XFILLER_106_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10250_ _04300_ _04563_ net890 vssd1 vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07007__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout690_X net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout788_X net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10181_ _04882_ _05016_ vssd1 vssd1 vccd1 vccd1 _05017_ sky130_fd_sc_hd__nand2b_1
Xfanout1205 net1213 vssd1 vssd1 vccd1 vccd1 net1205 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06766__B2 datapath.ru.latched_instruction\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1216 net1217 vssd1 vssd1 vccd1 vccd1 net1216 sky130_fd_sc_hd__clkbuf_4
Xfanout1227 net1231 vssd1 vssd1 vccd1 vccd1 net1227 sky130_fd_sc_hd__clkbuf_4
Xfanout240 net242 vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__clkbuf_2
Xfanout1238 net1251 vssd1 vssd1 vccd1 vccd1 net1238 sky130_fd_sc_hd__buf_2
XANTENNA_fanout955_X net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1249 net1250 vssd1 vssd1 vccd1 vccd1 net1249 sky130_fd_sc_hd__clkbuf_4
Xfanout251 net252 vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11148__S net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout262 _05575_ vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_89_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13940_ clknet_leaf_95_clk _00718_ net1216 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_89_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout273 _05564_ vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__buf_1
XFILLER_87_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout284 net285 vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07715__B1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout295 net297 vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13871_ clknet_leaf_53_clk _00675_ net1183 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10987__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12822_ net1937 net196 net492 vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__mux2_1
XANTENNA__09468__B1 _03205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11275__A0 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12753_ net1975 net210 net402 vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__mux2_1
XFILLER_42_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11704_ mmio.wishbone.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1 _05888_ sky130_fd_sc_hd__nand2_1
X_12684_ _06514_ _06515_ _06512_ vssd1 vssd1 vccd1 vccd1 _06517_ sky130_fd_sc_hd__o21a_1
XFILLER_30_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14423_ clknet_leaf_124_clk _01128_ net1208 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11635_ _05809_ _05815_ _05816_ _05817_ vssd1 vssd1 vccd1 vccd1 _05859_ sky130_fd_sc_hd__or4b_1
XFILLER_128_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09288__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07246__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14354_ clknet_leaf_30_clk _01059_ net1135 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11566_ net1009 _05775_ vssd1 vssd1 vccd1 vccd1 _05790_ sky130_fd_sc_hd__nor2_1
XFILLER_156_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13305_ clknet_leaf_30_clk _00115_ net1131 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10517_ net1279 net1274 net1270 screen.counter.ct\[20\] _05344_ vssd1 vssd1 vccd1
+ vccd1 _05347_ sky130_fd_sc_hd__a41o_1
XFILLER_6_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14285_ clknet_leaf_123_clk _00990_ net1199 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11497_ net235 net1716 net512 vssd1 vssd1 vccd1 vccd1 _00533_ sky130_fd_sc_hd__mux2_1
XFILLER_143_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13236_ clknet_leaf_128_clk _00046_ net1117 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10448_ _05282_ _05283_ vssd1 vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__and2_1
XANTENNA__12712__A_N _05894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13167_ net1968 vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__clkbuf_1
X_10379_ _03720_ _04682_ _04685_ _05214_ _05213_ vssd1 vssd1 vccd1 vccd1 _05215_ sky130_fd_sc_hd__a41o_1
XANTENNA__06757__B2 datapath.ru.latched_instruction\[29\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_97_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07954__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11750__B2 _02876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12118_ net1277 _05907_ _06154_ vssd1 vssd1 vccd1 vccd1 _06155_ sky130_fd_sc_hd__and3_1
XFILLER_112_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13098_ net303 net2212 net472 vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__mux2_1
XFILLER_78_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11058__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12049_ screen.register.currentXbus\[12\] _05768_ _06019_ screen.register.currentYbus\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06090_ sky130_fd_sc_hd__a22o_1
XFILLER_66_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10305__A2 _04580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07706__B1 _02536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06610_ mmio.key_data\[4\] net1049 _01448_ vssd1 vssd1 vccd1 vccd1 _01449_ sky130_fd_sc_hd__o21ai_1
X_07590_ datapath.rf.registers\[17\]\[19\] net748 net724 datapath.rf.registers\[18\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__a22o_1
XANTENNA__09459__B1 _03718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12397__B net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11805__A2 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08131__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09260_ net374 _03836_ _03833_ net376 vssd1 vssd1 vccd1 vccd1 _04096_ sky130_fd_sc_hd__a211oi_1
XFILLER_21_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07485__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08211_ datapath.rf.registers\[11\]\[6\] net882 net860 datapath.rf.registers\[16\]\[6\]
+ _03046_ vssd1 vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__a221o_1
X_09191_ _03584_ _04024_ net578 vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__o21a_1
X_08142_ datapath.rf.registers\[24\]\[8\] net768 net667 datapath.rf.registers\[15\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__a22o_1
XFILLER_146_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07237__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07938__C net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload120 clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 clkload120/Y sky130_fd_sc_hd__clkinv_4
X_08073_ datapath.rf.registers\[16\]\[9\] net862 net854 datapath.rf.registers\[19\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__a22o_1
Xclkload131 clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 clkload131/Y sky130_fd_sc_hd__inv_6
Xclkload142 clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 clkload142/Y sky130_fd_sc_hd__clkinvlp_4
X_07024_ _01859_ vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__inv_2
XFILLER_143_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08198__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06748__A1 _01443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11741__B2 _03357_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08975_ net448 _03810_ vssd1 vssd1 vccd1 vccd1 _03811_ sky130_fd_sc_hd__nand2_1
Xhold15 screen.screenEdge.enable2 vssd1 vssd1 vccd1 vccd1 net1363 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout483_A _06554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold26 datapath.pc_module.i_ack1 vssd1 vssd1 vccd1 vccd1 net1374 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold37 datapath.i_ack vssd1 vssd1 vccd1 vccd1 net1385 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07018__Y _01854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07926_ datapath.rf.registers\[23\]\[12\] net701 net674 datapath.rf.registers\[7\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__a22o_1
XFILLER_130_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold48 net68 vssd1 vssd1 vccd1 vccd1 net1396 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 net70 vssd1 vssd1 vccd1 vccd1 net1407 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_68_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07857_ datapath.rf.registers\[8\]\[13\] net877 net798 datapath.rf.registers\[29\]\[13\]
+ _02692_ vssd1 vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout650_A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout369_X net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout748_A net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06808_ datapath.ru.latched_instruction\[7\] net1028 net993 _01642_ vssd1 vssd1 vccd1
+ vccd1 _01644_ sky130_fd_sc_hd__a22o_1
XFILLER_84_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07788_ datapath.rf.registers\[30\]\[15\] net759 net672 datapath.rf.registers\[7\]\[15\]
+ _02621_ vssd1 vssd1 vccd1 vccd1 _02624_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_84_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09527_ net357 _04359_ vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__nand2_1
XANTENNA__14178__RESET_B net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06739_ _01486_ net1014 vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout1180_X net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout915_A net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout536_X net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09458_ net574 _04285_ _04286_ _04293_ vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__a22o_1
XFILLER_52_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08409_ datapath.rf.registers\[26\]\[2\] net979 _01720_ vssd1 vssd1 vccd1 vccd1 _03245_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout703_X net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09389_ net328 _03983_ _03623_ vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__o21a_1
XANTENNA__11431__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11420_ net272 net2303 net516 vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__mux2_1
XANTENNA__07228__A2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07848__C net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07210__A _02045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11351_ net280 net2299 net521 vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_115_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10302_ _01702_ _04580_ _05137_ net1040 vssd1 vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__o211a_1
X_14070_ clknet_leaf_111_clk _00837_ net1196 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11282_ net279 net1922 net525 vssd1 vssd1 vccd1 vccd1 _00330_ sky130_fd_sc_hd__mux2_1
XFILLER_4_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08189__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13021_ net2270 net194 net391 vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__mux2_1
XFILLER_140_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10233_ _04829_ _04892_ vssd1 vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__and2b_1
XANTENNA__10571__A _02804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07936__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07209__X _02045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10164_ _04177_ _04584_ _04999_ vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__o21ai_1
Xfanout1002 net1004 vssd1 vssd1 vccd1 vccd1 net1002 sky130_fd_sc_hd__buf_4
Xfanout1013 _05433_ vssd1 vssd1 vccd1 vccd1 net1013 sky130_fd_sc_hd__buf_2
Xfanout1024 _05890_ vssd1 vssd1 vccd1 vccd1 net1024 sky130_fd_sc_hd__clkbuf_2
XFILLER_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1035 _05887_ vssd1 vssd1 vccd1 vccd1 net1035 sky130_fd_sc_hd__buf_2
X_10095_ net225 _04885_ _04930_ vssd1 vssd1 vccd1 vccd1 _04931_ sky130_fd_sc_hd__nand3_1
Xfanout1057 net1058 vssd1 vssd1 vccd1 vccd1 net1057 sky130_fd_sc_hd__clkbuf_2
Xfanout1068 net1075 vssd1 vssd1 vccd1 vccd1 net1068 sky130_fd_sc_hd__clkbuf_4
Xfanout1079 net1084 vssd1 vssd1 vccd1 vccd1 net1079 sky130_fd_sc_hd__clkbuf_2
X_13923_ clknet_leaf_109_clk _00701_ net1218 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06767__Y _01604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13093__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13854_ clknet_leaf_49_clk _00658_ net1176 vssd1 vssd1 vccd1 vccd1 keypad.apps.app_c\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12805_ net1721 net281 net493 vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__mux2_1
X_13785_ clknet_leaf_52_clk _00594_ net1183 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08982__Y _03818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10997_ net1669 net178 net437 vssd1 vssd1 vccd1 vccd1 _00062_ sky130_fd_sc_hd__mux2_1
XANTENNA__11799__B2 _01441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12736_ net1944 net295 net402 vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__mux2_1
XANTENNA__07467__A2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12667_ datapath.mulitply_result\[26\] datapath.multiplication_module.multiplicand_i\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06503_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_13_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14406_ clknet_leaf_17_clk _01111_ net1107 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_128_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11618_ _05839_ _05841_ _05766_ vssd1 vssd1 vccd1 vccd1 _05842_ sky130_fd_sc_hd__and3b_1
XANTENNA__07219__A2 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07758__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12598_ net2513 net505 net501 _06445_ vssd1 vssd1 vccd1 vccd1 _00924_ sky130_fd_sc_hd__a22o_1
X_14337_ clknet_leaf_37_clk _01042_ net1137 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11549_ _05751_ net1006 vssd1 vssd1 vccd1 vccd1 _05773_ sky130_fd_sc_hd__nor2_4
XFILLER_116_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold507 datapath.rf.registers\[9\]\[6\] vssd1 vssd1 vccd1 vccd1 net1855 sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 datapath.rf.registers\[18\]\[26\] vssd1 vssd1 vccd1 vccd1 net1866 sky130_fd_sc_hd__dlygate4sd3_1
Xhold529 datapath.rf.registers\[3\]\[19\] vssd1 vssd1 vccd1 vccd1 net1877 sky130_fd_sc_hd__dlygate4sd3_1
X_14268_ clknet_leaf_9_clk _00973_ net1074 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_143_246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13219_ clknet_leaf_120_clk _00029_ net1192 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_14199_ clknet_leaf_66_clk datapath.multiplication_module.multiplicand_i_n\[10\]
+ net1237 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07927__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1207 datapath.rf.registers\[10\]\[17\] vssd1 vssd1 vccd1 vccd1 net2555 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12900__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08760_ _03487_ _03489_ _03594_ _03485_ vssd1 vssd1 vccd1 vccd1 _03596_ sky130_fd_sc_hd__a31oi_1
XTAP_TAPCELL_ROW_146_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_29_Left_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1218 datapath.rf.registers\[31\]\[26\] vssd1 vssd1 vccd1 vccd1 net2566 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06958__X _01794_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1229 datapath.rf.registers\[29\]\[28\] vssd1 vssd1 vccd1 vccd1 net2577 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08886__A _01611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07711_ datapath.rf.registers\[26\]\[16\] net974 net937 vssd1 vssd1 vccd1 vccd1 _02547_
+ sky130_fd_sc_hd__and3_1
X_08691_ _02751_ _02772_ vssd1 vssd1 vccd1 vccd1 _03527_ sky130_fd_sc_hd__nor2_1
X_07642_ datapath.rf.registers\[2\]\[18\] net742 net718 datapath.rf.registers\[20\]\[18\]
+ _02477_ vssd1 vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__a221o_1
XFILLER_19_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07573_ datapath.rf.registers\[1\]\[19\] net847 _02392_ _02400_ _02404_ vssd1 vssd1
+ vccd1 vccd1 _02409_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08104__B1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09312_ net630 _04147_ vssd1 vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__nor2_1
XFILLER_34_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09510__A _03205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09243_ _03505_ net627 _04078_ net644 vssd1 vssd1 vccd1 vccd1 _04079_ sky130_fd_sc_hd__a211oi_1
XANTENNA__07949__B net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_38_Left_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11251__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09174_ _03801_ _03803_ net448 vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__mux2_1
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07668__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08125_ _02960_ vssd1 vssd1 vccd1 vccd1 _02961_ sky130_fd_sc_hd__clkinv_4
XFILLER_147_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1238_A net1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07091__B1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08056_ datapath.rf.registers\[26\]\[9\] net977 net937 vssd1 vssd1 vccd1 vccd1 _02892_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout698_A net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07007_ datapath.rf.registers\[14\]\[31\] net774 net676 datapath.rf.registers\[29\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__a22o_1
XANTENNA__07602__A2_N net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput49 net49 vssd1 vssd1 vccd1 vccd1 ADR_O[18] sky130_fd_sc_hd__buf_2
XFILLER_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07918__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08499__C _01816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout486_X net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout865_A _01726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12810__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08958_ net561 _02613_ net445 vssd1 vssd1 vccd1 vccd1 _03794_ sky130_fd_sc_hd__mux2_1
X_07909_ datapath.rf.registers\[22\]\[12\] net822 net820 datapath.rf.registers\[5\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__a22o_1
X_08889_ net904 _01859_ _03698_ _03723_ _03724_ vssd1 vssd1 vccd1 vccd1 _03725_ sky130_fd_sc_hd__o2111a_1
XFILLER_56_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11426__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10920_ datapath.mulitply_result\[27\] net597 net618 vssd1 vssd1 vccd1 vccd1 _05663_
+ sky130_fd_sc_hd__a21o_1
XFILLER_45_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07697__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10851_ datapath.mulitply_result\[17\] net597 _05603_ vssd1 vssd1 vccd1 vccd1 _05604_
+ sky130_fd_sc_hd__a21bo_1
XANTENNA_fanout820_X net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout918_X net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13570_ clknet_leaf_150_clk _00380_ net1053 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10782_ _04495_ _05544_ net901 vssd1 vssd1 vccd1 vccd1 _05545_ sky130_fd_sc_hd__mux2_1
X_12521_ datapath.mulitply_result\[2\] datapath.multiplication_module.multiplicand_i\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06381_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_40_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11161__S net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12452_ net167 _05952_ net129 net2654 vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__a2bb2o_1
X_11403_ net2071 net192 net410 vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12383_ _05940_ net159 vssd1 vssd1 vccd1 vccd1 _06339_ sky130_fd_sc_hd__nor2_1
XFILLER_126_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10756__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14122_ clknet_leaf_21_clk _00879_ net1163 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07082__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11334_ net2213 net197 net416 vssd1 vssd1 vccd1 vccd1 _00379_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_55_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13088__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09359__C1 _02612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14053_ clknet_leaf_101_clk _00820_ net1228 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11265_ net200 net1560 net419 vssd1 vssd1 vccd1 vccd1 _00314_ sky130_fd_sc_hd__mux2_1
XFILLER_137_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07909__B1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13004_ net1977 net274 net392 vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__mux2_1
X_10216_ _04966_ _05009_ _05051_ vssd1 vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__or3_2
XFILLER_140_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11196_ net210 net2193 net422 vssd1 vssd1 vccd1 vccd1 _00248_ sky130_fd_sc_hd__mux2_1
XANTENNA__08202__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08582__B1 _03384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10147_ _04625_ _04982_ _04981_ net226 vssd1 vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__a211o_1
XFILLER_67_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_113_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10078_ _03752_ _04913_ net1044 vssd1 vssd1 vccd1 vccd1 _04914_ sky130_fd_sc_hd__o21a_1
XANTENNA__08334__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11336__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13906_ clknet_leaf_42_clk net1369 net1149 vssd1 vssd1 vccd1 vccd1 keypad.debounce.debounce\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14029__RESET_B net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07688__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13837_ clknet_leaf_115_clk _00646_ net1187 vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_128_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13768_ clknet_leaf_82_clk _00577_ net1256 vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__dfrtp_1
X_12719_ columns.count\[6\] _06538_ columns.count\[7\] vssd1 vssd1 vccd1 vccd1 _06542_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_44_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_13699_ clknet_leaf_120_clk _00509_ net1200 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_44_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14131__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07860__A2 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10763__X _05529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold304 datapath.rf.registers\[11\]\[30\] vssd1 vssd1 vccd1 vccd1 net1652 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07073__B1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold315 datapath.rf.registers\[22\]\[1\] vssd1 vssd1 vccd1 vccd1 net1663 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold326 datapath.rf.registers\[6\]\[8\] vssd1 vssd1 vccd1 vccd1 net1674 sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 datapath.rf.registers\[16\]\[3\] vssd1 vssd1 vccd1 vccd1 net1685 sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 datapath.rf.registers\[4\]\[20\] vssd1 vssd1 vccd1 vccd1 net1696 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09930_ datapath.PC\[7\] _03029_ vssd1 vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__and2_1
Xhold359 datapath.rf.registers\[13\]\[29\] vssd1 vssd1 vccd1 vccd1 net1707 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout806 _01768_ vssd1 vssd1 vccd1 vccd1 net806 sky130_fd_sc_hd__clkbuf_8
Xfanout817 net818 vssd1 vssd1 vccd1 vccd1 net817 sky130_fd_sc_hd__buf_4
X_09861_ _02827_ _02881_ _03435_ _04674_ vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__o22a_1
Xfanout828 _01749_ vssd1 vssd1 vccd1 vccd1 net828 sky130_fd_sc_hd__clkbuf_8
XFILLER_98_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout839 net840 vssd1 vssd1 vccd1 vccd1 net839 sky130_fd_sc_hd__clkbuf_8
X_08812_ _01636_ _03644_ vssd1 vssd1 vccd1 vccd1 _03648_ sky130_fd_sc_hd__nand2_1
XFILLER_86_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_783 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1004 datapath.rf.registers\[26\]\[12\] vssd1 vssd1 vccd1 vccd1 net2352 sky130_fd_sc_hd__dlygate4sd3_1
X_09792_ _04627_ vssd1 vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__inv_2
Xhold1015 datapath.rf.registers\[8\]\[14\] vssd1 vssd1 vccd1 vccd1 net2363 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10380__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1026 datapath.rf.registers\[22\]\[15\] vssd1 vssd1 vccd1 vccd1 net2374 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09505__A _03009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08743_ _03518_ _03521_ _03576_ _03517_ _03515_ vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__a311o_1
Xhold1037 datapath.rf.registers\[1\]\[0\] vssd1 vssd1 vccd1 vccd1 net2385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1048 datapath.rf.registers\[3\]\[26\] vssd1 vssd1 vccd1 vccd1 net2396 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07951__C net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1059 datapath.rf.registers\[24\]\[27\] vssd1 vssd1 vccd1 vccd1 net2407 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11246__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout279_A _05554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07679__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08674_ _02466_ _02488_ vssd1 vssd1 vccd1 vccd1 _03510_ sky130_fd_sc_hd__nand2_1
XANTENNA__08876__A1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07625_ datapath.rf.registers\[4\]\[18\] net864 net790 datapath.rf.registers\[18\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout446_A net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1188_A net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_46_Left_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07556_ datapath.rf.registers\[12\]\[19\] net955 net920 vssd1 vssd1 vccd1 vccd1 _02392_
+ sky130_fd_sc_hd__and3_1
X_07487_ datapath.rf.registers\[14\]\[21\] net774 net710 datapath.rf.registers\[11\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02323_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout613_A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09226_ net364 _03986_ vssd1 vssd1 vccd1 vccd1 _04062_ sky130_fd_sc_hd__nand2_1
XFILLER_21_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09157_ net461 _03773_ _03992_ vssd1 vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout401_X net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12805__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06870__Y _01706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07064__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08108_ datapath.rf.registers\[10\]\[8\] net881 net797 datapath.rf.registers\[29\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__a22o_1
X_09088_ net377 _03923_ _03623_ vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout982_A net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08039_ _02872_ _02873_ _02874_ vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_55_Left_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold860 datapath.rf.registers\[20\]\[23\] vssd1 vssd1 vccd1 vccd1 net2208 sky130_fd_sc_hd__dlygate4sd3_1
Xhold871 datapath.rf.registers\[0\]\[28\] vssd1 vssd1 vccd1 vccd1 net2219 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold882 mmio.memload_or_instruction\[30\] vssd1 vssd1 vccd1 vccd1 net2230 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold893 datapath.rf.registers\[0\]\[6\] vssd1 vssd1 vccd1 vccd1 net2241 sky130_fd_sc_hd__dlygate4sd3_1
X_11050_ net264 net2310 net431 vssd1 vssd1 vccd1 vccd1 _00110_ sky130_fd_sc_hd__mux2_1
XANTENNA__11699__B1 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout770_X net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10001_ _04784_ _04786_ vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11945__A _01954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09108__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07119__A1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11156__S net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11952_ net134 _05998_ _05997_ vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__o21ai_1
XFILLER_85_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10903_ net1264 _05636_ datapath.PC\[25\] vssd1 vssd1 vccd1 vccd1 _05648_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10995__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Left_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14671_ clknet_leaf_30_clk _01376_ net1132 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_123_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11883_ net137 _05952_ _05951_ vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_123_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13622_ clknet_leaf_142_clk _00432_ net1094 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10834_ datapath.PC\[15\] _05583_ vssd1 vssd1 vccd1 vccd1 _05589_ sky130_fd_sc_hd__xor2_1
XFILLER_16_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13553_ clknet_leaf_41_clk _00363_ net1140 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10765_ datapath.PC\[5\] _05524_ vssd1 vssd1 vccd1 vccd1 _05530_ sky130_fd_sc_hd__and2_1
XANTENNA__08095__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12504_ net192 net2566 net506 vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__mux2_1
XANTENNA__07842__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13484_ clknet_leaf_16_clk _00294_ net1106 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10696_ net1450 _03357_ net570 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i_n\[1\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12435_ _05992_ net156 vssd1 vssd1 vccd1 vccd1 _06365_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07055__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_73_Left_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12366_ _06326_ _06328_ datapath.PC\[30\] net309 vssd1 vssd1 vccd1 vccd1 _00809_
+ sky130_fd_sc_hd__a2bb2o_1
XPHY_EDGE_ROW_136_Right_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14105_ clknet_leaf_95_clk _00871_ net1226 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_141_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11317_ net1858 net278 net416 vssd1 vssd1 vccd1 vccd1 _00362_ sky130_fd_sc_hd__mux2_1
X_12297_ datapath.PC\[11\] _06278_ net307 vssd1 vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__mux2_1
X_14036_ clknet_leaf_85_clk _00805_ net1259 vssd1 vssd1 vccd1 vccd1 datapath.PC\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11248_ net285 net1757 net420 vssd1 vssd1 vccd1 vccd1 _00297_ sky130_fd_sc_hd__mux2_1
XFILLER_110_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11179_ net294 net1576 net422 vssd1 vssd1 vccd1 vccd1 _00231_ sky130_fd_sc_hd__mux2_1
XANTENNA__10362__B1 net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06949__A _01593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08307__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11066__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08858__A1 _01889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09979__B net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08883__B _03718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07410_ datapath.rf.registers\[21\]\[22\] net815 net813 datapath.rf.registers\[23\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__a22o_1
X_08390_ datapath.rf.registers\[0\]\[3\] net783 _03216_ _03225_ vssd1 vssd1 vccd1
+ vccd1 _03226_ sky130_fd_sc_hd__o22ai_4
X_07341_ datapath.rf.registers\[11\]\[24\] net711 net680 datapath.rf.registers\[6\]\[24\]
+ _02176_ vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__a221o_1
XANTENNA__08086__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07294__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07272_ datapath.rf.registers\[25\]\[25\] net978 net943 vssd1 vssd1 vccd1 vccd1 _02108_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07833__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09011_ net350 _03842_ _03845_ _03846_ net359 vssd1 vssd1 vccd1 vccd1 _03847_ sky130_fd_sc_hd__o311ai_2
XTAP_TAPCELL_ROW_154_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07046__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold101 mmio.key_data\[1\] vssd1 vssd1 vccd1 vccd1 net1449 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold112 net117 vssd1 vssd1 vccd1 vccd1 net1460 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07946__C net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold123 datapath.multiplication_module.multiplier_i\[5\] vssd1 vssd1 vccd1 vccd1
+ net1471 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold134 net90 vssd1 vssd1 vccd1 vccd1 net1482 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_103_Right_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold145 net101 vssd1 vssd1 vccd1 vccd1 net1493 sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 datapath.multiplication_module.multiplicand_i\[26\] vssd1 vssd1 vccd1 vccd1
+ net1504 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 net73 vssd1 vssd1 vccd1 vccd1 net1515 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_99_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09913_ _04748_ vssd1 vssd1 vccd1 vccd1 _04749_ sky130_fd_sc_hd__inv_2
Xhold178 net97 vssd1 vssd1 vccd1 vccd1 net1526 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout603 _06169_ vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_74_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold189 datapath.rf.registers\[13\]\[17\] vssd1 vssd1 vccd1 vccd1 net1537 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout614 _01781_ vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout396_A _06555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout625 _03721_ vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__clkbuf_4
Xfanout636 _01627_ vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09743__C1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09844_ _03420_ _03548_ _04339_ _04678_ vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__or4_1
Xfanout647 _01609_ vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__clkbuf_4
XFILLER_113_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout658 net659 vssd1 vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1103_A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout669 _01832_ vssd1 vssd1 vccd1 vccd1 net669 sky130_fd_sc_hd__buf_4
X_09775_ _03592_ _04610_ net579 vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__o21ai_1
XFILLER_39_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout563_A _02264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06987_ net991 _01637_ _01647_ net972 vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__and4_2
XFILLER_85_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08726_ _03559_ _03561_ _03541_ vssd1 vssd1 vccd1 vccd1 _03562_ sky130_fd_sc_hd__a21o_1
XANTENNA__08849__A1 _01981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08657_ _02126_ _02146_ vssd1 vssd1 vccd1 vccd1 _03493_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout730_A _01811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout828_A _01749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07608_ datapath.rf.registers\[25\]\[18\] net841 vssd1 vssd1 vccd1 vccd1 _02444_
+ sky130_fd_sc_hd__nand2_1
X_08588_ _03230_ _03423_ _03231_ vssd1 vssd1 vccd1 vccd1 _03424_ sky130_fd_sc_hd__a21oi_2
X_07539_ datapath.rf.registers\[3\]\[20\] net772 net766 datapath.rf.registers\[24\]\[20\]
+ _02372_ vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__a221o_1
XFILLER_139_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout616_X net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10550_ keypad.debounce.debounce\[13\] keypad.debounce.debounce\[12\] keypad.debounce.debounce\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05377_ sky130_fd_sc_hd__and3_1
XANTENNA__07285__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07824__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06881__X _01717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09209_ net649 _04044_ net439 vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__a21o_1
X_10481_ screen.controlBus\[21\] screen.controlBus\[20\] screen.controlBus\[23\] screen.controlBus\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05311_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_20_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12220_ net2148 _06221_ net602 vssd1 vssd1 vccd1 vccd1 _06224_ sky130_fd_sc_hd__o21ai_1
XFILLER_6_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11659__B _05874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06760__C net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08785__A0 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12151_ net1606 _06180_ _06181_ vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__o21a_1
XFILLER_150_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11102_ net183 net1819 net534 vssd1 vssd1 vccd1 vccd1 _00159_ sky130_fd_sc_hd__mux2_1
X_12082_ screen.register.currentYbus\[22\] _05837_ _06018_ screen.register.currentYbus\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06121_ sky130_fd_sc_hd__a22o_1
Xhold690 datapath.rf.registers\[9\]\[30\] vssd1 vssd1 vccd1 vccd1 net2038 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08968__B net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11033_ net181 net2198 net539 vssd1 vssd1 vccd1 vccd1 _00095_ sky130_fd_sc_hd__mux2_1
XANTENNA__06769__A _01571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12984_ net210 net2616 net478 vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__mux2_1
X_11935_ net2564 net162 vssd1 vssd1 vccd1 vccd1 _05987_ sky130_fd_sc_hd__nand2_1
XFILLER_33_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14654_ clknet_leaf_149_clk _01359_ net1061 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_28_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11866_ net2550 net163 vssd1 vssd1 vccd1 vccd1 _05941_ sky130_fd_sc_hd__nand2_1
X_13605_ clknet_leaf_139_clk _00415_ net1099 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06935__C _01656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10817_ _01480_ net655 _05573_ _05574_ vssd1 vssd1 vccd1 vccd1 _05575_ sky130_fd_sc_hd__o22a_2
X_14585_ clknet_leaf_31_clk _01290_ net1122 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08068__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11797_ datapath.ru.latched_instruction\[3\] net334 net314 _01461_ vssd1 vssd1 vccd1
+ vccd1 _00663_ sky130_fd_sc_hd__a22o_1
XFILLER_13_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13536_ clknet_leaf_137_clk _00346_ net1090 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10748_ _05513_ _05514_ vssd1 vssd1 vccd1 vccd1 _05515_ sky130_fd_sc_hd__or2_1
X_13467_ clknet_leaf_37_clk _00277_ net1138 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10679_ _05428_ _05494_ _05482_ vssd1 vssd1 vccd1 vccd1 _05497_ sky130_fd_sc_hd__o21a_1
XANTENNA__10754__A net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06951__B net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12418_ net1419 net131 _06356_ vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__a21o_1
XANTENNA__09568__A2 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13398_ clknet_leaf_140_clk _00208_ net1093 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_127_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12349_ net638 _04624_ _06315_ vssd1 vssd1 vccd1 vccd1 _06316_ sky130_fd_sc_hd__a21oi_1
XFILLER_5_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08528__B1 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14019_ clknet_leaf_80_clk _00788_ net1254 vssd1 vssd1 vccd1 vccd1 datapath.PC\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_06910_ net974 net919 vssd1 vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__and2_1
XFILLER_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07890_ net613 _02725_ net564 vssd1 vssd1 vccd1 vccd1 _02726_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07200__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06841_ datapath.ru.latched_instruction\[15\] _01510_ net1015 vssd1 vssd1 vccd1 vccd1
+ _01677_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09560_ _04393_ _04394_ _04338_ vssd1 vssd1 vccd1 vccd1 _04396_ sky130_fd_sc_hd__a21bo_1
XFILLER_110_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06772_ _01575_ _01607_ vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__or2_2
XFILLER_83_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06966__X _01802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08511_ datapath.rf.registers\[26\]\[1\] net781 net716 datapath.rf.registers\[4\]\[1\]
+ _03346_ vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__a221o_1
XANTENNA__09342__X _04178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09491_ net376 _04321_ _04326_ net379 vssd1 vssd1 vccd1 vccd1 _04327_ sky130_fd_sc_hd__a31o_1
X_08442_ datapath.rf.registers\[9\]\[2\] net705 _03269_ _03271_ _03272_ vssd1 vssd1
+ vccd1 vccd1 _03278_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_156_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_max_cap950_X net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08373_ datapath.rf.registers\[29\]\[3\] net677 net670 datapath.rf.registers\[21\]\[3\]
+ _03208_ vssd1 vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_156_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout144_A net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07324_ datapath.rf.registers\[14\]\[24\] net831 net799 datapath.rf.registers\[15\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__a22o_1
XANTENNA__07797__X _02633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07806__A2 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07255_ net612 _02090_ net564 vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__a21oi_4
XANTENNA_fanout1053_A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout409_A _05733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07186_ datapath.rf.registers\[8\]\[27\] net877 net800 datapath.rf.registers\[15\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__a22o_1
XFILLER_105_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08231__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout680_A _01828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout400 net401 vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__clkbuf_8
Xfanout411 _05730_ vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__buf_4
XANTENNA__08788__B net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout422 net425 vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__buf_6
XANTENNA_fanout778_A _01794_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout399_X net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_6_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout433 _05711_ vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__buf_4
Xfanout444 net445 vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__clkbuf_4
Xfanout455 net456 vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__buf_1
Xfanout466 _01701_ vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__clkbuf_4
X_09827_ net608 _04646_ _04662_ net556 vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__o211a_1
Xfanout477 _06559_ vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_107_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout488 _06552_ vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout566_X net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout945_A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout499 net501 vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__buf_2
X_09758_ net337 _04553_ vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__nor2_1
XFILLER_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08709_ _03263_ _03296_ vssd1 vssd1 vccd1 vccd1 _03545_ sky130_fd_sc_hd__nor2_1
XANTENNA__11942__B screen.counter.ack vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09689_ _04259_ _04440_ net373 vssd1 vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout733_X net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11434__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ net6 net1034 net1024 net1453 vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_120_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11651_ keypad.decode.sticky_n\[2\] keypad.decode.sticky_n\[3\] _05873_ vssd1 vssd1
+ vccd1 vccd1 _05874_ sky130_fd_sc_hd__nor3_4
X_10602_ screen.register.currentYbus\[25\] screen.register.currentYbus\[24\] screen.register.currentYbus\[27\]
+ screen.register.currentYbus\[26\] vssd1 vssd1 vccd1 vccd1 _05423_ sky130_fd_sc_hd__or4_1
X_14370_ clknet_leaf_151_clk _01075_ net1052 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11582_ screen.counter.ct\[4\] screen.counter.ct\[5\] vssd1 vssd1 vccd1 vccd1 _05806_
+ sky130_fd_sc_hd__nand2_2
XFILLER_156_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13321_ clknet_leaf_62_clk _00131_ net1234 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10533_ _05351_ _05353_ _05356_ _05360_ _05362_ vssd1 vssd1 vccd1 vccd1 _05363_ sky130_fd_sc_hd__o2111a_1
XANTENNA__10574__A _03009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08470__A2 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06771__B _01607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12003__B1 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13252_ clknet_leaf_22_clk _00062_ net1156 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_118_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10464_ _05292_ _05293_ vssd1 vssd1 vccd1 vccd1 _05294_ sky130_fd_sc_hd__or2_1
XANTENNA__08044__A _02856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12203_ net1523 _06210_ _06212_ vssd1 vssd1 vccd1 vccd1 _00762_ sky130_fd_sc_hd__a21oi_1
X_13183_ net2520 vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08222__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10395_ _03612_ net575 vssd1 vssd1 vccd1 vccd1 _05231_ sky130_fd_sc_hd__nand2_1
XFILLER_135_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07430__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12134_ _06168_ net601 vssd1 vssd1 vccd1 vccd1 _06171_ sky130_fd_sc_hd__nor2_1
XFILLER_89_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13096__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09707__C1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12065_ _05806_ _05856_ _05860_ _05846_ vssd1 vssd1 vccd1 vccd1 _06105_ sky130_fd_sc_hd__a211o_1
X_11016_ net265 net2309 net541 vssd1 vssd1 vccd1 vccd1 _00078_ sky130_fd_sc_hd__mux2_1
XFILLER_37_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11817__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12967_ net295 net2143 net478 vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__mux2_1
XANTENNA__13437__RESET_B net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11344__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11918_ _02385_ net656 vssd1 vssd1 vccd1 vccd1 _05976_ sky130_fd_sc_hd__nand2_1
X_12898_ net1909 net288 net485 vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__mux2_1
X_11849_ _05336_ _05919_ _05922_ _05343_ vssd1 vssd1 vccd1 vccd1 _05928_ sky130_fd_sc_hd__a2bb2o_1
X_14637_ clknet_leaf_125_clk _01342_ net1205 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09238__A1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07249__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14568_ clknet_leaf_59_clk _01273_ net1235 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06962__A net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13519_ clknet_leaf_27_clk _00329_ net1133 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_14499_ clknet_leaf_120_clk _01204_ net1193 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08461__A2 _03294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload10 clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clkload10/Y sky130_fd_sc_hd__inv_6
Xclkload21 clknet_leaf_149_clk vssd1 vssd1 vccd1 vccd1 clkload21/Y sky130_fd_sc_hd__clkinv_4
X_07040_ datapath.rf.registers\[23\]\[30\] net941 net925 vssd1 vssd1 vccd1 vccd1 _01876_
+ sky130_fd_sc_hd__and3_1
Xclkload32 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 clkload32/Y sky130_fd_sc_hd__clkinv_2
Xclkload43 clknet_leaf_145_clk vssd1 vssd1 vccd1 vccd1 clkload43/Y sky130_fd_sc_hd__bufinv_16
Xclkload54 clknet_leaf_135_clk vssd1 vssd1 vccd1 vccd1 clkload54/Y sky130_fd_sc_hd__bufinv_16
Xclkload65 clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 clkload65/Y sky130_fd_sc_hd__inv_8
Xclkload76 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 clkload76/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__10771__X _05536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload87 clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 clkload87/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__08213__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12903__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload98 clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 clkload98/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__07421__B1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08991_ _03822_ _03826_ vssd1 vssd1 vccd1 vccd1 _03827_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_10_Left_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07942_ datapath.rf.registers\[29\]\[11\] net979 net918 vssd1 vssd1 vccd1 vccd1 _02778_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08401__B net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07873_ datapath.rf.registers\[12\]\[13\] net755 net660 datapath.rf.registers\[5\]\[13\]
+ _02708_ vssd1 vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__a221o_1
X_09612_ net905 _03558_ net627 _03542_ _04447_ vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__a221o_1
X_06824_ net1029 _01659_ vssd1 vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__nor2_1
XANTENNA__13860__RESET_B net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09543_ _04377_ _04378_ net366 vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__mux2_1
XANTENNA__09513__A _02704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06755_ net652 vssd1 vssd1 vccd1 vccd1 MemRead sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_69_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08134__D1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11254__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07488__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09474_ net463 net452 _04304_ net460 vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__o211a_1
X_06686_ datapath.ru.latched_instruction\[16\] _01524_ vssd1 vssd1 vccd1 vccd1 _01525_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_52_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08425_ _03251_ _03256_ _03260_ vssd1 vssd1 vccd1 vccd1 _03261_ sky130_fd_sc_hd__or3_2
XFILLER_12_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout526_A _05721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout147_X net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1170_A net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08356_ datapath.rf.registers\[20\]\[3\] net840 net792 datapath.rf.registers\[18\]\[3\]
+ _03183_ vssd1 vssd1 vccd1 vccd1 _03192_ sky130_fd_sc_hd__a221o_1
XANTENNA__06872__A _01656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload4 clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clkload4/Y sky130_fd_sc_hd__clkinvlp_4
X_07307_ _02129_ _02131_ _02141_ _02142_ vssd1 vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__or4_1
XFILLER_138_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08287_ _03114_ _03118_ _03122_ net784 datapath.rf.registers\[0\]\[5\] vssd1 vssd1
+ vccd1 vccd1 _03123_ sky130_fd_sc_hd__o32a_4
XFILLER_50_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08452__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07238_ datapath.rf.registers\[4\]\[26\] net714 net679 datapath.rf.registers\[6\]\[26\]
+ _02073_ vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout895_A net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07169_ datapath.rf.registers\[2\]\[27\] net888 net846 datapath.rf.registers\[1\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__a22o_1
XANTENNA__12813__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10180_ _04831_ _04881_ vssd1 vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout683_X net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11429__S net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1206 net1213 vssd1 vssd1 vccd1 vccd1 net1206 sky130_fd_sc_hd__clkbuf_2
Xfanout1217 net1262 vssd1 vssd1 vccd1 vccd1 net1217 sky130_fd_sc_hd__buf_2
Xfanout230 _04712_ vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__clkbuf_4
Xfanout1228 net1230 vssd1 vssd1 vccd1 vccd1 net1228 sky130_fd_sc_hd__clkbuf_4
Xfanout241 net242 vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__clkbuf_2
XFILLER_87_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1239 net1240 vssd1 vssd1 vccd1 vccd1 net1239 sky130_fd_sc_hd__clkbuf_4
Xfanout252 _05588_ vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_89_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout850_X net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout263 _05575_ vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_89_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout274 net277 vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__clkbuf_2
Xfanout285 _05547_ vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout948_X net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout296 net297 vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__clkbuf_2
X_13870_ clknet_leaf_75_clk _00674_ net1247 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07191__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12821_ net1813 net201 net491 vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__mux2_1
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11164__S net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07479__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12752_ net2370 net215 net402 vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__mux2_1
XANTENNA__12472__B1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11814__A3 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11703_ mmio.wishbone.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1 _05887_ sky130_fd_sc_hd__and2_1
X_12683_ net2595 net503 net499 _06516_ vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__a22o_1
XANTENNA__10856__X _05608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14422_ clknet_leaf_140_clk _01127_ net1094 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_11634_ net998 _05857_ vssd1 vssd1 vccd1 vccd1 _05858_ sky130_fd_sc_hd__nor2_1
XANTENNA__06782__A _01614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14353_ clknet_leaf_40_clk _01058_ net1140 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11565_ net1009 _05777_ vssd1 vssd1 vccd1 vccd1 _05789_ sky130_fd_sc_hd__nor2_1
XANTENNA__08443__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13304_ clknet_leaf_6_clk _00114_ net1067 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10516_ _05344_ _05345_ vssd1 vssd1 vccd1 vccd1 _05346_ sky130_fd_sc_hd__nand2_1
XFILLER_144_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14284_ clknet_leaf_133_clk _00989_ net1105 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_109_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11496_ net218 net2062 net510 vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__mux2_1
XFILLER_6_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13235_ clknet_leaf_34_clk _00045_ net1128 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10447_ _05240_ _05270_ _05211_ vssd1 vssd1 vccd1 vccd1 _05283_ sky130_fd_sc_hd__or3b_1
XFILLER_3_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13166_ datapath.rf.registers\[0\]\[3\] vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__clkbuf_1
XFILLER_112_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10378_ _01859_ _04705_ vssd1 vssd1 vccd1 vccd1 _05214_ sky130_fd_sc_hd__nand2_1
XFILLER_112_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06757__A2 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11339__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12117_ _05780_ _05806_ vssd1 vssd1 vccd1 vccd1 _06154_ sky130_fd_sc_hd__nor2_1
XANTENNA__12317__A2_N _06253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13097_ net286 net1642 net472 vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__mux2_1
X_12048_ _05775_ _05852_ _05847_ vssd1 vssd1 vccd1 vccd1 _06089_ sky130_fd_sc_hd__o21a_1
XFILLER_38_615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07706__A1 datapath.rf.registers\[0\]\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06957__A _01637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07182__A2 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13999_ clknet_leaf_113_clk _00776_ net1195 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11074__S net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08210_ datapath.rf.registers\[1\]\[6\] net845 net829 datapath.rf.registers\[14\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03046_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_16_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07890__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09190_ _03584_ _04024_ vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__nand2_1
XFILLER_147_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10485__Y _05315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08141_ datapath.rf.registers\[14\]\[8\] net777 net745 datapath.rf.registers\[2\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02977_ sky130_fd_sc_hd__a22o_1
XANTENNA__10777__B1 _05539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload110 clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 clkload110/Y sky130_fd_sc_hd__inv_6
XANTENNA__07642__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08072_ datapath.rf.registers\[14\]\[9\] net830 net812 datapath.rf.registers\[13\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02908_ sky130_fd_sc_hd__a22o_1
Xclkload121 clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 clkload121/X sky130_fd_sc_hd__clkbuf_8
Xclkload132 clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 clkload132/Y sky130_fd_sc_hd__inv_8
Xclkload143 clknet_leaf_79_clk vssd1 vssd1 vccd1 vccd1 clkload143/Y sky130_fd_sc_hd__inv_8
XANTENNA__10364__D _05199_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07023_ _01857_ _01858_ vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__or2_2
XFILLER_136_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06748__A2 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11741__A2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11249__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08974_ _03263_ _03320_ net446 vssd1 vssd1 vccd1 vccd1 _03810_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1016_A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold16 keypad.debounce.debounce\[3\] vssd1 vssd1 vccd1 vccd1 net1364 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold27 datapath.ru.n_memread vssd1 vssd1 vccd1 vccd1 net1375 sky130_fd_sc_hd__dlygate4sd3_1
X_07925_ datapath.rf.registers\[26\]\[12\] net781 net729 datapath.rf.registers\[25\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02761_ sky130_fd_sc_hd__a22o_1
Xhold38 screen.controlBus\[21\] vssd1 vssd1 vccd1 vccd1 net1386 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07158__C1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold49 net69 vssd1 vssd1 vccd1 vccd1 net1397 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout476_A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07856_ datapath.rf.registers\[16\]\[13\] net861 net833 datapath.rf.registers\[30\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__a22o_1
XFILLER_84_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07173__A2 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08370__B2 _01647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06807_ datapath.ru.latched_instruction\[7\] net1028 net993 _01642_ vssd1 vssd1 vccd1
+ vccd1 _01643_ sky130_fd_sc_hd__a22oi_4
XFILLER_45_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10797__A2_N _05556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07787_ datapath.rf.registers\[17\]\[15\] net747 net676 datapath.rf.registers\[29\]\[15\]
+ _02622_ vssd1 vssd1 vccd1 vccd1 _02623_ sky130_fd_sc_hd__a221o_1
XFILLER_25_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09526_ net360 _04361_ vssd1 vssd1 vccd1 vccd1 _04362_ sky130_fd_sc_hd__nand2_1
X_06738_ datapath.ru.latched_instruction\[6\] net1028 vssd1 vssd1 vccd1 vccd1 _01577_
+ sky130_fd_sc_hd__and2_1
XFILLER_52_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09457_ net379 _03838_ _04287_ _04292_ _03614_ vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__a221o_1
XANTENNA__07969__Y _02805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06669_ _01409_ _01502_ _01507_ vssd1 vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__a21bo_1
XFILLER_40_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout810_A net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout431_X net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12808__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout529_X net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08408_ datapath.rf.registers\[8\]\[2\] net956 _01712_ vssd1 vssd1 vccd1 vccd1 _03244_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07881__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09388_ net650 _04223_ net439 vssd1 vssd1 vccd1 vccd1 _04224_ sky130_fd_sc_hd__a21oi_1
X_08339_ datapath.rf.registers\[4\]\[3\] net960 net936 vssd1 vssd1 vccd1 vccd1 _03175_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07633__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11350_ net284 net1893 net520 vssd1 vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_115_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10301_ datapath.PC\[12\] net467 vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__or2_1
XANTENNA__11948__A _01908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11281_ net282 net1988 net524 vssd1 vssd1 vccd1 vccd1 _00329_ sky130_fd_sc_hd__mux2_1
XFILLER_106_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13020_ net1603 net197 net392 vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__mux2_1
XFILLER_4_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10232_ net638 _04626_ _05067_ _05066_ net224 vssd1 vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__a311o_1
XFILLER_152_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10571__B _02856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07936__A1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11159__S net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10163_ net890 _04585_ vssd1 vssd1 vccd1 vccd1 _04999_ sky130_fd_sc_hd__nor2_1
Xfanout1003 net1004 vssd1 vssd1 vccd1 vccd1 net1003 sky130_fd_sc_hd__clkbuf_2
XFILLER_79_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1014 net1015 vssd1 vssd1 vccd1 vccd1 net1014 sky130_fd_sc_hd__buf_2
XANTENNA__08041__B _01784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1025 _05889_ vssd1 vssd1 vccd1 vccd1 net1025 sky130_fd_sc_hd__buf_2
Xfanout1036 _05887_ vssd1 vssd1 vccd1 vccd1 net1036 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input37_A gpio_in[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10094_ _04882_ _04884_ vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__or2_1
XANTENNA__10998__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1058 net1121 vssd1 vssd1 vccd1 vccd1 net1058 sky130_fd_sc_hd__clkbuf_2
Xfanout1069 net1075 vssd1 vssd1 vccd1 vccd1 net1069 sky130_fd_sc_hd__clkbuf_4
X_13922_ clknet_leaf_109_clk _00700_ net1220 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06777__A _01613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13853_ clknet_leaf_49_clk _00657_ net1177 vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__dfrtp_1
XFILLER_63_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06911__A2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12804_ net1870 net284 net492 vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__mux2_1
X_13784_ clknet_leaf_52_clk _00593_ net1181 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10996_ net2311 net185 net434 vssd1 vssd1 vccd1 vccd1 _00061_ sky130_fd_sc_hd__mux2_1
XFILLER_90_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12735_ net1708 net300 net402 vssd1 vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__mux2_1
XFILLER_30_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06783__Y _01620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12666_ datapath.mulitply_result\[26\] datapath.multiplication_module.multiplicand_i\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06502_ sky130_fd_sc_hd__nand2_1
XANTENNA__07872__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11617_ _05294_ _05760_ _05762_ _05838_ net1006 vssd1 vssd1 vccd1 vccd1 _05841_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_13_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14405_ clknet_leaf_117_clk _01110_ net1190 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08416__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12597_ _06442_ _06443_ vssd1 vssd1 vccd1 vccd1 _06445_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11548_ net1009 _05770_ vssd1 vssd1 vccd1 vccd1 _05772_ sky130_fd_sc_hd__nor2_4
X_14336_ clknet_leaf_136_clk _01041_ net1088 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_144_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11858__A _03417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold508 datapath.rf.registers\[6\]\[15\] vssd1 vssd1 vccd1 vccd1 net1856 sky130_fd_sc_hd__dlygate4sd3_1
X_14267_ clknet_leaf_45_clk _00972_ net1146 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold519 datapath.rf.registers\[24\]\[16\] vssd1 vssd1 vccd1 vccd1 net1867 sky130_fd_sc_hd__dlygate4sd3_1
X_11479_ net258 net1550 net513 vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__mux2_1
XFILLER_143_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13218_ clknet_leaf_150_clk _00028_ net1053 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_98_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14198_ clknet_leaf_66_clk datapath.multiplication_module.multiplicand_i_n\[9\] net1237
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[9\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11069__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11723__A2 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13149_ net1887 net216 net382 vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__mux2_1
XFILLER_32_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1208 screen.register.currentYbus\[25\] vssd1 vssd1 vccd1 vccd1 net2556 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1219 datapath.rf.registers\[25\]\[26\] vssd1 vssd1 vccd1 vccd1 net2567 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07710_ datapath.rf.registers\[4\]\[16\] net957 net931 vssd1 vssd1 vccd1 vccd1 _02546_
+ sky130_fd_sc_hd__and3_1
XFILLER_111_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08690_ _02705_ _02726_ vssd1 vssd1 vccd1 vccd1 _03526_ sky130_fd_sc_hd__nor2_1
XANTENNA__07155__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07641_ datapath.rf.registers\[31\]\[18\] net687 net664 datapath.rf.registers\[15\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__a22o_1
XFILLER_25_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07572_ datapath.rf.registers\[30\]\[19\] net834 _02391_ _02402_ _02403_ vssd1 vssd1
+ vccd1 vccd1 _02408_ sky130_fd_sc_hd__a2111o_1
X_09311_ _03447_ _03518_ vssd1 vssd1 vccd1 vccd1 _04147_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09242_ _02364_ _02386_ net624 vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__o21a_1
XANTENNA__07863__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07949__C net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07311__A _02125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09173_ _04008_ vssd1 vssd1 vccd1 vccd1 _04009_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout224_A net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08124_ _02950_ net584 datapath.rf.registers\[0\]\[8\] net867 vssd1 vssd1 vccd1 vccd1
+ _02960_ sky130_fd_sc_hd__o2bb2a_4
XANTENNA__07615__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07030__B net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08055_ datapath.rf.registers\[7\]\[9\] net941 net934 vssd1 vssd1 vccd1 vccd1 _02891_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1133_A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07006_ datapath.rf.registers\[24\]\[31\] net767 net692 datapath.rf.registers\[13\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01842_ sky130_fd_sc_hd__a22o_1
XFILLER_89_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11714__A2 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08040__B1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07394__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08957_ _03792_ vssd1 vssd1 vccd1 vccd1 _03793_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout760_A _01802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08328__D1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout479_X net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout858_A net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07908_ datapath.rf.registers\[4\]\[12\] net865 net840 datapath.rf.registers\[20\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__a22o_1
XANTENNA__06597__A net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08888_ _03665_ _03668_ net317 _03715_ vssd1 vssd1 vccd1 vccd1 _03724_ sky130_fd_sc_hd__o22a_1
XANTENNA__09540__A0 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07146__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07839_ datapath.rf.registers\[26\]\[14\] net779 _02674_ net787 vssd1 vssd1 vccd1
+ vccd1 _02675_ sky130_fd_sc_hd__a211o_1
XANTENNA__10150__A1 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10850_ _04146_ _05602_ net902 vssd1 vssd1 vccd1 vccd1 _05603_ sky130_fd_sc_hd__mux2_2
XANTENNA__06884__X _01720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09509_ net464 _03149_ net452 vssd1 vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout813_X net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10781_ _05542_ _05543_ vssd1 vssd1 vccd1 vccd1 _05544_ sky130_fd_sc_hd__nor2_1
X_12520_ datapath.mulitply_result\[2\] datapath.multiplication_module.multiplicand_i\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06380_ sky130_fd_sc_hd__and2_1
XANTENNA__07854__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_117_Right_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12451_ net165 _05950_ net127 net2648 vssd1 vssd1 vccd1 vccd1 _00853_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_12_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11402_ net1557 net198 net412 vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__mux2_1
X_12382_ net2636 net133 _06338_ vssd1 vssd1 vccd1 vccd1 _00815_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_97_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14121_ clknet_leaf_60_clk _00878_ net1169 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11333_ net1777 net200 net415 vssd1 vssd1 vccd1 vccd1 _00378_ sky130_fd_sc_hd__mux2_1
XFILLER_4_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09359__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14052_ clknet_leaf_100_clk _00819_ net1228 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11264_ net204 net2417 net418 vssd1 vssd1 vccd1 vccd1 _00313_ sky130_fd_sc_hd__mux2_1
X_13003_ net1762 net278 net393 vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__mux2_1
X_10215_ _05019_ _05031_ _05041_ _05050_ vssd1 vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__or4_1
XANTENNA__08031__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11195_ net215 net2244 net422 vssd1 vssd1 vccd1 vccd1 _00247_ sky130_fd_sc_hd__mux2_1
XFILLER_79_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07385__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07891__A _02704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10146_ net637 _04624_ _04928_ _04606_ vssd1 vssd1 vccd1 vccd1 _04982_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_128_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10077_ datapath.PC\[30\] _03751_ vssd1 vssd1 vccd1 vccd1 _04913_ sky130_fd_sc_hd__and2_1
XANTENNA__12302__A net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07137__A2 _01756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09531__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13905_ clknet_leaf_43_clk net1359 net1149 vssd1 vssd1 vccd1 vccd1 keypad.debounce.debounce\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_63_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload2_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06794__X _01630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13836_ clknet_leaf_113_clk _00645_ net1197 vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__dfrtp_1
XFILLER_35_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13767_ clknet_leaf_81_clk _00576_ net1255 vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__dfrtp_1
X_10979_ net1665 net271 net436 vssd1 vssd1 vccd1 vccd1 _00044_ sky130_fd_sc_hd__mux2_1
XANTENNA__11352__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07402__Y _02238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12718_ columns.count\[7\] columns.count\[6\] _06538_ vssd1 vssd1 vccd1 vccd1 _06541_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07845__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13698_ clknet_leaf_151_clk _00508_ net1053 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_44_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12649_ _06486_ _06487_ vssd1 vssd1 vccd1 vccd1 _06488_ sky130_fd_sc_hd__or2_1
XANTENNA__06970__A _01800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07073__A1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold305 datapath.rf.registers\[8\]\[17\] vssd1 vssd1 vccd1 vccd1 net1653 sky130_fd_sc_hd__dlygate4sd3_1
X_14319_ clknet_leaf_27_clk _01024_ net1133 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08270__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold316 datapath.rf.registers\[21\]\[24\] vssd1 vssd1 vccd1 vccd1 net1664 sky130_fd_sc_hd__dlygate4sd3_1
Xhold327 datapath.rf.registers\[20\]\[30\] vssd1 vssd1 vccd1 vccd1 net1675 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_wire561_A _02568_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold338 datapath.rf.registers\[5\]\[2\] vssd1 vssd1 vccd1 vccd1 net1686 sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 datapath.rf.registers\[3\]\[10\] vssd1 vssd1 vccd1 vccd1 net1697 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout807 net809 vssd1 vssd1 vccd1 vccd1 net807 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08022__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09860_ _03231_ _03298_ _04695_ _03230_ vssd1 vssd1 vccd1 vccd1 _04696_ sky130_fd_sc_hd__o31a_1
XANTENNA__12911__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout818 _01758_ vssd1 vssd1 vccd1 vccd1 net818 sky130_fd_sc_hd__clkbuf_8
Xfanout829 net831 vssd1 vssd1 vccd1 vccd1 net829 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07376__A2 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09770__B1 _03978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08811_ _03228_ _03644_ _03645_ vssd1 vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__o21ai_1
X_09791_ _01957_ _03471_ vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__and2b_1
XANTENNA__10380__A1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1005 datapath.rf.registers\[15\]\[10\] vssd1 vssd1 vccd1 vccd1 net2353 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1016 datapath.multiplication_module.multiplicand_i\[2\] vssd1 vssd1 vccd1 vccd1
+ net2364 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1027 datapath.rf.registers\[2\]\[19\] vssd1 vssd1 vccd1 vccd1 net2375 sky130_fd_sc_hd__dlygate4sd3_1
X_08742_ _03518_ _03521_ _03576_ _03517_ vssd1 vssd1 vccd1 vccd1 _03578_ sky130_fd_sc_hd__a31o_1
Xhold1038 datapath.rf.registers\[10\]\[10\] vssd1 vssd1 vccd1 vccd1 net2386 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 datapath.rf.registers\[21\]\[11\] vssd1 vssd1 vccd1 vccd1 net2397 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_916 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08673_ _02419_ _02440_ vssd1 vssd1 vccd1 vccd1 _03509_ sky130_fd_sc_hd__nor2_1
XANTENNA__10132__A1 _01702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout174_A _05684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07624_ datapath.rf.registers\[2\]\[18\] net887 _02449_ _02452_ _02459_ vssd1 vssd1
+ vccd1 vccd1 _02460_ sky130_fd_sc_hd__a2111oi_1
XTAP_TAPCELL_ROW_37_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07025__B net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11880__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08089__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07555_ datapath.rf.registers\[27\]\[19\] net977 net938 vssd1 vssd1 vccd1 vccd1 _02391_
+ sky130_fd_sc_hd__and3_1
XFILLER_81_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11262__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1083_A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07836__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07486_ datapath.rf.registers\[17\]\[21\] net746 net722 datapath.rf.registers\[18\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__a22o_1
XANTENNA__07300__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09225_ net372 _03766_ _03627_ net377 vssd1 vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__a211o_1
XFILLER_22_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1250_A net1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout227_X net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09156_ net461 _03926_ _03927_ vssd1 vssd1 vccd1 vccd1 _03992_ sky130_fd_sc_hd__nand3_1
XANTENNA__06880__A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_726 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08107_ datapath.rf.registers\[24\]\[8\] net858 net791 datapath.rf.registers\[18\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__a22o_1
X_09087_ net372 _03766_ _03922_ vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__o21a_1
XFILLER_135_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_110_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_110_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_2_Left_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08038_ datapath.rf.registers\[3\]\[10\] net772 net764 datapath.rf.registers\[1\]\[10\]
+ _02860_ vssd1 vssd1 vccd1 vccd1 _02874_ sky130_fd_sc_hd__a221o_1
Xhold850 datapath.rf.registers\[27\]\[29\] vssd1 vssd1 vccd1 vccd1 net2198 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold861 datapath.rf.registers\[20\]\[6\] vssd1 vssd1 vccd1 vccd1 net2209 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout975_A net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout596_X net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold872 datapath.rf.registers\[3\]\[24\] vssd1 vssd1 vccd1 vccd1 net2220 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12821__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold883 datapath.rf.registers\[10\]\[19\] vssd1 vssd1 vccd1 vccd1 net2231 sky130_fd_sc_hd__dlygate4sd3_1
Xhold894 datapath.rf.registers\[23\]\[26\] vssd1 vssd1 vccd1 vccd1 net2242 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06879__X _01715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07367__A2 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10000_ _04771_ _04792_ vssd1 vssd1 vccd1 vccd1 _04836_ sky130_fd_sc_hd__xor2_1
XFILLER_49_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09989_ net1263 net594 vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout763_X net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10371__A1 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11437__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07119__A2 _01954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10123__A1 _03729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11951_ _01854_ screen.counter.ack vssd1 vssd1 vccd1 vccd1 _05998_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout930_X net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10902_ net1264 datapath.PC\[25\] _05636_ vssd1 vssd1 vccd1 vccd1 _05647_ sky130_fd_sc_hd__and3_1
X_14670_ clknet_leaf_0_clk _01375_ net1055 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11871__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11882_ _02980_ net658 vssd1 vssd1 vccd1 vccd1 _05952_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_123_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10833_ net251 net2588 net542 vssd1 vssd1 vccd1 vccd1 _00016_ sky130_fd_sc_hd__mux2_1
X_13621_ clknet_leaf_127_clk _00431_ net1211 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_25_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10577__A _02025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11172__S net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07827__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10764_ net301 net2276 net544 vssd1 vssd1 vccd1 vccd1 _00006_ sky130_fd_sc_hd__mux2_1
X_13552_ clknet_leaf_24_clk _00362_ net1155 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_12503_ net196 net2132 net507 vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__mux2_1
X_13483_ clknet_leaf_47_clk _00293_ net1174 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10695_ net1444 _03417_ net570 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i_n\[0\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_145_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12434_ net1412 net131 _06364_ vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__a21o_1
XFILLER_138_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08334__X _03170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13099__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12365_ _05680_ _06254_ _06327_ net190 vssd1 vssd1 vccd1 vccd1 _06328_ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_101_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_101_clk
+ sky130_fd_sc_hd__clkbuf_8
X_14104_ clknet_leaf_95_clk _00870_ net1217 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_11316_ net1605 net282 net416 vssd1 vssd1 vccd1 vccd1 _00361_ sky130_fd_sc_hd__mux2_1
X_12296_ _04300_ _06277_ net890 vssd1 vssd1 vccd1 vccd1 _06278_ sky130_fd_sc_hd__mux2_1
XFILLER_99_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14035_ clknet_leaf_84_clk _00804_ net1259 vssd1 vssd1 vccd1 vccd1 datapath.PC\[25\]
+ sky130_fd_sc_hd__dfstp_2
X_11247_ net293 net2184 net418 vssd1 vssd1 vccd1 vccd1 _00296_ sky130_fd_sc_hd__mux2_1
XANTENNA__08004__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12731__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07358__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11178_ net299 net2235 net423 vssd1 vssd1 vccd1 vccd1 _00230_ sky130_fd_sc_hd__mux2_1
XFILLER_121_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10362__A1 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11347__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06949__B _01784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10129_ _04954_ _04964_ vssd1 vssd1 vccd1 vccd1 _04965_ sky130_fd_sc_hd__nand2_1
XANTENNA__09504__A0 _02912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12103__A2 _05773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06965__A net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07530__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13819_ clknet_leaf_115_clk _00628_ net1189 vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__dfrtp_1
XFILLER_51_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09807__A1 _03607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11082__S net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07340_ datapath.rf.registers\[4\]\[24\] net715 net707 datapath.rf.registers\[10\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__a22o_1
XANTENNA__07818__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07499__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07271_ datapath.rf.registers\[15\]\[25\] net987 net916 vssd1 vssd1 vccd1 vccd1 _02107_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12906__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap659_X net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09010_ _03295_ _03644_ net458 _03659_ _03648_ vssd1 vssd1 vccd1 vccd1 _03846_ sky130_fd_sc_hd__o221ai_4
XFILLER_145_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold102 datapath.multiplication_module.multiplier_i\[2\] vssd1 vssd1 vccd1 vccd1
+ net1450 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold113 net102 vssd1 vssd1 vccd1 vccd1 net1461 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08404__B net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold124 mmio.key_data\[5\] vssd1 vssd1 vccd1 vccd1 net1472 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07597__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold135 keypad.decode.sticky\[1\] vssd1 vssd1 vccd1 vccd1 net1483 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold146 net78 vssd1 vssd1 vccd1 vccd1 net1494 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 datapath.multiplication_module.multiplier_i\[9\] vssd1 vssd1 vccd1 vccd1
+ net1505 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 datapath.multiplication_module.multiplicand_i\[23\] vssd1 vssd1 vccd1 vccd1
+ net1516 sky130_fd_sc_hd__dlygate4sd3_1
X_09912_ datapath.PC\[13\] net604 _04747_ vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__or3_2
Xhold179 screen.controlBus\[4\] vssd1 vssd1 vccd1 vccd1 net1527 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_74_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout604 _04727_ vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__buf_2
Xfanout615 net616 vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__buf_4
Xfanout626 net629 vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__clkbuf_4
Xfanout637 net639 vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__buf_2
X_09843_ _01859_ _01911_ vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__nand2_1
Xfanout648 net650 vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__buf_2
XANTENNA__11257__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06986_ net969 net911 net908 vssd1 vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__and3_1
X_09774_ _03494_ _03591_ _03492_ vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__a21oi_1
X_08725_ _03080_ _03081_ vssd1 vssd1 vccd1 vccd1 _03561_ sky130_fd_sc_hd__nand2b_2
XANTENNA__10949__X _05688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ _02092_ _02094_ vssd1 vssd1 vccd1 vccd1 _03492_ sky130_fd_sc_hd__nand2_2
XFILLER_82_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06875__A _01630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07521__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_54_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07607_ _02442_ vssd1 vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_105_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08587_ _03297_ _03360_ _03421_ _03298_ vssd1 vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__a31o_2
XANTENNA_fanout723_A net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07809__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07538_ datapath.rf.registers\[17\]\[20\] net746 net742 datapath.rf.registers\[2\]\[20\]
+ _02373_ vssd1 vssd1 vccd1 vccd1 _02374_ sky130_fd_sc_hd__a221o_1
XFILLER_149_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout511_X net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07469_ datapath.rf.registers\[20\]\[21\] net839 net824 datapath.rf.registers\[6\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02305_ sky130_fd_sc_hd__a22o_1
XANTENNA__12816__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_69_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout609_X net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09208_ net345 _04043_ vssd1 vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__or2_1
X_10480_ _05308_ _05309_ vssd1 vssd1 vccd1 vccd1 _05310_ sky130_fd_sc_hd__nor2_1
XFILLER_6_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_112_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09139_ _01620_ _03951_ _03974_ net318 _03973_ vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__o221a_1
XANTENNA__08234__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08785__A1 _03228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07588__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12150_ net1279 _06180_ _06178_ vssd1 vssd1 vccd1 vccd1 _06181_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout880_X net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11101_ net176 net1695 net534 vssd1 vssd1 vccd1 vccd1 _00158_ sky130_fd_sc_hd__mux2_1
XFILLER_151_857 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12081_ screen.register.currentYbus\[6\] _05778_ net996 screen.register.currentXbus\[30\]
+ vssd1 vssd1 vccd1 vccd1 _06120_ sky130_fd_sc_hd__a22o_1
XFILLER_123_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold680 datapath.rf.registers\[17\]\[15\] vssd1 vssd1 vccd1 vccd1 net2028 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_127_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold691 datapath.rf.registers\[28\]\[30\] vssd1 vssd1 vccd1 vccd1 net2039 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11032_ net177 net1952 net541 vssd1 vssd1 vccd1 vccd1 _00094_ sky130_fd_sc_hd__mux2_1
XFILLER_2_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11167__S net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07760__A2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12983_ net215 net2534 net478 vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__mux2_1
XFILLER_91_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11934_ net136 _05986_ _05985_ vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06785__A _01610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07233__X _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14653_ clknet_leaf_149_clk _01358_ net1060 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11865_ net137 _05940_ _05939_ vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_28_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13604_ clknet_leaf_17_clk _00414_ net1109 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10816_ datapath.mulitply_result\[12\] net599 net621 vssd1 vssd1 vccd1 vccd1 _05574_
+ sky130_fd_sc_hd__a21o_1
X_11796_ datapath.ru.latched_instruction\[2\] net333 net313 _01443_ vssd1 vssd1 vccd1
+ vccd1 _00662_ sky130_fd_sc_hd__a22o_1
XFILLER_13_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14584_ clknet_leaf_6_clk _01289_ net1067 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13535_ clknet_leaf_13_clk _00345_ net1102 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10747_ _01643_ _01663_ vssd1 vssd1 vccd1 vccd1 _05514_ sky130_fd_sc_hd__or2_1
XFILLER_146_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10678_ _05440_ _05493_ _05495_ vssd1 vssd1 vccd1 vccd1 _05496_ sky130_fd_sc_hd__o21ai_1
X_13466_ clknet_leaf_3_clk _00276_ net1076 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_136_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12417_ _05974_ net158 vssd1 vssd1 vccd1 vccd1 _06356_ sky130_fd_sc_hd__nor2_1
XANTENNA__08225__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13397_ clknet_leaf_18_clk _00207_ net1108 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07579__A2 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12348_ _05656_ _06254_ _06314_ net191 vssd1 vssd1 vccd1 vccd1 _06315_ sky130_fd_sc_hd__o22a_1
XFILLER_114_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12279_ net892 _04495_ vssd1 vssd1 vccd1 vccd1 _06265_ sky130_fd_sc_hd__or2_1
XFILLER_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14018_ clknet_leaf_79_clk _00787_ net1254 vssd1 vssd1 vccd1 vccd1 datapath.PC\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__10335__A1 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11077__S net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06840_ _01463_ net1003 net1019 net1026 datapath.ru.latched_instruction\[24\] vssd1
+ vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_52_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06771_ _01575_ _01607_ vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__nor2_1
XFILLER_49_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10769__X _05534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08510_ datapath.rf.registers\[16\]\[1\] net970 net912 _01636_ net990 vssd1 vssd1
+ vccd1 vccd1 _03346_ sky130_fd_sc_hd__o2111a_1
XFILLER_64_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09490_ net362 _04325_ _04324_ net371 vssd1 vssd1 vccd1 vccd1 _04326_ sky130_fd_sc_hd__a211o_1
XFILLER_82_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14013__RESET_B net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08441_ datapath.rf.registers\[28\]\[2\] net753 net737 datapath.rf.registers\[22\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__a22o_1
XANTENNA__06625__C_N mmio.memload_or_instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08372_ datapath.rf.registers\[24\]\[3\] net769 net753 datapath.rf.registers\[28\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03208_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_156_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07323_ net872 _02154_ _02156_ _02158_ vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__or4_2
XFILLER_20_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout137_A _05934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07254_ datapath.rf.registers\[0\]\[26\] net782 _02085_ _02089_ vssd1 vssd1 vccd1
+ vccd1 _02090_ sky130_fd_sc_hd__o22a_4
XFILLER_149_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08415__A net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08216__B1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07185_ datapath.rf.registers\[25\]\[27\] net841 net792 datapath.rf.registers\[18\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__a22o_1
XANTENNA__08767__A1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_857 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1213_A net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12315__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout401 _06553_ vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__buf_4
Xfanout412 _05730_ vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__clkbuf_8
Xfanout423 net425 vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__buf_4
XFILLER_99_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout434 net435 vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__buf_4
XFILLER_58_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout445 net446 vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_92_Left_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout673_A net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_max_cap1046_X net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout456 _03652_ vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__clkbuf_2
Xfanout467 _01701_ vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__buf_2
X_09826_ net905 _03482_ _04658_ _04660_ _04661_ vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10877__A2 _04057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1001_X net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout478 _06556_ vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__clkbuf_8
XFILLER_101_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_107_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout489 _06552_ vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__buf_4
XANTENNA__07742__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout840_A _01740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09757_ _04005_ _04009_ net341 vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__mux2_1
X_06969_ _01636_ net990 net965 vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout559_X net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06876__Y _01712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout938_A net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08708_ _03205_ _03228_ vssd1 vssd1 vccd1 vccd1 _03544_ sky130_fd_sc_hd__nor2_1
XFILLER_15_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09688_ net648 _04523_ net438 vssd1 vssd1 vccd1 vccd1 _04524_ sky130_fd_sc_hd__a21o_1
XANTENNA__09495__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ _03471_ _03474_ _01957_ vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout726_X net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11650_ keypad.decode.sticky\[1\] keypad.decode.sticky\[2\] net1022 keypad.decode.push
+ vssd1 vssd1 vccd1 vccd1 _05873_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_25_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07988__X _02824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10601_ screen.register.currentYbus\[29\] screen.register.currentYbus\[28\] screen.register.currentYbus\[31\]
+ screen.register.currentYbus\[30\] vssd1 vssd1 vccd1 vccd1 _05422_ sky130_fd_sc_hd__or4_1
X_11581_ screen.counter.ct\[20\] screen.counter.ct\[22\] screen.counter.ct\[21\] vssd1
+ vssd1 vccd1 vccd1 _05805_ sky130_fd_sc_hd__or3b_1
XFILLER_22_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11450__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10532_ _05329_ _05350_ _05361_ vssd1 vssd1 vccd1 vccd1 _05362_ sky130_fd_sc_hd__or3_1
XFILLER_80_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13320_ clknet_leaf_62_clk _00130_ net1234 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10574__B net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13251_ clknet_leaf_138_clk _00061_ net1100 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08207__B1 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10463_ screen.counter.ct\[3\] screen.counter.ct\[2\] vssd1 vssd1 vccd1 vccd1 _05293_
+ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_118_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12202_ screen.counter.currentCt\[4\] _06210_ net603 vssd1 vssd1 vccd1 vccd1 _06212_
+ sky130_fd_sc_hd__o21ai_1
X_13182_ net2162 vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__clkbuf_1
X_10394_ net360 _04498_ _05229_ vssd1 vssd1 vccd1 vccd1 _05230_ sky130_fd_sc_hd__o21ai_1
X_12133_ _06167_ net1012 vssd1 vssd1 vccd1 vccd1 _06170_ sky130_fd_sc_hd__and2b_1
XFILLER_124_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12064_ screen.register.currentYbus\[29\] _05757_ _05837_ screen.register.currentYbus\[21\]
+ vssd1 vssd1 vccd1 vccd1 _06104_ sky130_fd_sc_hd__a22o_1
XFILLER_49_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11015_ net269 datapath.rf.registers\[27\]\[11\] net540 vssd1 vssd1 vccd1 vccd1 _00077_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07194__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07733__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout990 _01646_ vssd1 vssd1 vccd1 vccd1 net990 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06941__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12966_ net298 net2484 net478 vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__mux2_1
XANTENNA__09486__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11917_ net2628 net160 vssd1 vssd1 vccd1 vccd1 _05975_ sky130_fd_sc_hd__nand2_1
X_12897_ net2357 net260 net485 vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__mux2_1
X_14636_ clknet_leaf_17_clk _01341_ net1108 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07123__B _01707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11848_ _05303_ _05795_ _05331_ vssd1 vssd1 vccd1 vccd1 _05927_ sky130_fd_sc_hd__a21oi_1
XFILLER_61_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14567_ clknet_leaf_145_clk _01272_ net1087 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11779_ net123 _05442_ _05894_ vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__mux2_1
XANTENNA__11360__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06962__B _01797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10253__B1 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13518_ clknet_leaf_5_clk _00328_ net1067 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_147_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14498_ clknet_leaf_152_clk _01203_ net1052 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_151_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload11 clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clkload11/Y sky130_fd_sc_hd__inv_6
Xclkload22 clknet_leaf_150_clk vssd1 vssd1 vccd1 vccd1 clkload22/X sky130_fd_sc_hd__clkbuf_4
X_13449_ clknet_leaf_92_clk _00259_ net1234 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_62_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload33 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 clkload33/Y sky130_fd_sc_hd__inv_8
Xclkload44 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 clkload44/Y sky130_fd_sc_hd__inv_8
XFILLER_115_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload55 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 clkload55/Y sky130_fd_sc_hd__clkinv_2
Xclkload66 clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 clkload66/Y sky130_fd_sc_hd__inv_6
XANTENNA__08522__X _03358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload77 clknet_leaf_56_clk vssd1 vssd1 vccd1 vccd1 clkload77/Y sky130_fd_sc_hd__clkinv_2
Xclkload88 clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 clkload88/Y sky130_fd_sc_hd__bufinv_16
XFILLER_126_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload99 clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 clkload99/X sky130_fd_sc_hd__clkbuf_8
XFILLER_5_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08990_ _03823_ _03825_ net600 vssd1 vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_71_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07972__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07941_ datapath.rf.registers\[18\]\[11\] net976 net949 vssd1 vssd1 vccd1 vccd1 _02777_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08401__C net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07872_ datapath.rf.registers\[28\]\[13\] net753 net733 datapath.rf.registers\[19\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__a22o_1
XANTENNA__07185__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07724__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09611_ net464 _03126_ net623 vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__a21oi_1
X_06823_ _01536_ net1016 net993 vssd1 vssd1 vccd1 vccd1 _01659_ sky130_fd_sc_hd__and3_1
X_09542_ _03009_ net560 net441 vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__mux2_1
X_06754_ _01572_ _01591_ vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__or2_1
XFILLER_37_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06685_ net1286 net1285 mmio.memload_or_instruction\[16\] vssd1 vssd1 vccd1 vccd1
+ _01524_ sky130_fd_sc_hd__or3b_1
X_09473_ net349 _04282_ _04277_ net358 vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_102_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_90_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_90_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07033__B net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08424_ _03257_ _03258_ _03259_ vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__or3_1
XFILLER_51_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08844__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08355_ datapath.rf.registers\[16\]\[3\] net862 net830 datapath.rf.registers\[14\]\[3\]
+ _03182_ vssd1 vssd1 vccd1 vccd1 _03191_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_82_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout421_A _05722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11270__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout519_A net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10244__B1 net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07306_ datapath.rf.registers\[24\]\[25\] net768 net673 datapath.rf.registers\[7\]\[25\]
+ _02132_ vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__a221o_1
Xclkload5 clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clkload5/X sky130_fd_sc_hd__clkbuf_8
X_08286_ _03107_ _03108_ _03120_ _03121_ vssd1 vssd1 vccd1 vccd1 _03122_ sky130_fd_sc_hd__or4_1
X_07237_ datapath.rf.registers\[12\]\[26\] net754 net702 datapath.rf.registers\[9\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout307_X net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07168_ _01981_ _02003_ vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout790_A net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout888_A net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07099_ datapath.rf.registers\[0\]\[29\] net871 _01920_ net592 vssd1 vssd1 vccd1
+ vccd1 _01935_ sky130_fd_sc_hd__a2bb2o_4
XANTENNA__07963__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1207 net1213 vssd1 vssd1 vccd1 vccd1 net1207 sky130_fd_sc_hd__clkbuf_4
Xfanout1218 net1219 vssd1 vssd1 vccd1 vccd1 net1218 sky130_fd_sc_hd__clkbuf_4
Xfanout220 net221 vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__clkbuf_2
XFILLER_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1229 net1230 vssd1 vssd1 vccd1 vccd1 net1229 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout676_X net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout231 net234 vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__clkbuf_2
Xfanout242 _05605_ vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout253 _05588_ vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__clkbuf_2
Xfanout264 _05575_ vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_89_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06887__X _01723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout275 net276 vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07715__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout286 _05706_ vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11953__B net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout297 _05536_ vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__clkbuf_2
X_09809_ _01706_ _04629_ _04631_ _04644_ vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__o22ai_4
XFILLER_46_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout843_X net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11445__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12820_ net2115 net203 net490 vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__mux2_1
XFILLER_61_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12751_ net1607 net232 net404 vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_81_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_clk sky130_fd_sc_hd__clkbuf_8
X_11702_ _04909_ net154 net149 net1405 vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__a22o_1
X_12682_ _06514_ _06515_ vssd1 vssd1 vccd1 vccd1 _06516_ sky130_fd_sc_hd__xor2_1
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14421_ clknet_leaf_129_clk _01126_ net1117 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_91_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11633_ _05759_ _05851_ _05854_ _05855_ _05813_ vssd1 vssd1 vccd1 vccd1 _05857_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10585__A _03028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11180__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06782__B _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14352_ clknet_leaf_57_clk _01057_ net1160 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11564_ net1008 _05787_ vssd1 vssd1 vccd1 vccd1 _05788_ sky130_fd_sc_hd__nor2_1
XFILLER_7_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07100__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11983__B1 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13303_ clknet_leaf_124_clk _00113_ net1208 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10515_ net1279 net1274 net1270 screen.counter.ct\[20\] vssd1 vssd1 vccd1 vccd1 _05345_
+ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_133_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11495_ net240 net1662 net512 vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__mux2_1
X_14283_ clknet_leaf_64_clk _00988_ net1236 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_133_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13234_ clknet_leaf_32_clk _00044_ net1126 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10446_ _05271_ _05281_ vssd1 vssd1 vccd1 vccd1 _05282_ sky130_fd_sc_hd__nand2_1
XFILLER_6_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13165_ net2147 vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__clkbuf_1
X_10377_ _03716_ _04706_ vssd1 vssd1 vccd1 vccd1 _05213_ sky130_fd_sc_hd__nor2_1
XANTENNA__08502__B net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07954__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12116_ net1271 net1272 screen.counter.ct\[16\] vssd1 vssd1 vccd1 vccd1 _06153_ sky130_fd_sc_hd__and3_1
X_13096_ net259 net1588 net472 vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__mux2_1
XFILLER_105_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12047_ net1393 _06017_ _06088_ vssd1 vssd1 vccd1 vccd1 _00730_ sky130_fd_sc_hd__a21o_1
XANTENNA__08929__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07167__B1 _01787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07706__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09614__A net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06914__B1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11355__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06957__B net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_148_Left_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13998_ clknet_leaf_113_clk _00775_ net1195 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06676__C datapath.ru.latched_instruction\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07134__A net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12949_ net234 net1702 net396 vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_72_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08131__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06973__A _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14619_ clknet_leaf_38_clk _01324_ net1145 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07890__A1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11090__S net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08140_ _02964_ _02966_ _02973_ _02975_ vssd1 vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__or4_1
XANTENNA__10226__B1 _01702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload100 clknet_leaf_121_clk vssd1 vssd1 vccd1 vccd1 clkload100/Y sky130_fd_sc_hd__bufinv_16
X_08071_ datapath.rf.registers\[8\]\[9\] net878 _02882_ _02885_ _02893_ vssd1 vssd1
+ vccd1 vccd1 _02907_ sky130_fd_sc_hd__a2111o_1
XANTENNA__14117__D datapath.multiplication_module.zero_multi vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xclkload111 clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 clkload111/Y sky130_fd_sc_hd__inv_8
XANTENNA__10782__X _05545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload122 clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 clkload122/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__12914__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload133 clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 clkload133/Y sky130_fd_sc_hd__inv_8
X_07022_ net566 _01856_ vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__and2b_1
Xclkload144 clknet_leaf_80_clk vssd1 vssd1 vccd1 vccd1 clkload144/Y sky130_fd_sc_hd__inv_6
XFILLER_127_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08198__A2 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06748__A3 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08973_ _03204_ net446 _03808_ vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__a21o_1
Xhold17 keypad.debounce.debounce\[14\] vssd1 vssd1 vccd1 vccd1 net1365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 datapath.ru.ack_mul_reg vssd1 vssd1 vccd1 vccd1 net1376 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07924_ datapath.rf.registers\[22\]\[12\] net735 net669 datapath.rf.registers\[21\]\[12\]
+ _02759_ vssd1 vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__a221o_1
XFILLER_152_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold39 screen.controlBus\[30\] vssd1 vssd1 vccd1 vccd1 net1387 sky130_fd_sc_hd__dlygate4sd3_1
X_07855_ datapath.rf.registers\[13\]\[13\] net810 _02689_ _02690_ net873 vssd1 vssd1
+ vccd1 vccd1 _02691_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__10701__A1 _03076_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11265__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout469_A _01701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06806_ _01438_ net1014 vssd1 vssd1 vccd1 vccd1 _01642_ sky130_fd_sc_hd__and2_1
X_07786_ datapath.rf.registers\[20\]\[15\] net718 net699 datapath.rf.registers\[23\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02622_ sky130_fd_sc_hd__a22o_1
XFILLER_84_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09525_ net355 _04213_ _04360_ vssd1 vssd1 vccd1 vccd1 _04361_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_84_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06737_ _01571_ _01574_ vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__nand2_2
Xclkbuf_leaf_63_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_101_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06668_ datapath.ru.latched_instruction\[26\] _01504_ _01506_ datapath.ru.latched_instruction\[21\]
+ vssd1 vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__o22a_1
X_09456_ net376 _04291_ net379 vssd1 vssd1 vccd1 vccd1 _04292_ sky130_fd_sc_hd__a21oi_1
XFILLER_52_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07330__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08407_ datapath.rf.registers\[31\]\[2\] net980 net916 vssd1 vssd1 vccd1 vccd1 _03243_
+ sky130_fd_sc_hd__and3_1
XFILLER_40_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06599_ net1287 net1282 mmio.memload_or_instruction\[7\] vssd1 vssd1 vccd1 vccd1
+ _01438_ sky130_fd_sc_hd__nor3b_2
XANTENNA_fanout424_X net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09387_ _04221_ _04222_ net346 _04220_ vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout803_A _01769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09083__A0 _02025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08338_ _03149_ _03171_ vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__nor2_1
XFILLER_137_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08269_ datapath.rf.registers\[30\]\[5\] net759 net751 datapath.rf.registers\[28\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03105_ sky130_fd_sc_hd__a22o_1
XANTENNA__12824__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10300_ datapath.PC\[5\] _05135_ net1252 vssd1 vssd1 vccd1 vccd1 _05136_ sky130_fd_sc_hd__mux2_1
XFILLER_153_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11280_ net291 net2431 net522 vssd1 vssd1 vccd1 vccd1 _00328_ sky130_fd_sc_hd__mux2_1
XFILLER_146_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout793_X net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08189__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10231_ _03865_ _04625_ _03827_ vssd1 vssd1 vccd1 vccd1 _05067_ sky130_fd_sc_hd__o21ai_1
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10344__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07397__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10571__C _02912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07936__A2 _02771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10162_ net890 _04177_ vssd1 vssd1 vccd1 vccd1 _04998_ sky130_fd_sc_hd__nor2_1
XFILLER_106_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout960_X net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1004 net1005 vssd1 vssd1 vccd1 vccd1 net1004 sky130_fd_sc_hd__buf_4
Xfanout1015 _01562_ vssd1 vssd1 vccd1 vccd1 net1015 sky130_fd_sc_hd__buf_2
XFILLER_86_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1026 net1028 vssd1 vssd1 vccd1 vccd1 net1026 sky130_fd_sc_hd__buf_4
X_10093_ net225 _04923_ _04926_ _04927_ vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__or4_1
Xfanout1048 net1049 vssd1 vssd1 vccd1 vccd1 net1048 sky130_fd_sc_hd__buf_2
XFILLER_48_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07149__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1059 net1061 vssd1 vssd1 vccd1 vccd1 net1059 sky130_fd_sc_hd__clkbuf_4
X_13921_ clknet_leaf_109_clk _00699_ net1220 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09434__A _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12131__Y _06168_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11175__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13852_ clknet_leaf_49_clk _00656_ net1177 vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__dfrtp_1
X_12803_ net1842 net293 net490 vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__mux2_1
XFILLER_74_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13783_ clknet_leaf_52_clk _00592_ net1181 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10995_ net1722 net194 net435 vssd1 vssd1 vccd1 vccd1 _00060_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_54_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09310__A1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12734_ net2044 net304 net405 vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__mux2_1
XANTENNA__07321__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12665_ net498 _06500_ _06501_ net502 net2559 vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__a32o_1
XFILLER_31_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14404_ clknet_leaf_22_clk _01109_ net1156 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11616_ net1007 _05760_ vssd1 vssd1 vccd1 vccd1 _05840_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_13_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09074__B1 _03721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12596_ _06442_ _06443_ vssd1 vssd1 vccd1 vccd1 _06444_ sky130_fd_sc_hd__nand2b_1
X_14335_ clknet_leaf_14_clk _01040_ net1079 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12734__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11547_ _05770_ vssd1 vssd1 vccd1 vccd1 _05771_ sky130_fd_sc_hd__inv_2
XFILLER_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold509 datapath.rf.registers\[27\]\[6\] vssd1 vssd1 vccd1 vccd1 net1857 sky130_fd_sc_hd__dlygate4sd3_1
X_14266_ clknet_leaf_2_clk _00971_ net1078 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11858__B net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11478_ _05700_ net2256 net513 vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__mux2_1
XFILLER_125_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13217_ clknet_leaf_56_clk _00027_ net1159 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10429_ _03770_ _05262_ vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__or2_1
X_14197_ clknet_leaf_66_clk datapath.multiplication_module.multiplicand_i_n\[8\] net1237
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[8\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__07388__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07927__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08585__C1 _03419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13148_ net2301 net231 net383 vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__mux2_1
XANTENNA__08800__X _03636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13079_ net1956 net239 net386 vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__mux2_1
Xhold1209 datapath.rf.registers\[28\]\[9\] vssd1 vssd1 vccd1 vccd1 net2557 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11085__S net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07640_ _02469_ _02471_ _02473_ _02475_ vssd1 vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__or4_1
XFILLER_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07571_ datapath.rf.registers\[10\]\[19\] net881 net838 datapath.rf.registers\[26\]\[19\]
+ _02390_ vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__a221o_1
XFILLER_80_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10777__X _05541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12909__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_45_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08104__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09310_ net632 _04120_ _04122_ _04145_ vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__a22oi_4
XANTENNA__07312__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09241_ net337 _03807_ _04076_ _03673_ vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__o211a_1
XFILLER_22_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08407__B net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09172_ _03796_ _03800_ net450 vssd1 vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__mux2_1
X_08123_ _02951_ _02952_ _02956_ _02958_ vssd1 vssd1 vccd1 vccd1 _02959_ sky130_fd_sc_hd__nor4_1
XFILLER_108_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07030__C _01712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout217_A _05628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09078__X _03914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08054_ datapath.rf.registers\[21\]\[9\] net947 net924 vssd1 vssd1 vccd1 vccd1 _02890_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07091__A2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07005_ datapath.rf.registers\[2\]\[31\] net743 net684 datapath.rf.registers\[27\]\[31\]
+ _01840_ vssd1 vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__a221o_1
XANTENNA__09368__A1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07379__B1 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1126_A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07918__A2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08040__B2 datapath.rf.registers\[0\]\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08591__A2 _03423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08956_ _03789_ _03791_ net450 vssd1 vssd1 vccd1 vccd1 _03792_ sky130_fd_sc_hd__mux2_1
XFILLER_130_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07907_ datapath.rf.registers\[10\]\[12\] net879 net848 datapath.rf.registers\[1\]\[12\]
+ _02742_ vssd1 vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout753_A _01804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08887_ _01857_ net623 _03719_ net642 vssd1 vssd1 vccd1 vccd1 _03723_ sky130_fd_sc_hd__o211a_1
XANTENNA__09540__A1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07838_ datapath.rf.registers\[1\]\[14\] net763 net715 datapath.rf.registers\[4\]\[14\]
+ _02662_ vssd1 vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__a221o_1
XFILLER_84_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout920_A _01744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12819__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07769_ datapath.rf.registers\[16\]\[15\] net861 net855 datapath.rf.registers\[19\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout541_X net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout639_X net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_36_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_8
X_09508_ net458 _04340_ _04343_ vssd1 vssd1 vccd1 vccd1 _04344_ sky130_fd_sc_hd__a21o_1
X_10780_ net1268 _05530_ datapath.PC\[7\] vssd1 vssd1 vccd1 vccd1 _05543_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07303__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09439_ net633 _04274_ vssd1 vssd1 vccd1 vccd1 _04275_ sky130_fd_sc_hd__and2_1
XFILLER_13_858 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout806_X net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12450_ net165 _05948_ net127 net2600 vssd1 vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_10_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11401_ net1625 net202 net410 vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__mux2_1
XFILLER_138_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12381_ _05938_ net159 vssd1 vssd1 vccd1 vccd1 _06338_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_97_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14120_ clknet_leaf_78_clk net1376 net1245 vssd1 vssd1 vccd1 vccd1 datapath.ru.ack_mul_reg2
+ sky130_fd_sc_hd__dfrtp_1
X_11332_ net1803 net204 net414 vssd1 vssd1 vccd1 vccd1 _00377_ sky130_fd_sc_hd__mux2_1
XANTENNA__09429__A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07082__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14051_ clknet_leaf_101_clk _00818_ net1228 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11263_ net212 net2177 net418 vssd1 vssd1 vccd1 vccd1 _00312_ sky130_fd_sc_hd__mux2_1
XFILLER_106_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08052__B net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07909__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13002_ net1711 net283 net392 vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__mux2_1
X_10214_ datapath.PC\[18\] net1256 _05047_ _05049_ vssd1 vssd1 vccd1 vccd1 _05050_
+ sky130_fd_sc_hd__o22a_1
XFILLER_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11194_ net233 net2111 net422 vssd1 vssd1 vccd1 vccd1 _00246_ sky130_fd_sc_hd__mux2_1
X_10145_ _04978_ _04979_ _04980_ net1044 net638 vssd1 vssd1 vccd1 vccd1 _04981_ sky130_fd_sc_hd__a221oi_1
XANTENNA__08582__A2 _03417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10802__S net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06788__A _01579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07790__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10076_ datapath.PC\[30\] net468 net1038 vssd1 vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__o21a_1
XFILLER_153_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09531__A1 _03263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13904_ clknet_leaf_43_clk net1367 net1149 vssd1 vssd1 vccd1 vccd1 keypad.debounce.debounce\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_36_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07542__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12796__Y _06551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13835_ clknet_leaf_141_clk _00644_ net1187 vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_141_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_27_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_90_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13766_ clknet_leaf_82_clk _00575_ net1256 vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09295__B1 _02522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10978_ net1654 net276 net436 vssd1 vssd1 vccd1 vccd1 _00043_ sky130_fd_sc_hd__mux2_1
XFILLER_16_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12717_ _05893_ _06539_ _06540_ _06530_ vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__a31o_1
XFILLER_15_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10249__S net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13697_ clknet_leaf_45_clk _00507_ net1147 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_44_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12648_ datapath.mulitply_result\[23\] datapath.multiplication_module.multiplicand_i\[23\]
+ vssd1 vssd1 vccd1 vccd1 _06487_ sky130_fd_sc_hd__nor2_1
XFILLER_12_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12579_ net500 _06428_ _06429_ net504 net1802 vssd1 vssd1 vccd1 vccd1 _00921_ sky130_fd_sc_hd__a32o_1
XANTENNA__06970__B net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14318_ clknet_leaf_0_clk _01023_ net1055 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07073__A2 _01908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold306 datapath.rf.registers\[7\]\[9\] vssd1 vssd1 vccd1 vccd1 net1654 sky130_fd_sc_hd__dlygate4sd3_1
Xhold317 datapath.rf.registers\[7\]\[10\] vssd1 vssd1 vccd1 vccd1 net1665 sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 datapath.rf.registers\[14\]\[0\] vssd1 vssd1 vccd1 vccd1 net1676 sky130_fd_sc_hd__dlygate4sd3_1
Xhold339 datapath.rf.registers\[12\]\[28\] vssd1 vssd1 vccd1 vccd1 net1687 sky130_fd_sc_hd__dlygate4sd3_1
X_14249_ clknet_leaf_20_clk _00954_ net1165 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout808 net809 vssd1 vssd1 vccd1 vccd1 net808 sky130_fd_sc_hd__clkbuf_4
XFILLER_124_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout819 net820 vssd1 vssd1 vccd1 vccd1 net819 sky130_fd_sc_hd__buf_4
XANTENNA__09770__A1 _03947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08810_ _03228_ _03644_ _03645_ vssd1 vssd1 vccd1 vccd1 _03646_ sky130_fd_sc_hd__o21a_1
XANTENNA__10712__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09790_ _03822_ _03826_ _03865_ _04625_ vssd1 vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__a211o_1
XANTENNA__07781__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1006 datapath.rf.registers\[19\]\[28\] vssd1 vssd1 vccd1 vccd1 net2354 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10380__A2 _03418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1017 datapath.rf.registers\[25\]\[18\] vssd1 vssd1 vccd1 vccd1 net2365 sky130_fd_sc_hd__dlygate4sd3_1
X_08741_ _03518_ _03521_ _03576_ vssd1 vssd1 vccd1 vccd1 _03577_ sky130_fd_sc_hd__and3_1
Xhold1028 datapath.rf.registers\[13\]\[7\] vssd1 vssd1 vccd1 vccd1 net2376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1039 datapath.rf.registers\[30\]\[10\] vssd1 vssd1 vccd1 vccd1 net2387 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08325__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08672_ _02419_ _02440_ vssd1 vssd1 vccd1 vccd1 _03508_ sky130_fd_sc_hd__nand2_1
XANTENNA__10132__A2 _04023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07533__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07623_ datapath.rf.registers\[20\]\[18\] net839 net824 datapath.rf.registers\[6\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__a22o_1
XFILLER_54_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07025__C net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_18_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout167_A _05288_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07554_ datapath.rf.registers\[2\]\[19\] net985 net949 vssd1 vssd1 vccd1 vccd1 _02390_
+ sky130_fd_sc_hd__and3_1
X_07485_ datapath.rf.registers\[29\]\[21\] net675 _02319_ _02320_ net786 vssd1 vssd1
+ vccd1 vccd1 _02321_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout1076_A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09224_ _03583_ _04059_ net578 vssd1 vssd1 vccd1 vccd1 _04060_ sky130_fd_sc_hd__o21ai_1
X_09155_ net360 net351 net458 _03772_ vssd1 vssd1 vccd1 vccd1 _03991_ sky130_fd_sc_hd__or4_1
XANTENNA__12374__S net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1243_A net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_885 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06880__B net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08106_ datapath.rf.registers\[8\]\[8\] net956 _01712_ vssd1 vssd1 vccd1 vccd1 _02942_
+ sky130_fd_sc_hd__and3_1
XFILLER_108_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07064__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09086_ net372 _03921_ vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__nand2_1
X_08037_ datapath.rf.registers\[2\]\[10\] net744 net666 datapath.rf.registers\[15\]\[10\]
+ _02859_ vssd1 vssd1 vccd1 vccd1 _02873_ sky130_fd_sc_hd__a221o_1
XFILLER_123_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold840 datapath.rf.registers\[21\]\[8\] vssd1 vssd1 vccd1 vccd1 net2188 sky130_fd_sc_hd__dlygate4sd3_1
Xhold851 mmio.memload_or_instruction\[20\] vssd1 vssd1 vccd1 vccd1 net2199 sky130_fd_sc_hd__dlygate4sd3_1
Xhold862 datapath.rf.registers\[16\]\[24\] vssd1 vssd1 vccd1 vccd1 net2210 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold873 datapath.rf.registers\[21\]\[31\] vssd1 vssd1 vccd1 vccd1 net2221 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold884 datapath.rf.registers\[19\]\[22\] vssd1 vssd1 vccd1 vccd1 net2232 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap592 net593 vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__clkbuf_1
XANTENNA_fanout491_X net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout870_A net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold895 datapath.rf.registers\[13\]\[19\] vssd1 vssd1 vccd1 vccd1 net2243 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08564__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout968_A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09988_ datapath.PC\[27\] net594 vssd1 vssd1 vccd1 vccd1 _04824_ sky130_fd_sc_hd__xnor2_1
XFILLER_130_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07772__B1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08939_ net352 _03774_ vssd1 vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_150_Right_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout756_X net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11950_ net2490 net160 vssd1 vssd1 vccd1 vccd1 _05997_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_4_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07524__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10901_ net201 net2035 net542 vssd1 vssd1 vccd1 vccd1 _00026_ sky130_fd_sc_hd__mux2_1
XANTENNA__11871__A2 _05944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11881_ net2487 net163 vssd1 vssd1 vccd1 vccd1 _05951_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout923_X net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11453__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13620_ clknet_leaf_93_clk _00430_ net1211 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10832_ _01513_ net619 _05586_ _05587_ vssd1 vssd1 vccd1 vccd1 _05588_ sky130_fd_sc_hd__o2bb2a_4
XANTENNA__10577__B _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13551_ clknet_leaf_30_clk _00361_ net1131 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10763_ _01450_ net654 _05527_ _05528_ vssd1 vssd1 vccd1 vccd1 _05529_ sky130_fd_sc_hd__o22a_1
XANTENNA__08047__B net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12502_ net201 net2034 net509 vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__mux2_1
XFILLER_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10831__B1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13482_ clknet_leaf_59_clk _00292_ net1170 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10694_ _05507_ _05509_ vssd1 vssd1 vccd1 vccd1 keypad.decode.button_n\[4\] sky130_fd_sc_hd__nor2_1
XFILLER_139_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12433_ _05990_ net158 vssd1 vssd1 vccd1 vccd1 _06364_ sky130_fd_sc_hd__nor2_1
XFILLER_154_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07055__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12364_ net637 _04902_ vssd1 vssd1 vccd1 vccd1 _06327_ sky130_fd_sc_hd__nor2_1
X_14103_ clknet_leaf_110_clk _00869_ net1202 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_11315_ net2098 net292 net414 vssd1 vssd1 vccd1 vccd1 _00360_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_112_Left_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12295_ _04854_ _05567_ net227 vssd1 vssd1 vccd1 vccd1 _06277_ sky130_fd_sc_hd__mux2_1
XFILLER_107_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14034_ clknet_leaf_84_clk _00803_ net1260 vssd1 vssd1 vccd1 vccd1 datapath.PC\[24\]
+ sky130_fd_sc_hd__dfstp_1
X_11246_ net295 net1820 net419 vssd1 vssd1 vccd1 vccd1 _00295_ sky130_fd_sc_hd__mux2_1
XFILLER_79_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11177_ net304 net1613 net424 vssd1 vssd1 vccd1 vccd1 _00229_ sky130_fd_sc_hd__mux2_1
XFILLER_94_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10128_ datapath.PC\[21\] net1295 _04961_ _04963_ vssd1 vssd1 vccd1 vccd1 _04964_
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__08307__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09504__A1 _02960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10059_ datapath.PC\[29\] net595 vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_121_Left_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10768__A net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11363__S net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06965__B _01800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13818_ clknet_leaf_115_clk _00627_ net1189 vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__dfrtp_1
XFILLER_149_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13749_ clknet_leaf_88_clk _00558_ net1252 vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__dfrtp_1
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07270_ datapath.rf.registers\[11\]\[25\] net986 net938 vssd1 vssd1 vccd1 vccd1 _02106_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07294__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06981__A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_130_Left_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07046__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold103 datapath.multiplication_module.multiplier_i\[12\] vssd1 vssd1 vccd1 vccd1
+ net1451 sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 mmio.memload_or_instruction\[25\] vssd1 vssd1 vccd1 vccd1 net1462 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08404__C net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold125 datapath.multiplication_module.multiplier_i\[11\] vssd1 vssd1 vccd1 vccd1
+ net1473 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10790__X _05552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold136 keypad.decode.sticky_n\[1\] vssd1 vssd1 vccd1 vccd1 net1484 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12922__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_7_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_8
Xhold147 net75 vssd1 vssd1 vccd1 vccd1 net1495 sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 keypad.decode.push vssd1 vssd1 vccd1 vccd1 net1506 sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ _01618_ _03670_ vssd1 vssd1 vccd1 vccd1 _04747_ sky130_fd_sc_hd__and2b_1
Xhold169 datapath.multiplication_module.multiplicand_i\[25\] vssd1 vssd1 vccd1 vccd1
+ net1517 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08701__A _02912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout605 net606 vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09743__A1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout616 _01623_ vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__clkbuf_4
X_09842_ net558 _03419_ vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__nor2_1
Xfanout627 net629 vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__clkbuf_4
Xfanout638 net639 vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout649 net650 vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__clkbuf_4
XFILLER_113_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09773_ _01706_ _04608_ vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__nor2_1
X_06985_ net964 _01820_ vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__and2_1
XFILLER_67_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08724_ _03057_ _03079_ vssd1 vssd1 vccd1 vccd1 _03560_ sky130_fd_sc_hd__nand2_1
XANTENNA__07036__B net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_7_0_clk_X clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_831 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08655_ _02070_ _02091_ vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_1_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06875__B _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07606_ _02418_ _02440_ vssd1 vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_105_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08586_ _03360_ _03421_ vssd1 vssd1 vccd1 vccd1 _03422_ sky130_fd_sc_hd__nand2_1
XFILLER_35_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08148__A _02960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07537_ datapath.rf.registers\[20\]\[20\] net718 net698 datapath.rf.registers\[23\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout716_A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07285__A2 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07468_ datapath.rf.registers\[22\]\[21\] net821 net813 datapath.rf.registers\[23\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__a22o_1
XFILLER_139_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09207_ net356 _04041_ _04042_ _04036_ vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout504_X net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07399_ datapath.rf.registers\[3\]\[23\] net770 net762 datapath.rf.registers\[1\]\[23\]
+ _02234_ vssd1 vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__a221o_1
XFILLER_6_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09138_ net320 _03714_ vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_20_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09069_ _03709_ _03711_ net448 vssd1 vssd1 vccd1 vccd1 _03905_ sky130_fd_sc_hd__mux2_1
XANTENNA__12832__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11100_ net185 net1761 net534 vssd1 vssd1 vccd1 vccd1 _00157_ sky130_fd_sc_hd__mux2_1
XFILLER_78_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11956__B _05786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12080_ _06119_ net1442 _06017_ vssd1 vssd1 vccd1 vccd1 _00732_ sky130_fd_sc_hd__mux2_1
XFILLER_151_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout873_X net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold670 datapath.rf.registers\[10\]\[0\] vssd1 vssd1 vccd1 vccd1 net2018 sky130_fd_sc_hd__dlygate4sd3_1
Xhold681 datapath.rf.registers\[2\]\[18\] vssd1 vssd1 vccd1 vccd1 net2029 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11448__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08537__A2 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold692 datapath.rf.registers\[17\]\[11\] vssd1 vssd1 vccd1 vccd1 net2040 sky130_fd_sc_hd__dlygate4sd3_1
X_11031_ net187 net2413 net539 vssd1 vssd1 vccd1 vccd1 _00093_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07745__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12097__A2 _06018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12982_ net234 net1635 net480 vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__mux2_1
XANTENNA__09498__B1 _04328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input12_A DAT_I[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09442__A _02750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11933_ _02145_ net658 vssd1 vssd1 vccd1 vccd1 _05986_ sky130_fd_sc_hd__nand2_1
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06785__B net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11183__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14652_ clknet_leaf_8_clk _01357_ net1072 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11864_ _03292_ net658 vssd1 vssd1 vccd1 vccd1 _05940_ sky130_fd_sc_hd__nand2_1
XFILLER_72_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13603_ clknet_leaf_119_clk _00413_ net1191 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10815_ _04580_ _05572_ net899 vssd1 vssd1 vccd1 vccd1 _05573_ sky130_fd_sc_hd__mux2_1
X_14583_ clknet_leaf_133_clk _01288_ net1111 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11795_ datapath.ru.latched_instruction\[1\] net336 net316 _01502_ vssd1 vssd1 vccd1
+ vccd1 _00661_ sky130_fd_sc_hd__a22o_1
X_13534_ clknet_leaf_147_clk _00344_ net1062 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07276__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10746_ _01648_ _03264_ vssd1 vssd1 vccd1 vccd1 _05513_ sky130_fd_sc_hd__nand2_1
XANTENNA__10594__Y datapath.multiplication_module.zero_multi vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13465_ clknet_leaf_29_clk _00275_ net1131 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10677_ _05428_ _05443_ _05494_ _05490_ _05459_ vssd1 vssd1 vccd1 vccd1 _05495_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_136_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12416_ net1398 net131 _06355_ vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__a21o_1
XANTENNA__07028__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13396_ clknet_leaf_128_clk _00206_ net1210 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12742__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12347_ net637 _04888_ vssd1 vssd1 vccd1 vccd1 _06314_ sky130_fd_sc_hd__nor2_1
XANTENNA__07984__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12278_ net1268 net309 _06262_ _06264_ vssd1 vssd1 vccd1 vccd1 _00785_ sky130_fd_sc_hd__a22o_1
XANTENNA__11358__S net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09186__C1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14017_ clknet_leaf_86_clk _00786_ net1254 vssd1 vssd1 vccd1 vccd1 datapath.PC\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08528__A2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11229_ net216 net2000 net526 vssd1 vssd1 vccd1 vccd1 _00279_ sky130_fd_sc_hd__mux2_1
XFILLER_96_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07736__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07200__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11882__A _02980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09489__A0 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06770_ _01571_ _01579_ _01588_ vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__or3_4
XANTENNA__06976__A net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11093__S net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08161__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08440_ datapath.rf.registers\[2\]\[2\] net745 net682 datapath.rf.registers\[6\]\[2\]
+ _03274_ vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__a221o_1
X_08371_ _03206_ vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__inv_2
XANTENNA__12917__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07322_ datapath.rf.registers\[2\]\[24\] net887 net807 datapath.rf.registers\[27\]\[24\]
+ _02157_ vssd1 vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__a221o_1
X_07253_ _02076_ _02081_ _02087_ _02088_ vssd1 vssd1 vccd1 vccd1 _02089_ sky130_fd_sc_hd__or4_1
XFILLER_118_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07184_ datapath.rf.registers\[11\]\[27\] net883 net850 datapath.rf.registers\[17\]\[27\]
+ _02007_ vssd1 vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__a221o_1
XANTENNA__08767__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07975__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1039_A net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout499_A net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11268__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout402 _06549_ vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08519__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout413 _05730_ vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout424 net425 vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1206_A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout435 net437 vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08150__B net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout446 net447 vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__buf_2
XANTENNA_input4_A DAT_I[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout457 net458 vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__buf_2
X_09825_ _04652_ _04653_ _03700_ _04237_ vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__a2bb2o_1
Xfanout468 net469 vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__clkbuf_4
XFILLER_58_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout479 _06556_ vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout666_A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09756_ net575 _04590_ _04591_ _04589_ vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__a22o_1
XFILLER_104_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06886__A net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06968_ net964 net911 _01795_ vssd1 vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__and3_4
X_08707_ net463 _03172_ vssd1 vssd1 vccd1 vccd1 _03543_ sky130_fd_sc_hd__nor2_1
X_09687_ _03889_ _04522_ net326 vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout833_A net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06899_ net976 _01707_ net947 vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_87_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07053__Y _01889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08638_ _03470_ _03472_ _02004_ vssd1 vssd1 vccd1 vccd1 _03474_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_120_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11039__A0 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12827__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08569_ datapath.rf.registers\[9\]\[0\] net704 _03402_ _03403_ _03404_ vssd1 vssd1
+ vccd1 vccd1 _03405_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_25_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout719_X net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10600_ _05417_ _05418_ _05420_ vssd1 vssd1 vccd1 vccd1 _05421_ sky130_fd_sc_hd__or3_1
XFILLER_23_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11580_ net1277 screen.counter.ct\[11\] net1275 net1276 vssd1 vssd1 vccd1 vccd1 _05804_
+ sky130_fd_sc_hd__or4b_1
XANTENNA__08606__A _02750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09652__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10531_ net1273 net1272 screen.counter.ct\[18\] screen.counter.ct\[21\] vssd1 vssd1
+ vccd1 vccd1 _05361_ sky130_fd_sc_hd__and4_1
XFILLER_7_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10574__C net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13250_ clknet_leaf_0_clk _00060_ net1054 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10462_ screen.counter.ct\[1\] screen.counter.ct\[0\] vssd1 vssd1 vccd1 vccd1 _05292_
+ sky130_fd_sc_hd__nand2_2
XANTENNA__12003__A2 _05773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout990_X net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12201_ _06210_ _06211_ vssd1 vssd1 vccd1 vccd1 _00761_ sky130_fd_sc_hd__nor2_1
X_13181_ net2010 vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_135_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10393_ net351 _04418_ _05227_ _05228_ net358 vssd1 vssd1 vccd1 vccd1 _05229_ sky130_fd_sc_hd__a221o_1
XFILLER_108_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11762__B2 _02283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12132_ screen.counter.currentEnable _06167_ vssd1 vssd1 vccd1 vccd1 _06169_ sky130_fd_sc_hd__or2_1
XANTENNA__07430__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_131_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11178__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12063_ _06103_ net1460 _06017_ vssd1 vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__mux2_1
XANTENNA__07718__B1 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08060__B net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11973__Y _06018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11014_ net273 net2400 net540 vssd1 vssd1 vccd1 vccd1 _00076_ sky130_fd_sc_hd__mux2_1
XFILLER_93_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout980 _01651_ vssd1 vssd1 vccd1 vccd1 net980 sky130_fd_sc_hd__clkbuf_2
Xfanout991 net992 vssd1 vssd1 vccd1 vccd1 net991 sky130_fd_sc_hd__clkbuf_4
XFILLER_38_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12965_ net303 net1861 net481 vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__mux2_1
XANTENNA__09340__C1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11916_ net136 _05974_ _05973_ vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__o21ai_1
X_12896_ net2204 net209 net485 vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__mux2_1
XFILLER_61_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14635_ clknet_leaf_54_clk _01340_ net1179 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11847_ _05849_ _05925_ vssd1 vssd1 vccd1 vccd1 _05926_ sky130_fd_sc_hd__nor2_1
XANTENNA__07123__C net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12737__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07249__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14566_ clknet_leaf_23_clk _01271_ net1154 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11778_ net122 _05451_ _05894_ vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__mux2_1
XANTENNA__09643__B1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08075__X _02911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13517_ clknet_leaf_125_clk _00327_ net1207 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10729_ net2411 _02612_ net573 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[15\]
+ sky130_fd_sc_hd__mux2_1
X_14497_ clknet_leaf_45_clk _01202_ net1147 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_151_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13448_ clknet_leaf_65_clk _00258_ net1238 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload12 clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clkload12/Y sky130_fd_sc_hd__inv_12
Xclkload23 clknet_leaf_151_clk vssd1 vssd1 vccd1 vccd1 clkload23/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_58_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload34 clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 clkload34/Y sky130_fd_sc_hd__inv_6
Xclkload45 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 clkload45/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload56 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 clkload56/Y sky130_fd_sc_hd__inv_6
X_13379_ clknet_leaf_120_clk _00189_ net1193 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload67 clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 clkload67/Y sky130_fd_sc_hd__inv_6
XFILLER_55_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload78 clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 clkload78/Y sky130_fd_sc_hd__inv_6
Xclkload89 clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 clkload89/Y sky130_fd_sc_hd__inv_6
XANTENNA__11753__B2 _02725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_53_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09347__A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07421__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11088__S net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07940_ datapath.rf.registers\[8\]\[11\] net955 _01712_ vssd1 vssd1 vccd1 vccd1 _02776_
+ sky130_fd_sc_hd__and3_1
X_07871_ datapath.rf.registers\[16\]\[13\] net739 net707 datapath.rf.registers\[10\]\[13\]
+ _02706_ vssd1 vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__a221o_1
XFILLER_29_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08382__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09610_ _03667_ _04437_ _04438_ _04445_ vssd1 vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__o22ai_2
XANTENNA__09614__D_N _04446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_68_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06822_ _01655_ _01657_ datapath.ru.latched_instruction\[16\] vssd1 vssd1 vccd1 vccd1
+ _01658_ sky130_fd_sc_hd__mux2_1
XFILLER_84_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_111_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09541_ _02913_ _02961_ net441 vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__mux2_1
X_06753_ _01574_ _01579_ _01588_ vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__or3_1
XANTENNA__11808__A2 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07488__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07314__B net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09472_ _04305_ _04306_ net460 vssd1 vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_69_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06684_ mmio.memload_or_instruction\[16\] net1048 vssd1 vssd1 vccd1 vccd1 _01523_
+ sky130_fd_sc_hd__and2_1
XFILLER_91_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_102_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08423_ datapath.rf.registers\[12\]\[2\] net828 _03232_ _03234_ _03235_ vssd1 vssd1
+ vccd1 vccd1 _03259_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07033__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_126_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout247_A net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08354_ datapath.rf.registers\[13\]\[3\] net989 net918 vssd1 vssd1 vccd1 vccd1 _03190_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_82_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07305_ datapath.rf.registers\[14\]\[25\] net776 net681 datapath.rf.registers\[6\]\[25\]
+ _02140_ vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__a221o_1
XFILLER_138_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload6 clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clkload6/Y sky130_fd_sc_hd__clkinvlp_4
X_08285_ datapath.rf.registers\[24\]\[5\] net767 net672 datapath.rf.registers\[7\]\[5\]
+ _03109_ vssd1 vssd1 vccd1 vccd1 _03121_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout414_A _05726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1156_A net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08145__B _01784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07236_ datapath.rf.registers\[20\]\[26\] net718 net660 datapath.rf.registers\[5\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02072_ sky130_fd_sc_hd__a22o_1
XFILLER_145_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07167_ net610 _02001_ _01787_ vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__o21ai_2
XFILLER_3_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11744__B2 _03170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07098_ _01920_ net593 datapath.rf.registers\[0\]\[29\] net871 vssd1 vssd1 vccd1
+ vccd1 _01934_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_106_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout783_A net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout210 net211 vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__clkbuf_2
Xfanout1208 net1213 vssd1 vssd1 vccd1 vccd1 net1208 sky130_fd_sc_hd__buf_2
Xfanout1219 net1222 vssd1 vssd1 vccd1 vccd1 net1219 sky130_fd_sc_hd__buf_2
Xfanout221 _05610_ vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__clkbuf_2
Xfanout232 net234 vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__clkbuf_2
Xfanout243 net246 vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__clkbuf_2
Xfanout254 net257 vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__clkbuf_2
Xfanout265 _05575_ vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_89_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout669_X net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08373__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout276 net277 vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__clkbuf_2
Xfanout287 _05706_ vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__buf_1
X_09808_ _04643_ vssd1 vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__inv_2
XFILLER_86_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout298 net299 vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__clkbuf_2
XFILLER_75_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09739_ _04571_ _04574_ _03667_ _04570_ vssd1 vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08100__S net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout836_X net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12750_ net2378 net238 net404 vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__mux2_1
XANTENNA__07479__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11701_ _04919_ net154 net149 net1403 vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__a22o_1
XFILLER_70_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12681_ _06507_ _06509_ _06508_ vssd1 vssd1 vccd1 vccd1 _06515_ sky130_fd_sc_hd__o21ba_1
XANTENNA__11461__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14420_ clknet_leaf_93_clk _01125_ net1212 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11632_ _05855_ vssd1 vssd1 vccd1 vccd1 _05856_ sky130_fd_sc_hd__inv_2
XANTENNA__09625__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10585__B _03076_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10235__A1 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14351_ clknet_leaf_26_clk _01056_ net1137 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11563_ _05763_ _05774_ vssd1 vssd1 vccd1 vccd1 _05787_ sky130_fd_sc_hd__or2_1
XFILLER_11_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08055__B net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13302_ clknet_leaf_141_clk _00112_ net1095 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10514_ _05343_ vssd1 vssd1 vccd1 vccd1 _05344_ sky130_fd_sc_hd__inv_2
X_14282_ clknet_leaf_91_clk _00987_ net1241 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_137_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07651__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11494_ net243 net2384 net510 vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_133_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13233_ clknet_leaf_40_clk _00043_ net1140 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07894__B net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10445_ _05278_ _05280_ datapath.PC\[3\] net1292 vssd1 vssd1 vccd1 vccd1 _05281_
+ sky130_fd_sc_hd__a2bb2o_2
XANTENNA__10805__S net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13164_ net2267 vssd1 vssd1 vccd1 vccd1 _00986_ sky130_fd_sc_hd__clkbuf_1
XFILLER_156_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10376_ net466 net1039 net634 vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__a21o_1
XANTENNA__10943__C1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12115_ _06145_ _06146_ _06151_ vssd1 vssd1 vccd1 vccd1 _06152_ sky130_fd_sc_hd__nor3_1
XANTENNA__08502__C _01797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13095_ net208 net1577 net472 vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_15_0_clk_X clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12046_ _06017_ _06072_ _06087_ vssd1 vssd1 vccd1 vccd1 _06088_ sky130_fd_sc_hd__and3b_1
XANTENNA__07167__A1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08364__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10171__B1 _05002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13997_ clknet_leaf_113_clk _00774_ net1197 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_81_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08116__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13948__SET_B net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12948_ net235 net1877 net396 vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__mux2_1
XFILLER_33_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11671__B1 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12879_ net245 net2063 net398 vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__mux2_1
XANTENNA__11371__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06973__B _01647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14618_ clknet_leaf_14_clk _01323_ net1078 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07890__A2 _02725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14549_ clknet_leaf_130_clk _01254_ net1111 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10777__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08070_ _02902_ _02903_ _02904_ _02905_ vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__or4_1
XANTENNA__07642__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload101 clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 clkload101/Y sky130_fd_sc_hd__inv_6
Xclkload112 clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 clkload112/Y sky130_fd_sc_hd__clkinv_2
Xclkload123 clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 clkload123/Y sky130_fd_sc_hd__inv_8
Xclkload134 clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 clkload134/Y sky130_fd_sc_hd__clkinvlp_4
X_07021_ _01856_ net566 vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__and2b_1
Xclkload145 clknet_leaf_81_clk vssd1 vssd1 vccd1 vccd1 clkload145/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__06850__B1 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10934__C1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08972_ net463 net446 vssd1 vssd1 vccd1 vccd1 _03808_ sky130_fd_sc_hd__nor2_1
XANTENNA__12930__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06988__X _01824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07923_ datapath.rf.registers\[19\]\[12\] net733 _02758_ net786 vssd1 vssd1 vccd1
+ vccd1 _02759_ sky130_fd_sc_hd__a211o_1
Xhold18 keypad.debounce.debounce\[12\] vssd1 vssd1 vccd1 vccd1 net1366 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 mmio.memload_or_instruction\[6\] vssd1 vssd1 vccd1 vccd1 net1377 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08355__B1 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07854_ datapath.rf.registers\[24\]\[13\] net857 net807 datapath.rf.registers\[27\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__a22o_1
X_06805_ _01640_ vssd1 vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__inv_2
XFILLER_84_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07785_ datapath.rf.registers\[4\]\[15\] net715 net692 datapath.rf.registers\[13\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02621_ sky130_fd_sc_hd__a22o_1
XANTENNA__08107__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09304__C1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09524_ net461 _03929_ _03997_ net352 vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_84_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06736_ datapath.ru.latched_instruction\[5\] net1030 net994 _01441_ vssd1 vssd1 vccd1
+ vccd1 _01575_ sky130_fd_sc_hd__a22oi_4
X_09455_ net370 _04290_ _04288_ vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__o21ai_1
X_06667_ net1286 net1285 mmio.memload_or_instruction\[21\] vssd1 vssd1 vccd1 vccd1
+ _01506_ sky130_fd_sc_hd__or3b_1
XANTENNA_fanout531_A net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08427__Y _03263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11281__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06883__B net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08406_ datapath.rf.registers\[14\]\[2\] net988 _01745_ vssd1 vssd1 vccd1 vccd1 _03242_
+ sky130_fd_sc_hd__and3_1
XFILLER_24_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09386_ net357 _04218_ _04219_ net326 vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__o31ai_1
X_06598_ net1286 net1281 vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__nor2_1
XANTENNA__07881__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08337_ net463 _03171_ vssd1 vssd1 vccd1 vccd1 _03173_ sky130_fd_sc_hd__and2_1
XANTENNA__09083__A1 _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout417_X net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07094__B1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07633__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08268_ _03082_ _03103_ vssd1 vssd1 vccd1 vccd1 _03104_ sky130_fd_sc_hd__nand2_2
XANTENNA__06841__A0 datapath.ru.latched_instruction\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07219_ datapath.rf.registers\[11\]\[26\] net882 net807 datapath.rf.registers\[27\]\[26\]
+ _02054_ vssd1 vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__a221o_1
X_08199_ datapath.rf.registers\[19\]\[6\] net974 net927 vssd1 vssd1 vccd1 vccd1 _03035_
+ sky130_fd_sc_hd__and3_1
XFILLER_152_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13001__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10230_ _05062_ _05063_ _05065_ net638 vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__a211oi_1
XFILLER_3_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout786_X net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10571__D _02960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10161_ datapath.PC\[20\] _04996_ net1256 vssd1 vssd1 vccd1 vccd1 _04997_ sky130_fd_sc_hd__mux2_1
XANTENNA__12840__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1005 _01564_ vssd1 vssd1 vccd1 vccd1 net1005 sky130_fd_sc_hd__buf_2
XFILLER_121_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1016 net1017 vssd1 vssd1 vccd1 vccd1 net1016 sky130_fd_sc_hd__buf_4
Xfanout1027 net1028 vssd1 vssd1 vccd1 vccd1 net1027 sky130_fd_sc_hd__clkbuf_2
X_10092_ net637 _03868_ _03914_ vssd1 vssd1 vccd1 vccd1 _04928_ sky130_fd_sc_hd__and3_1
XFILLER_86_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout953_X net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1038 net1039 vssd1 vssd1 vccd1 vccd1 net1038 sky130_fd_sc_hd__buf_2
XFILLER_59_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1049 net1051 vssd1 vssd1 vccd1 vccd1 net1049 sky130_fd_sc_hd__buf_2
XANTENNA__11456__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13920_ clknet_leaf_109_clk _00698_ net1218 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_142_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13851_ clknet_leaf_49_clk _00655_ net1177 vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__dfrtp_1
XFILLER_142_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12802_ datapath.rf.registers\[1\]\[5\] net296 net490 vssd1 vssd1 vccd1 vccd1 _01054_
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13782_ clknet_leaf_51_clk _00591_ net1181 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10994_ net1632 net197 net436 vssd1 vssd1 vccd1 vccd1 _00059_ sky130_fd_sc_hd__mux2_1
X_12733_ net1660 net288 net405 vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__mux2_1
XANTENNA__11191__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12664_ _06498_ _06499_ _06497_ vssd1 vssd1 vccd1 vccd1 _06501_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07872__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14403_ clknet_leaf_138_clk _01108_ net1100 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11615_ _05755_ _05768_ _05769_ _05772_ vssd1 vssd1 vccd1 vccd1 _05839_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_13_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12595_ _06435_ _06436_ _06437_ vssd1 vssd1 vccd1 vccd1 _06443_ sky130_fd_sc_hd__a21boi_2
XFILLER_11_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14334_ clknet_leaf_1_clk _01039_ net1062 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07085__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11546_ screen.counter.ct\[3\] _05761_ vssd1 vssd1 vccd1 vccd1 _05770_ sky130_fd_sc_hd__or2_2
XANTENNA__07624__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14265_ clknet_leaf_29_clk _00970_ net1131 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_11477_ _05517_ _05734_ vssd1 vssd1 vccd1 vccd1 _05735_ sky130_fd_sc_hd__nand2_4
XANTENNA__12316__A net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13216_ clknet_leaf_137_clk _00026_ net1098 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_125_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10428_ net325 _04135_ _05255_ _05263_ vssd1 vssd1 vccd1 vccd1 _05264_ sky130_fd_sc_hd__o211ai_1
X_14196_ clknet_leaf_65_clk datapath.multiplication_module.multiplicand_i_n\[7\] net1237
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[7\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__08585__B1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13147_ net1990 net238 net384 vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__mux2_1
XANTENNA__12750__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10359_ net227 _05190_ _05194_ vssd1 vssd1 vccd1 vccd1 _05195_ sky130_fd_sc_hd__and3_1
XANTENNA__07793__D1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13078_ net2321 net243 net386 vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_146_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11366__S net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12029_ _06071_ net1431 _06017_ vssd1 vssd1 vccd1 vccd1 _00729_ sky130_fd_sc_hd__mux2_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10695__A1 _03417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07570_ datapath.rf.registers\[17\]\[19\] net851 net797 datapath.rf.registers\[29\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_66_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06984__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13808__RESET_B net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09240_ net321 _03798_ vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__or2_1
XFILLER_22_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07863__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08407__C net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09171_ net344 _04004_ _04006_ vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_32_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12925__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08122_ _02943_ _02944_ _02957_ vssd1 vssd1 vccd1 vccd1 _02958_ sky130_fd_sc_hd__or3b_1
XANTENNA__07615__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08704__A _03008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10080__C1 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08053_ datapath.rf.registers\[6\]\[9\] net952 net934 vssd1 vssd1 vccd1 vccd1 _02889_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12226__A _06168_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07004_ datapath.rf.registers\[9\]\[31\] net703 net661 datapath.rf.registers\[5\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_131_Right_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_110_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1119_A net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08955_ _02467_ _02523_ net445 vssd1 vssd1 vccd1 vccd1 _03791_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout481_A _06556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11276__S net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout579_A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07906_ datapath.rf.registers\[11\]\[12\] net883 net794 datapath.rf.registers\[31\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__a22o_1
X_08886_ _01611_ _03720_ vssd1 vssd1 vccd1 vccd1 _03722_ sky130_fd_sc_hd__nand2_1
XFILLER_57_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07000__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07837_ _02669_ _02670_ _02672_ vssd1 vssd1 vccd1 vccd1 _02673_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_16_Left_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout746_A net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07768_ datapath.rf.registers\[1\]\[15\] net846 net837 datapath.rf.registers\[26\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__a22o_1
XANTENNA__06894__A _01712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09507_ net457 _04341_ _04342_ vssd1 vssd1 vccd1 vccd1 _04343_ sky130_fd_sc_hd__nor3_1
X_06719_ mmio.memload_or_instruction\[30\] mmio.memload_or_instruction\[31\] mmio.memload_or_instruction\[27\]
+ mmio.memload_or_instruction\[29\] vssd1 vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__and4b_1
XANTENNA__07839__C1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout534_X net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07699_ datapath.rf.registers\[23\]\[17\] net700 _02534_ net788 vssd1 vssd1 vccd1
+ vccd1 _02535_ sky130_fd_sc_hd__a211o_1
XFILLER_13_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09438_ _03438_ _04273_ vssd1 vssd1 vccd1 vccd1 _04274_ sky130_fd_sc_hd__xor2_1
XFILLER_24_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07854__A2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09056__A1 _03666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout701_X net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09369_ net904 _04179_ _04202_ _04204_ vssd1 vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__o211a_1
XANTENNA__12835__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11400_ net2119 net205 net412 vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__mux2_1
XANTENNA__07067__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_25_Left_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12380_ net2598 net133 _06337_ vssd1 vssd1 vccd1 vccd1 _00814_ sky130_fd_sc_hd__a21o_1
XANTENNA__08173__X _03009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11331_ net2449 net210 net414 vssd1 vssd1 vccd1 vccd1 _00376_ sky130_fd_sc_hd__mux2_1
XFILLER_4_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10355__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14050_ clknet_leaf_101_clk _00817_ net1228 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11262_ net217 net2154 net418 vssd1 vssd1 vccd1 vccd1 _00311_ sky130_fd_sc_hd__mux2_1
XFILLER_97_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13001_ net1770 net290 net391 vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__mux2_1
XANTENNA__08052__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10213_ net225 _05048_ net1295 vssd1 vssd1 vccd1 vccd1 _05049_ sky130_fd_sc_hd__a21o_1
XFILLER_97_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08031__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11193_ net237 net2231 net424 vssd1 vssd1 vccd1 vccd1 _00245_ sky130_fd_sc_hd__mux2_1
XANTENNA__10374__B1 net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10144_ net1263 _03748_ vssd1 vssd1 vccd1 vccd1 _04980_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08319__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11186__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_128_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_34_Left_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10075_ _04649_ _04663_ _01702_ _04647_ vssd1 vssd1 vccd1 vccd1 _04911_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_128_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13903_ clknet_leaf_43_clk net1361 net1149 vssd1 vssd1 vccd1 vccd1 keypad.debounce.debounce\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09531__A2 _03296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13834_ clknet_leaf_115_clk _00643_ net1195 vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_141_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13765_ clknet_leaf_81_clk _00574_ net1255 vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__dfrtp_1
X_10977_ net1875 net278 net437 vssd1 vssd1 vccd1 vccd1 _00042_ sky130_fd_sc_hd__mux2_1
XANTENNA__08098__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08508__B _01797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12716_ columns.count\[6\] _06538_ vssd1 vssd1 vccd1 vccd1 _06540_ sky130_fd_sc_hd__nand2_1
XANTENNA__07412__B net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13696_ clknet_leaf_138_clk _00506_ net1097 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07845__A2 _02680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12647_ datapath.mulitply_result\[23\] datapath.multiplication_module.multiplicand_i\[23\]
+ vssd1 vssd1 vccd1 vccd1 _06486_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_61_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12745__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07058__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12051__B1 _06018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11869__B net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12578_ _06425_ _06426_ _06427_ vssd1 vssd1 vccd1 vccd1 _06429_ sky130_fd_sc_hd__or3_1
XANTENNA__08524__A net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11529_ screen.counter.ct\[1\] screen.counter.ct\[0\] vssd1 vssd1 vccd1 vccd1 _05753_
+ sky130_fd_sc_hd__nand2b_2
X_14317_ clknet_leaf_131_clk _01022_ net1205 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08270__A2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold307 datapath.rf.registers\[4\]\[2\] vssd1 vssd1 vccd1 vccd1 net1655 sky130_fd_sc_hd__dlygate4sd3_1
Xhold318 datapath.rf.registers\[23\]\[14\] vssd1 vssd1 vccd1 vccd1 net1666 sky130_fd_sc_hd__dlygate4sd3_1
Xhold329 datapath.rf.registers\[1\]\[18\] vssd1 vssd1 vccd1 vccd1 net1677 sky130_fd_sc_hd__dlygate4sd3_1
X_14248_ clknet_leaf_60_clk _00953_ net1235 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11885__A _02934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14179_ clknet_leaf_47_clk _00934_ net1175 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08022__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12480__S net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout809 _01766_ vssd1 vssd1 vccd1 vccd1 net809 sky130_fd_sc_hd__clkbuf_8
XFILLER_140_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07230__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11096__S net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08740_ _03524_ _03525_ _03573_ _03522_ _03520_ vssd1 vssd1 vccd1 vccd1 _03576_ sky130_fd_sc_hd__a311o_1
Xhold1007 datapath.rf.registers\[2\]\[2\] vssd1 vssd1 vccd1 vccd1 net2355 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1018 datapath.rf.registers\[19\]\[4\] vssd1 vssd1 vccd1 vccd1 net2366 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10117__B1 net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1029 screen.counter.currentCt\[7\] vssd1 vssd1 vccd1 vccd1 net2377 sky130_fd_sc_hd__dlygate4sd3_1
X_08671_ _03506_ vssd1 vssd1 vccd1 vccd1 _03507_ sky130_fd_sc_hd__inv_2
XFILLER_94_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07622_ datapath.rf.registers\[29\]\[18\] net796 _02451_ _02453_ _02457_ vssd1 vssd1
+ vccd1 vccd1 _02458_ sky130_fd_sc_hd__a2111oi_1
XFILLER_94_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09090__A _02025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07603__A _02438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07553_ datapath.rf.registers\[19\]\[19\] net976 net928 vssd1 vssd1 vccd1 vccd1 _02389_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08089__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07297__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07484_ datapath.rf.registers\[2\]\[21\] net742 net698 datapath.rf.registers\[23\]\[21\]
+ _02314_ vssd1 vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__a221o_1
XANTENNA__07836__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09223_ _03508_ _03582_ _03507_ vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__a21oi_1
XFILLER_21_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1069_A net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07049__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12042__B1 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09154_ net311 _03989_ vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_79_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_3_0_clk_X clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08105_ datapath.rf.registers\[3\]\[8\] net988 net927 vssd1 vssd1 vccd1 vccd1 _02941_
+ sky130_fd_sc_hd__and3_1
XFILLER_148_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09085_ _03919_ _03920_ net368 vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__mux2_1
XANTENNA__08261__A2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08153__B net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08036_ _02868_ _02869_ _02870_ _02871_ vssd1 vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__or4_1
XFILLER_135_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold830 datapath.rf.registers\[6\]\[14\] vssd1 vssd1 vccd1 vccd1 net2178 sky130_fd_sc_hd__dlygate4sd3_1
Xhold841 datapath.rf.registers\[9\]\[31\] vssd1 vssd1 vccd1 vccd1 net2189 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout696_A net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold852 datapath.rf.registers\[23\]\[8\] vssd1 vssd1 vccd1 vccd1 net2200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold863 datapath.rf.registers\[15\]\[29\] vssd1 vssd1 vccd1 vccd1 net2211 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09210__A1 _03666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08013__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07992__B net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold874 datapath.rf.registers\[14\]\[15\] vssd1 vssd1 vccd1 vccd1 net2222 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap582 net583 vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__clkbuf_1
Xhold885 datapath.rf.registers\[31\]\[28\] vssd1 vssd1 vccd1 vccd1 net2233 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06889__A _01630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold896 datapath.rf.registers\[10\]\[21\] vssd1 vssd1 vccd1 vccd1 net2244 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07221__B1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09987_ _04821_ _04822_ vssd1 vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout484_X net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08938_ _03772_ _03773_ net461 vssd1 vssd1 vccd1 vccd1 _03774_ sky130_fd_sc_hd__mux2_1
XFILLER_85_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08869_ _02913_ _02961_ net446 vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout651_X net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout749_X net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10900_ _01463_ net618 _05644_ _05645_ vssd1 vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_4_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11880_ net135 _05950_ _05949_ vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__o21ai_1
XFILLER_17_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07072__X _01908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10831_ datapath.mulitply_result\[14\] net599 net619 vssd1 vssd1 vccd1 vccd1 _05587_
+ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout916_X net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10577__C _02125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13550_ clknet_leaf_0_clk _00360_ net1057 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12281__B1 _06253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10762_ datapath.mulitply_result\[4\] net599 net619 vssd1 vssd1 vccd1 vccd1 _05528_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__07827__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12501_ net205 net1895 net507 vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__mux2_1
XANTENNA__08047__C net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13481_ clknet_leaf_91_clk _00291_ net1232 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10693_ _01430_ _05459_ _05508_ net1013 _05455_ vssd1 vssd1 vccd1 vccd1 _05509_ sky130_fd_sc_hd__a32o_1
X_12432_ net1399 net131 _06363_ vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__a21o_1
XFILLER_8_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12363_ net893 _04664_ vssd1 vssd1 vccd1 vccd1 _06326_ sky130_fd_sc_hd__nor2_1
XANTENNA__08252__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14102_ clknet_leaf_111_clk _00868_ net1218 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_154_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11314_ datapath.rf.registers\[12\]\[5\] net294 net414 vssd1 vssd1 vccd1 vccd1 _00359_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07460__B1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12294_ datapath.PC\[10\] net308 _06274_ _06276_ vssd1 vssd1 vccd1 vccd1 _00789_
+ sky130_fd_sc_hd__a22o_1
XFILLER_5_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14033_ clknet_leaf_84_clk _00802_ net1260 vssd1 vssd1 vccd1 vccd1 datapath.PC\[23\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_4_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11245_ net300 net1891 net418 vssd1 vssd1 vccd1 vccd1 _00294_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08004__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10898__A1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11176_ net287 net1591 net425 vssd1 vssd1 vccd1 vccd1 _00228_ sky130_fd_sc_hd__mux2_1
XFILLER_110_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08960__A0 _02660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10127_ net225 _04877_ _04962_ net1294 vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__a31oi_1
XANTENNA__07407__B net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10058_ _04718_ _04828_ _04717_ vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_34_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13817_ clknet_leaf_115_clk _00626_ net1189 vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__dfrtp_1
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07279__B1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07818__A2 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13748_ clknet_leaf_88_clk _00557_ net1252 vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__dfrtp_1
XFILLER_149_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13679_ clknet_leaf_25_clk _00489_ net1138 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06981__B _01816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold104 net53 vssd1 vssd1 vccd1 vccd1 net1452 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold115 net83 vssd1 vssd1 vccd1 vccd1 net1463 sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 net79 vssd1 vssd1 vccd1 vccd1 net1474 sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 net88 vssd1 vssd1 vccd1 vccd1 net1485 sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 mmio.memload_or_instruction\[7\] vssd1 vssd1 vccd1 vccd1 net1496 sky130_fd_sc_hd__dlygate4sd3_1
X_09910_ datapath.PC\[14\] _04744_ vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__xor2_2
Xhold159 net80 vssd1 vssd1 vccd1 vccd1 net1507 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout606 _03610_ vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__clkbuf_2
Xfanout617 net618 vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__buf_2
XANTENNA__07203__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09841_ _03558_ _04675_ _04676_ vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__or3_1
XFILLER_113_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout628 net629 vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__clkbuf_2
Xfanout639 net641 vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkload14_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07317__B net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09772_ _03468_ _03492_ vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__xnor2_1
X_06984_ net991 _01637_ net990 _01666_ vssd1 vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__and4_1
XANTENNA__06996__X _01832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08723_ _03557_ _03558_ _03542_ vssd1 vssd1 vccd1 vccd1 _03559_ sky130_fd_sc_hd__a21o_1
XANTENNA__07036__C net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout277_A _05558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08654_ _02070_ _02091_ vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__nor2_1
XFILLER_94_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07605_ _02418_ _02440_ vssd1 vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_105_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08585_ net559 _03358_ net558 _03419_ vssd1 vssd1 vccd1 vccd1 _03421_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_105_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1186_A _00004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07536_ datapath.rf.registers\[28\]\[20\] net752 net728 datapath.rf.registers\[25\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__a22o_1
XANTENNA__07809__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07467_ datapath.rf.registers\[4\]\[21\] net864 _02290_ _02291_ _02292_ vssd1 vssd1
+ vccd1 vccd1 _02303_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout611_A _01782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09206_ net456 _03843_ _03844_ _03886_ net353 vssd1 vssd1 vccd1 vccd1 _04042_ sky130_fd_sc_hd__a311oi_2
XFILLER_139_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07690__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07398_ datapath.rf.registers\[7\]\[23\] net671 net664 datapath.rf.registers\[15\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__a22o_1
XFILLER_154_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09137_ _03498_ net627 net624 _03499_ net644 vssd1 vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__a221oi_1
XTAP_TAPCELL_ROW_20_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08234__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07442__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09068_ _03903_ vssd1 vssd1 vccd1 vccd1 _03904_ sky130_fd_sc_hd__inv_2
XFILLER_135_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout699_X net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08019_ _02846_ _02850_ _02854_ vssd1 vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__or3_4
XFILLER_118_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11956__C net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold660 datapath.rf.registers\[30\]\[6\] vssd1 vssd1 vccd1 vccd1 net2008 sky130_fd_sc_hd__dlygate4sd3_1
Xhold671 datapath.rf.registers\[22\]\[18\] vssd1 vssd1 vccd1 vccd1 net2019 sky130_fd_sc_hd__dlygate4sd3_1
X_11030_ net193 net2317 net538 vssd1 vssd1 vccd1 vccd1 _00092_ sky130_fd_sc_hd__mux2_1
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold682 datapath.rf.registers\[8\]\[6\] vssd1 vssd1 vccd1 vccd1 net2030 sky130_fd_sc_hd__dlygate4sd3_1
Xhold693 datapath.rf.registers\[19\]\[21\] vssd1 vssd1 vccd1 vccd1 net2041 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout866_X net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09282__X _04118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09723__A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12981_ net235 net2236 net480 vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__mux2_1
XANTENNA__11464__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09498__B2 _03614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11932_ net2556 net162 vssd1 vssd1 vccd1 vccd1 _05985_ sky130_fd_sc_hd__nand2_1
XANTENNA__10588__B _02090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11863_ net2514 net163 vssd1 vssd1 vccd1 vccd1 _05939_ sky130_fd_sc_hd__nand2_1
X_14651_ clknet_leaf_37_clk _01356_ net1136 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10814_ _05571_ vssd1 vssd1 vccd1 vccd1 _05572_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_28_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13602_ clknet_leaf_152_clk _00412_ net1054 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11794_ _01500_ net1014 net313 net333 datapath.ru.latched_instruction\[0\] vssd1
+ vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__a32o_1
X_14582_ clknet_leaf_137_clk _01287_ net1097 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10745_ net1530 net569 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[31\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__12295__S net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13533_ clknet_leaf_144_clk _00343_ net1085 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10280__A2 net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12006__B1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13464_ clknet_leaf_4_clk _00274_ net1069 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10676_ net1013 _05436_ _05490_ _05430_ vssd1 vssd1 vccd1 vccd1 _05494_ sky130_fd_sc_hd__o31a_1
X_12415_ _05972_ net158 vssd1 vssd1 vccd1 vccd1 _06355_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_136_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08225__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09422__A1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13395_ clknet_leaf_35_clk _00205_ net1129 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_153_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12346_ datapath.PC\[25\] _06313_ net306 vssd1 vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__mux2_1
XANTENNA__07433__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08802__A _01603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12277_ _05537_ _06254_ _06263_ vssd1 vssd1 vccd1 vccd1 _06264_ sky130_fd_sc_hd__o21ai_1
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14016_ clknet_leaf_86_clk _00785_ net1254 vssd1 vssd1 vccd1 vccd1 datapath.PC\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11228_ net233 net1583 net526 vssd1 vssd1 vccd1 vccd1 _00278_ sky130_fd_sc_hd__mux2_1
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08933__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11159_ net220 net2013 net530 vssd1 vssd1 vccd1 vccd1 _00212_ sky130_fd_sc_hd__mux2_1
XFILLER_110_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11882__B net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09489__A1 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11374__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10498__B _05315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08370_ _01649_ _01703_ _01783_ _01647_ vssd1 vssd1 vccd1 vccd1 _03206_ sky130_fd_sc_hd__a22o_1
X_07321_ datapath.rf.registers\[16\]\[24\] net861 net857 datapath.rf.registers\[24\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__a22o_1
XFILLER_149_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07252_ datapath.rf.registers\[24\]\[26\] net766 net742 datapath.rf.registers\[2\]\[26\]
+ _02077_ vssd1 vssd1 vccd1 vccd1 _02088_ sky130_fd_sc_hd__a221o_1
XANTENNA__07672__B1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07183_ datapath.rf.registers\[24\]\[27\] net857 _02005_ _02017_ _02018_ vssd1 vssd1
+ vccd1 vccd1 _02019_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08216__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12933__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14022__RESET_B net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08712__A net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12234__A _06168_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08431__B net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout403 _06549_ vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09716__A2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout414 _05726_ vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__clkbuf_8
Xfanout425 _05719_ vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__buf_4
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11523__A2 _05747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout394_A _06555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08150__C net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout436 net437 vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08924__B1 _03759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout447 _03679_ vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__clkbuf_4
X_09824_ _03481_ net627 _04659_ net645 vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout1101_A net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout458 _03652_ vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__buf_2
XFILLER_98_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout469 _01701_ vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__buf_4
XFILLER_86_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_107_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09755_ net649 _04590_ net438 vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__a21o_1
XFILLER_74_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06967_ net968 net911 _01795_ vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__and3_1
XANTENNA__11284__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06886__B _01712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07334__Y _02170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08706_ net464 _03126_ vssd1 vssd1 vccd1 vccd1 _03542_ sky130_fd_sc_hd__nor2_1
X_09686_ _04134_ _04521_ net359 vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__mux2_1
XFILLER_73_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06898_ datapath.rf.registers\[8\]\[31\] net877 net853 datapath.rf.registers\[19\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_87_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08637_ _03471_ _03472_ _01957_ vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__a21o_1
XFILLER_55_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_120_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout826_A net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout447_X net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08568_ datapath.rf.registers\[18\]\[0\] net910 _01805_ vssd1 vssd1 vccd1 vccd1 _03404_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_25_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07519_ datapath.rf.registers\[10\]\[20\] net879 net849 datapath.rf.registers\[17\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__a22o_1
X_08499_ datapath.rf.registers\[27\]\[1\] net965 _01816_ vssd1 vssd1 vccd1 vccd1 _03335_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09652__A1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout614_X net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13004__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10530_ screen.counter.ct\[9\] _05359_ vssd1 vssd1 vccd1 vccd1 _05360_ sky130_fd_sc_hd__nand2_1
XANTENNA__07510__B net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10574__D _03149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10461_ keypad.decode.sticky\[4\] keypad.decode.sticky\[3\] net1022 vssd1 vssd1 vccd1
+ vccd1 keypad.decode.sticky_n\[3\] sky130_fd_sc_hd__mux2_1
XANTENNA__08207__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12843__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12200_ net2335 _06209_ net603 vssd1 vssd1 vccd1 vccd1 _06211_ sky130_fd_sc_hd__o21ai_1
XFILLER_109_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07415__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13180_ datapath.rf.registers\[0\]\[17\] vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__clkbuf_1
X_10392_ net460 _05226_ net351 vssd1 vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__a21oi_1
XFILLER_89_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout983_X net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12131_ screen.counter.currentEnable _06167_ vssd1 vssd1 vccd1 vccd1 _06168_ sky130_fd_sc_hd__nor2_4
XANTENNA__11459__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10216__X _05052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10970__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08341__B net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12062_ _05858_ _06089_ _06094_ _06102_ vssd1 vssd1 vccd1 vccd1 _06103_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_78_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold490 datapath.rf.registers\[18\]\[9\] vssd1 vssd1 vccd1 vccd1 net1838 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08060__C net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11013_ net275 datapath.rf.registers\[27\]\[9\] net540 vssd1 vssd1 vccd1 vccd1 _00075_
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_8_Left_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07194__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout970 net971 vssd1 vssd1 vccd1 vccd1 net970 sky130_fd_sc_hd__buf_2
Xfanout981 net983 vssd1 vssd1 vccd1 vccd1 net981 sky130_fd_sc_hd__clkbuf_4
XFILLER_77_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout992 _01632_ vssd1 vssd1 vccd1 vccd1 net992 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_51_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11194__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06941__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12964_ net289 net2094 net481 vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__mux2_1
XANTENNA__11817__A3 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1190 datapath.mulitply_result\[3\] vssd1 vssd1 vccd1 vccd1 net2538 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11915_ _02438_ screen.counter.ack vssd1 vssd1 vccd1 vccd1 _05974_ sky130_fd_sc_hd__or2_1
XANTENNA__10886__X _05634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12895_ _05517_ _05693_ vssd1 vssd1 vccd1 vccd1 _06554_ sky130_fd_sc_hd__and2_2
XFILLER_61_857 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14634_ clknet_leaf_21_clk _01339_ net1164 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11846_ _05795_ _05912_ _05924_ _05752_ vssd1 vssd1 vccd1 vccd1 _05925_ sky130_fd_sc_hd__a22o_1
XFILLER_54_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_11_0_clk_X clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11777_ net121 _05483_ _05894_ vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__mux2_1
X_14565_ clknet_leaf_118_clk _01270_ net1191 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08516__B net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13516_ clknet_leaf_16_clk _00326_ net1106 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10728_ net1553 _02660_ net573 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[14\]
+ sky130_fd_sc_hd__mux2_1
X_14496_ clknet_leaf_137_clk _01201_ net1090 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10659_ net1037 _05474_ _05475_ _05477_ vssd1 vssd1 vccd1 vccd1 _05478_ sky130_fd_sc_hd__a211o_1
X_13447_ clknet_leaf_137_clk _00257_ net1089 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12753__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload13 clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clkload13/Y sky130_fd_sc_hd__clkinv_8
Xclkload24 clknet_leaf_152_clk vssd1 vssd1 vccd1 vccd1 clkload24/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload35 clknet_leaf_136_clk vssd1 vssd1 vccd1 vccd1 clkload35/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_58_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09187__X _04023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload46 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 clkload46/X sky130_fd_sc_hd__clkbuf_8
X_13378_ clknet_leaf_150_clk _00188_ net1053 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06604__X _01443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload57 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 clkload57/Y sky130_fd_sc_hd__inv_8
Xclkload68 clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 clkload68/Y sky130_fd_sc_hd__inv_8
XANTENNA__11369__S net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload79 clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 clkload79/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_141_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12329_ datapath.PC\[20\] net310 _06301_ vssd1 vssd1 vccd1 vccd1 _00799_ sky130_fd_sc_hd__a21o_1
XANTENNA__09159__B1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07870_ datapath.rf.registers\[25\]\[13\] net727 net719 datapath.rf.registers\[20\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__a22o_1
XANTENNA__06987__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07185__A2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06821_ net1002 net1018 _01654_ net1026 datapath.ru.latched_instruction\[16\] vssd1
+ vssd1 vccd1 vccd1 _01657_ sky130_fd_sc_hd__a32oi_4
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09540_ net464 net463 net441 vssd1 vssd1 vccd1 vccd1 _04376_ sky130_fd_sc_hd__mux2_1
XFILLER_110_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06752_ _01572_ _01589_ vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__nor2_1
XFILLER_48_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09650__X _04486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09471_ _02961_ _03009_ net452 vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__mux2_1
X_06683_ datapath.ru.latched_instruction\[17\] _01452_ _01506_ datapath.ru.latched_instruction\[21\]
+ vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__a22o_1
XANTENNA__07314__C net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07342__C1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08422_ datapath.rf.registers\[10\]\[2\] net881 net852 datapath.rf.registers\[17\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03258_ sky130_fd_sc_hd__a22o_1
XANTENNA__08707__A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08353_ datapath.rf.registers\[8\]\[3\] net956 _01712_ vssd1 vssd1 vccd1 vccd1 _03189_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout142_A _05891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09634__A1 _03673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14203__RESET_B net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07304_ datapath.rf.registers\[4\]\[25\] net716 net662 datapath.rf.registers\[5\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__a22o_1
XFILLER_138_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10244__A2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07645__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08284_ datapath.rf.registers\[14\]\[5\] net775 net688 datapath.rf.registers\[31\]\[5\]
+ _03119_ vssd1 vssd1 vccd1 vccd1 _03120_ sky130_fd_sc_hd__a221o_1
Xclkload7 clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clkload7/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_149_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07235_ datapath.rf.registers\[22\]\[26\] net734 net668 datapath.rf.registers\[21\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02071_ sky130_fd_sc_hd__a22o_1
XFILLER_149_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout407_A _05733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire951_X net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07166_ _02001_ vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__inv_2
XANTENNA__11279__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07097_ _01922_ _01926_ _01929_ _01932_ vssd1 vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__nor4_1
XTAP_TAPCELL_ROW_113_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout200 net202 vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__clkbuf_2
Xfanout211 net213 vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__clkbuf_2
Xfanout1209 net1210 vssd1 vssd1 vccd1 vccd1 net1209 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout776_A _01796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout397_X net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout222 _04713_ vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__buf_2
Xfanout233 net234 vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__clkbuf_2
Xfanout244 net246 vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout255 net257 vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06897__A net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout266 net267 vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09807_ _03607_ _04629_ _04642_ net605 vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__a211oi_1
Xfanout277 _05558_ vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout288 _05706_ vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__clkbuf_2
XFILLER_46_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout299 net301 vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__clkbuf_2
X_07999_ datapath.rf.registers\[7\]\[10\] net941 net935 vssd1 vssd1 vccd1 vccd1 _02835_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout564_X net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout943_A _01715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07505__B net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09738_ net381 _03768_ _04573_ _03614_ vssd1 vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__a211o_1
XANTENNA__09322__A0 _02419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout731_X net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09669_ net329 _04504_ vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__or2_1
XANTENNA__12838__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09873__A1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout829_X net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11700_ _05061_ net154 net149 net1402 vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__a22o_1
XANTENNA__11680__A1 _05116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12680_ _06512_ _06513_ vssd1 vssd1 vccd1 vccd1 _06514_ sky130_fd_sc_hd__nand2_1
XANTENNA__07884__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11631_ _05751_ _05853_ vssd1 vssd1 vccd1 vccd1 _05855_ sky130_fd_sc_hd__nor2_1
XFILLER_42_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09625__A1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10585__C _03123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_145_Right_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07636__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14350_ clknet_leaf_1_clk _01055_ net1062 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11562_ net1006 _05785_ vssd1 vssd1 vccd1 vccd1 _05786_ sky130_fd_sc_hd__nor2_4
XANTENNA__07100__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10513_ screen.controlBus\[4\] screen.controlBus\[5\] _05314_ _05327_ vssd1 vssd1
+ vccd1 vccd1 _05343_ sky130_fd_sc_hd__and4b_2
X_13301_ clknet_leaf_133_clk _00111_ net1111 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08055__C net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14281_ clknet_leaf_91_clk _00986_ net1232 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_11493_ net248 net2051 net510 vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_133_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13232_ clknet_leaf_24_clk _00042_ net1155 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10444_ _04839_ _05279_ net1254 vssd1 vssd1 vccd1 vccd1 _05280_ sky130_fd_sc_hd__o21ai_1
XFILLER_136_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07894__C net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11735__A2 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11189__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13163_ net2344 vssd1 vssd1 vccd1 vccd1 _00985_ sky130_fd_sc_hd__clkbuf_1
X_10375_ net1269 net1292 _05209_ _05210_ vssd1 vssd1 vccd1 vccd1 _05211_ sky130_fd_sc_hd__a22o_1
XFILLER_124_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10943__B1 _05682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12114_ screen.counter.currentCt\[10\] _06148_ _06150_ vssd1 vssd1 vccd1 vccd1 _06151_
+ sky130_fd_sc_hd__or3_1
XFILLER_151_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13094_ _05518_ _05725_ vssd1 vssd1 vccd1 vccd1 _06561_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_53_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12045_ _05332_ _06081_ _06086_ _06044_ _06075_ vssd1 vssd1 vccd1 vccd1 _06087_ sky130_fd_sc_hd__a2111o_1
XFILLER_78_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07167__A2 _02001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06914__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12448__B1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13996_ clknet_leaf_112_clk _00773_ net1197 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12947_ net221 net2142 net394 vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__mux2_1
XANTENNA__12748__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11671__A1 _05240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06678__B2 datapath.ru.latched_instruction\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__07875__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12878_ net249 net2247 net399 vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__mux2_1
XFILLER_21_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14617_ clknet_leaf_8_clk _01322_ net1072 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_11829_ net1274 screen.counter.ct\[17\] _05907_ vssd1 vssd1 vccd1 vccd1 _05908_ sky130_fd_sc_hd__and3_1
XANTENNA__08419__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09077__C1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08246__B net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07627__B1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14548_ clknet_leaf_128_clk _01253_ net1209 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_112_Right_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11888__A _02876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12483__S net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload102 clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 clkload102/Y sky130_fd_sc_hd__clkinv_8
X_14479_ clknet_leaf_26_clk _01184_ net1158 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload113 clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 clkload113/Y sky130_fd_sc_hd__bufinv_16
X_07020_ net610 _01854_ _01787_ vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__o21ai_1
Xclkload124 clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 clkload124/Y sky130_fd_sc_hd__inv_12
Xclkload135 clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 clkload135/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__06850__B2 datapath.ru.latched_instruction\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xclkload146 clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 clkload146/Y sky130_fd_sc_hd__inv_6
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11726__A2 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11099__S net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08971_ _03802_ _03806_ net340 vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__mux2_1
XFILLER_103_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07922_ datapath.rf.registers\[3\]\[12\] net771 net715 datapath.rf.registers\[4\]\[12\]
+ _02757_ vssd1 vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__a221o_1
Xhold19 keypad.debounce.debounce\[5\] vssd1 vssd1 vccd1 vccd1 net1367 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07158__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07165__X _02001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07853_ datapath.rf.registers\[2\]\[13\] net887 net885 datapath.rf.registers\[9\]\[13\]
+ _02688_ vssd1 vssd1 vccd1 vccd1 _02689_ sky130_fd_sc_hd__a221o_1
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07606__A _02418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06804_ _01474_ net1016 net994 net1030 datapath.ru.latched_instruction\[11\] vssd1
+ vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__a32oi_4
XFILLER_84_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07784_ datapath.rf.registers\[8\]\[15\] net695 net688 datapath.rf.registers\[31\]\[15\]
+ _02619_ vssd1 vssd1 vccd1 vccd1 _02620_ sky130_fd_sc_hd__a221o_1
XFILLER_72_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09523_ net352 _03993_ _04358_ vssd1 vssd1 vccd1 vccd1 _04359_ sky130_fd_sc_hd__o21a_1
X_06735_ _01441_ _01564_ net1021 net1030 datapath.ru.latched_instruction\[5\] vssd1
+ vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__a32o_1
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09454_ _04257_ _04289_ net367 vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__mux2_1
X_06666_ mmio.memload_or_instruction\[21\] net1049 vssd1 vssd1 vccd1 vccd1 _01505_
+ sky130_fd_sc_hd__and2_2
XFILLER_101_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10686__B _01435_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07330__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08405_ datapath.rf.registers\[22\]\[2\] net953 net926 vssd1 vssd1 vccd1 vccd1 _03241_
+ sky130_fd_sc_hd__and3_1
XFILLER_40_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09385_ net360 _03998_ _03999_ vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__nor3_1
X_06597_ net1294 vssd1 vssd1 vccd1 vccd1 _00004_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout524_A _05723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08336_ _03171_ vssd1 vssd1 vccd1 vccd1 _03172_ sky130_fd_sc_hd__inv_2
XFILLER_137_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08267_ _03089_ _03093_ _03102_ vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__or3_2
XANTENNA__07995__B net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10906__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_140_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_140_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_20_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07218_ datapath.rf.registers\[20\]\[26\] net957 net921 vssd1 vssd1 vccd1 vccd1 _02054_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_115_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08198_ datapath.rf.registers\[10\]\[6\] net879 net856 datapath.rf.registers\[24\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03034_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout893_A net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_89_Left_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07149_ datapath.rf.registers\[17\]\[28\] net749 net705 datapath.rf.registers\[9\]\[28\]
+ _01982_ vssd1 vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__a221o_1
XFILLER_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07397__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10160_ _04993_ _04995_ net225 vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__mux2_1
XANTENNA__12390__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout681_X net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1006 _05756_ vssd1 vssd1 vccd1 vccd1 net1006 sky130_fd_sc_hd__buf_4
XANTENNA_fanout779_X net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1017 _01562_ vssd1 vssd1 vccd1 vccd1 net1017 sky130_fd_sc_hd__clkbuf_4
X_10091_ net641 _03916_ _04607_ vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__and3_1
Xfanout1028 net1032 vssd1 vssd1 vccd1 vccd1 net1028 sky130_fd_sc_hd__buf_4
Xfanout1039 net1042 vssd1 vssd1 vccd1 vccd1 net1039 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07149__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12142__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout946_X net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13850_ clknet_leaf_49_clk _00654_ net1177 vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__dfstp_1
XFILLER_142_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_98_Left_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12801_ net1630 net299 net491 vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__mux2_1
XFILLER_142_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13781_ clknet_leaf_51_clk _00590_ net1182 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10993_ net1703 net199 net434 vssd1 vssd1 vccd1 vccd1 _00058_ sky130_fd_sc_hd__mux2_1
XANTENNA__11472__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07857__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12732_ net1551 net258 net405 vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_52_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07321__A2 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12663_ _06497_ _06498_ _06499_ vssd1 vssd1 vccd1 vccd1 _06500_ sky130_fd_sc_hd__or3_1
XFILLER_31_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14402_ clknet_leaf_1_clk _01107_ net1056 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11614_ _05758_ _05761_ _05764_ vssd1 vssd1 vccd1 vccd1 _05838_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_46_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12594_ _06440_ _06441_ vssd1 vssd1 vccd1 vccd1 _06442_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14333_ clknet_leaf_147_clk _01038_ net1064 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11545_ net1008 _05764_ vssd1 vssd1 vccd1 vccd1 _05769_ sky130_fd_sc_hd__nor2_2
XFILLER_11_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08282__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_131_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_131_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_67_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13760__RESET_B net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14264_ clknet_leaf_3_clk _00969_ net1077 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11476_ _05513_ _05689_ vssd1 vssd1 vccd1 vccd1 _05734_ sky130_fd_sc_hd__nor2_2
XANTENNA_clkbuf_leaf_110_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11708__A2 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10427_ net647 _05262_ _03667_ vssd1 vssd1 vccd1 vccd1 _05263_ sky130_fd_sc_hd__o21ai_1
X_13215_ clknet_leaf_11_clk _00025_ net1082 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08034__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14195_ clknet_leaf_66_clk datapath.multiplication_module.multiplicand_i_n\[6\] net1236
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[6\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__07388__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08585__A1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13146_ net1614 net220 net382 vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__mux2_1
X_10358_ net1039 _05191_ _05193_ net634 vssd1 vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__a211o_1
XFILLER_97_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13077_ net1688 net247 net387 vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_125_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10404__X _05240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10289_ _05122_ _05124_ net224 vssd1 vssd1 vccd1 vccd1 _05125_ sky130_fd_sc_hd__mux2_1
XANTENNA__09534__A0 _02705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12028_ _05847_ _06069_ _06070_ vssd1 vssd1 vccd1 vccd1 _06071_ sky130_fd_sc_hd__o21a_1
XFILLER_54_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12478__S net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13979_ clknet_leaf_107_clk _00757_ net1221 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[22\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__11382__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06984__B _01637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07312__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09170_ net344 _04005_ vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_32_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08121_ datapath.rf.registers\[17\]\[8\] net852 _02938_ _02941_ _02942_ vssd1 vssd1
+ vccd1 vccd1 _02957_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__08273__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_122_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_122_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10726__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13102__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08052_ datapath.rf.registers\[23\]\[9\] net941 net924 vssd1 vssd1 vccd1 vccd1 _02888_
+ sky130_fd_sc_hd__and3_1
X_07003_ _01833_ _01836_ _01837_ _01838_ vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__or4_1
XANTENNA__08025__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12941__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07379__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10383__A1 _03383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12242__A _06168_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08954_ _03789_ vssd1 vssd1 vccd1 vccd1 _03790_ sky130_fd_sc_hd__inv_2
XFILLER_57_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07905_ datapath.rf.registers\[24\]\[12\] net859 _02736_ _02740_ vssd1 vssd1 vccd1
+ vccd1 _02741_ sky130_fd_sc_hd__a211oi_2
XFILLER_102_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08885_ _01611_ _03720_ vssd1 vssd1 vccd1 vccd1 _03721_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout474_A net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07836_ datapath.rf.registers\[24\]\[14\] net767 net702 datapath.rf.registers\[9\]\[14\]
+ _02671_ vssd1 vssd1 vccd1 vccd1 _02672_ sky130_fd_sc_hd__a221o_1
XFILLER_72_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07767_ datapath.rf.registers\[13\]\[15\] net811 net802 datapath.rf.registers\[3\]\[15\]
+ _02594_ vssd1 vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__a221o_1
XFILLER_84_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11292__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06894__B net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout739_A net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09506_ net554 net550 net560 vssd1 vssd1 vccd1 vccd1 _04342_ sky130_fd_sc_hd__o21a_1
X_06718_ _01449_ _01485_ _01500_ vssd1 vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__or3b_1
X_07698_ datapath.rf.registers\[1\]\[17\] net764 net662 datapath.rf.registers\[5\]\[17\]
+ _02533_ vssd1 vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__a221o_1
XANTENNA__07303__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06649_ _01445_ _01458_ _01473_ _01487_ vssd1 vssd1 vccd1 vccd1 _01488_ sky130_fd_sc_hd__or4bb_1
XANTENNA__10843__C1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09437_ _03531_ _03532_ vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__nand2_2
XANTENNA__07502__C net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout527_X net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09368_ net324 _03715_ _04203_ vssd1 vssd1 vccd1 vccd1 _04204_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_10_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08264__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08319_ datapath.rf.registers\[3\]\[4\] net771 net763 datapath.rf.registers\[1\]\[4\]
+ _03153_ vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__a221o_1
XFILLER_21_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_113_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_113_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09299_ _03888_ _04134_ net361 vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__mux2_1
XANTENNA__13012__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11330_ net1700 net214 net414 vssd1 vssd1 vccd1 vccd1 _00375_ sky130_fd_sc_hd__mux2_1
XANTENNA__06814__B2 datapath.ru.latched_instruction\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_126_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout896_X net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11261_ net232 net2371 net418 vssd1 vssd1 vccd1 vccd1 _00310_ sky130_fd_sc_hd__mux2_1
XANTENNA__08016__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12851__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10212_ _04868_ _04869_ vssd1 vssd1 vccd1 vccd1 _05048_ sky130_fd_sc_hd__xnor2_1
X_13000_ net1793 net294 net390 vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__mux2_1
XFILLER_122_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11192_ net218 net2103 net422 vssd1 vssd1 vccd1 vccd1 _00244_ sky130_fd_sc_hd__mux2_1
XANTENNA__10374__A1 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11467__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10143_ datapath.PC\[26\] net468 net1039 vssd1 vssd1 vccd1 vccd1 _04979_ sky130_fd_sc_hd__o21a_1
XFILLER_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07790__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input35_A gpio_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10074_ _04626_ _04645_ _04664_ vssd1 vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_128_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13902_ clknet_leaf_43_clk net1364 net1150 vssd1 vssd1 vccd1 vccd1 keypad.debounce.debounce\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11874__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07542__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13833_ clknet_leaf_113_clk _00642_ net1196 vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13764_ clknet_leaf_81_clk _00573_ net1256 vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__dfrtp_1
X_10976_ net1814 net282 net436 vssd1 vssd1 vccd1 vccd1 _00041_ sky130_fd_sc_hd__mux2_1
X_12715_ columns.count\[6\] _06538_ vssd1 vssd1 vccd1 vccd1 _06539_ sky130_fd_sc_hd__or2_1
XANTENNA__08508__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10894__X _05641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07412__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13695_ clknet_leaf_10_clk _00505_ net1080 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_148_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12646_ net498 _06484_ _06485_ net502 datapath.mulitply_result\[22\] vssd1 vssd1
+ vccd1 vccd1 _00932_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_61_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_104_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_104_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08255__B1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12577_ _06426_ _06427_ _06425_ vssd1 vssd1 vccd1 vccd1 _06428_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08524__B _03358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14316_ clknet_leaf_16_clk _01021_ net1103 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11528_ net1009 _05751_ vssd1 vssd1 vccd1 vccd1 _05752_ sky130_fd_sc_hd__or2_1
XFILLER_117_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_886 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold308 datapath.rf.registers\[24\]\[1\] vssd1 vssd1 vccd1 vccd1 net1656 sky130_fd_sc_hd__dlygate4sd3_1
Xhold319 datapath.rf.registers\[20\]\[28\] vssd1 vssd1 vccd1 vccd1 net1667 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08007__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14247_ clknet_leaf_94_clk datapath.multiplication_module.multiplier_i_n\[15\] net1217
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i\[15\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12761__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11459_ net2222 net248 net407 vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__mux2_1
XFILLER_125_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12354__A2 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11885__B net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14178_ clknet_leaf_48_clk _00933_ net1177 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[23\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__11377__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13129_ net1731 net259 net385 vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__mux2_1
XFILLER_30_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07781__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1008 datapath.rf.registers\[11\]\[13\] vssd1 vssd1 vccd1 vccd1 net2356 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10117__A1 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1019 datapath.rf.registers\[6\]\[24\] vssd1 vssd1 vccd1 vccd1 net2367 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08670_ _02387_ _03456_ vssd1 vssd1 vccd1 vccd1 _03506_ sky130_fd_sc_hd__and2b_1
XANTENNA__06995__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07533__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07621_ _02454_ _02455_ _02456_ vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__or3_1
XFILLER_19_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07552_ datapath.rf.registers\[3\]\[19\] net985 net928 vssd1 vssd1 vccd1 vccd1 _02388_
+ sky130_fd_sc_hd__and3_1
X_07483_ datapath.rf.registers\[25\]\[21\] net726 net687 datapath.rf.registers\[31\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__a22o_1
XANTENNA__12290__B2 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12936__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09222_ _03453_ _03507_ vssd1 vssd1 vccd1 vccd1 _04058_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09153_ net376 _03988_ _03984_ net380 vssd1 vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__a211o_1
XFILLER_21_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08104_ datapath.rf.registers\[6\]\[8\] net825 net818 datapath.rf.registers\[7\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__a22o_1
XANTENNA__08434__B net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09084_ _02125_ _02169_ net443 vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08035_ datapath.rf.registers\[16\]\[10\] net740 net720 datapath.rf.registers\[20\]\[10\]
+ _02861_ vssd1 vssd1 vccd1 vccd1 _02871_ sky130_fd_sc_hd__a221o_1
XANTENNA__08153__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold820 datapath.rf.registers\[11\]\[9\] vssd1 vssd1 vccd1 vccd1 net2168 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1131_A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold831 datapath.rf.registers\[0\]\[26\] vssd1 vssd1 vccd1 vccd1 net2179 sky130_fd_sc_hd__dlygate4sd3_1
Xhold842 datapath.rf.registers\[30\]\[29\] vssd1 vssd1 vccd1 vccd1 net2190 sky130_fd_sc_hd__dlygate4sd3_1
Xhold853 datapath.rf.registers\[26\]\[29\] vssd1 vssd1 vccd1 vccd1 net2201 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07992__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold864 datapath.rf.registers\[28\]\[3\] vssd1 vssd1 vccd1 vccd1 net2212 sky130_fd_sc_hd__dlygate4sd3_1
Xhold875 datapath.rf.registers\[26\]\[26\] vssd1 vssd1 vccd1 vccd1 net2223 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold886 datapath.rf.registers\[8\]\[16\] vssd1 vssd1 vccd1 vccd1 net2234 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11287__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout689_A net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold897 datapath.rf.registers\[23\]\[31\] vssd1 vssd1 vccd1 vccd1 net2245 sky130_fd_sc_hd__dlygate4sd3_1
X_09986_ datapath.PC\[25\] net594 vssd1 vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout1017_X net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07772__A2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08937_ _01935_ _01981_ net453 vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout856_A net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout477_X net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08221__A2_N net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08868_ _02805_ _02857_ net444 vssd1 vssd1 vccd1 vccd1 _03704_ sky130_fd_sc_hd__mux2_1
XANTENNA__07353__X _02189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07524__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07819_ datapath.rf.registers\[11\]\[14\] net883 net855 datapath.rf.registers\[19\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02655_ sky130_fd_sc_hd__a22o_1
XFILLER_45_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08799_ net379 _03634_ vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout644_X net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13007__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10830_ _04239_ _05585_ net899 vssd1 vssd1 vccd1 vccd1 _05586_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_123_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10577__D _02169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12281__A1 _05002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12846__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout811_X net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10761_ _04428_ _05526_ net899 vssd1 vssd1 vccd1 vccd1 _05527_ sky130_fd_sc_hd__mux2_1
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12500_ net211 net2470 net506 vssd1 vssd1 vccd1 vccd1 _00900_ sky130_fd_sc_hd__mux2_1
XFILLER_12_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10692_ _05433_ _05449_ _05464_ vssd1 vssd1 vccd1 vccd1 _05508_ sky130_fd_sc_hd__a21o_1
XFILLER_12_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13480_ clknet_leaf_64_clk _00290_ net1236 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10831__A2 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08237__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12431_ _05988_ net158 vssd1 vssd1 vccd1 vccd1 _06363_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_101_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08344__B net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12362_ datapath.PC\[29\] net306 _06324_ _06325_ vssd1 vssd1 vccd1 vccd1 _00808_
+ sky130_fd_sc_hd__o22a_1
XFILLER_126_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14101_ clknet_leaf_112_clk _00867_ net1218 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11313_ net1782 net298 net414 vssd1 vssd1 vccd1 vccd1 _00358_ sky130_fd_sc_hd__mux2_1
XFILLER_126_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12293_ net190 _06275_ _06253_ _05561_ vssd1 vssd1 vccd1 vccd1 _06276_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14032_ clknet_leaf_83_clk _00801_ net1260 vssd1 vssd1 vccd1 vccd1 datapath.PC\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07528__X _02364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11244_ net304 net2467 net420 vssd1 vssd1 vccd1 vccd1 _00293_ sky130_fd_sc_hd__mux2_1
XANTENNA__10347__A1 net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11197__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11175_ net258 net2146 net425 vssd1 vssd1 vccd1 vccd1 _00227_ sky130_fd_sc_hd__mux2_1
XFILLER_121_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10126_ _04874_ _04876_ vssd1 vssd1 vccd1 vccd1 _04962_ sky130_fd_sc_hd__or2_1
XANTENNA__08960__A1 _02704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07407__C net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10057_ _04892_ _04829_ vssd1 vssd1 vccd1 vccd1 _04893_ sky130_fd_sc_hd__and2b_1
XANTENNA__07515__A2 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload0_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13816_ clknet_leaf_115_clk _00625_ net1189 vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__dfrtp_1
XFILLER_35_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08476__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13747_ clknet_leaf_88_clk _00556_ net1252 vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12756__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10959_ _05691_ _05696_ vssd1 vssd1 vccd1 vccd1 _05697_ sky130_fd_sc_hd__nor2_1
XFILLER_149_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13678_ clknet_leaf_1_clk _00488_ net1057 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_12629_ datapath.mulitply_result\[20\] datapath.multiplication_module.multiplicand_i\[20\]
+ vssd1 vssd1 vccd1 vccd1 _06471_ sky130_fd_sc_hd__nand2_1
XFILLER_31_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08228__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold105 mmio.memload_or_instruction\[13\] vssd1 vssd1 vccd1 vccd1 net1453 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12491__S net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold116 datapath.multiplication_module.multiplier_i\[15\] vssd1 vssd1 vccd1 vccd1
+ net1464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 mmio.key_data\[0\] vssd1 vssd1 vccd1 vccd1 net1475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 keypad.decode.sticky\[4\] vssd1 vssd1 vccd1 vccd1 net1486 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14299__RESET_B net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold149 net87 vssd1 vssd1 vccd1 vccd1 net1497 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07739__C1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout607 _03608_ vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__clkbuf_4
X_09840_ _03556_ _03561_ _03563_ vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__or3_1
Xfanout618 net619 vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout629 _03717_ vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__clkbuf_2
XFILLER_101_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09771_ _03947_ _03949_ _03978_ _04604_ vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__a211o_1
XANTENNA__07317__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06983_ net969 net908 _01800_ vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__and3_1
XFILLER_101_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08722_ _03127_ _03128_ vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__nand2b_2
X_08653_ _02025_ _02047_ vssd1 vssd1 vccd1 vccd1 _03489_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_1_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout172_A _05684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07604_ net610 _02438_ _01787_ vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__o21a_1
XANTENNA__13863__RESET_B net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08584_ net558 _03419_ vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_105_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07535_ datapath.rf.registers\[12\]\[20\] net754 net694 datapath.rf.registers\[8\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__a22o_1
XFILLER_34_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1081_A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1179_A net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07466_ datapath.rf.registers\[24\]\[21\] net856 net853 datapath.rf.registers\[19\]\[21\]
+ _02301_ vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__a221o_1
XANTENNA__06891__C net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09205_ net454 _03961_ _03962_ _04039_ net349 vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__a311oi_2
XANTENNA__08219__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07397_ datapath.rf.registers\[27\]\[23\] net683 net786 vssd1 vssd1 vccd1 vccd1 _02233_
+ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout225_X net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout604_A _04727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09136_ net338 _03693_ _03971_ vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_20_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09067_ _03705_ _03708_ net451 vssd1 vssd1 vccd1 vccd1 _03903_ sky130_fd_sc_hd__mux2_1
XANTENNA__12318__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08018_ _02830_ _02851_ _02852_ _02853_ vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__or4_1
XFILLER_151_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold650 datapath.rf.registers\[26\]\[17\] vssd1 vssd1 vccd1 vccd1 net1998 sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 datapath.rf.registers\[29\]\[24\] vssd1 vssd1 vccd1 vccd1 net2009 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout973_A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold672 datapath.rf.registers\[18\]\[12\] vssd1 vssd1 vccd1 vccd1 net2020 sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 datapath.rf.registers\[18\]\[23\] vssd1 vssd1 vccd1 vccd1 net2031 sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 datapath.rf.registers\[8\]\[21\] vssd1 vssd1 vccd1 vccd1 net2042 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07508__B net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07745__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08942__A1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09969_ _04748_ _04804_ vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout761_X net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout859_X net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12980_ net220 net2255 net478 vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__mux2_1
XFILLER_58_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11931_ net136 _05984_ _05983_ vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__o21ai_1
XFILLER_85_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08339__B net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10588__C _02145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14650_ clknet_leaf_136_clk _01355_ net1102 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11862_ net137 _05938_ _05937_ vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__o21ai_1
XFILLER_73_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08058__C net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13601_ clknet_leaf_46_clk _00411_ net1147 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10813_ net1266 _05565_ vssd1 vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12254__A1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14581_ clknet_leaf_16_clk _01286_ net1108 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11793_ _05899_ net336 vssd1 vssd1 vccd1 vccd1 _05905_ sky130_fd_sc_hd__nor2_1
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11480__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13532_ clknet_leaf_8_clk _00342_ net1074 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10744_ net1534 net568 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[30\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__07130__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13463_ clknet_leaf_126_clk _00273_ net1206 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10675_ _05444_ _05445_ _05450_ _05492_ vssd1 vssd1 vccd1 vccd1 _05493_ sky130_fd_sc_hd__a31o_1
XFILLER_139_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12414_ net1410 net131 _06354_ vssd1 vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__a21o_1
XFILLER_127_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13394_ clknet_leaf_30_clk _00204_ net1125 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_153_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12345_ net895 _06312_ _04928_ vssd1 vssd1 vccd1 vccd1 _06313_ sky130_fd_sc_hd__a21oi_1
XFILLER_127_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08802__B _03600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07984__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12276_ net892 _04836_ net190 vssd1 vssd1 vccd1 vccd1 _06263_ sky130_fd_sc_hd__a21o_1
XFILLER_141_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09186__A1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14015_ clknet_leaf_87_clk _00784_ net1252 vssd1 vssd1 vccd1 vccd1 datapath.PC\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_56_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11227_ net235 net2151 net528 vssd1 vssd1 vccd1 vccd1 _00277_ sky130_fd_sc_hd__mux2_1
XANTENNA__07197__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07736__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11158_ net241 net1998 net530 vssd1 vssd1 vccd1 vccd1 _00211_ sky130_fd_sc_hd__mux2_1
XFILLER_110_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10109_ datapath.PC\[19\] _04118_ net469 vssd1 vssd1 vccd1 vccd1 _04945_ sky130_fd_sc_hd__mux2_1
XANTENNA__12340__A net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11089_ net243 net2079 net535 vssd1 vssd1 vccd1 vccd1 _00146_ sky130_fd_sc_hd__mux2_1
XFILLER_64_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06976__C _01800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08161__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08964__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12486__S net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08449__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11390__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07320_ datapath.rf.registers\[13\]\[24\] net810 net804 datapath.rf.registers\[28\]\[24\]
+ _02155_ vssd1 vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__a221o_1
XFILLER_20_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07251_ datapath.rf.registers\[3\]\[26\] net770 net762 datapath.rf.registers\[1\]\[26\]
+ _02086_ vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__a221o_1
XFILLER_136_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07182_ datapath.rf.registers\[16\]\[27\] net861 net853 datapath.rf.registers\[19\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02018_ sky130_fd_sc_hd__a22o_1
XFILLER_129_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_Left_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13110__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08712__B _03358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07975__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire562_X net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08431__C _01825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout404 _06549_ vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__clkbuf_8
Xfanout415 _05726_ vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__buf_4
Xfanout426 _05716_ vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07727__A2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09823_ _01888_ _01909_ net625 vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__o21a_1
Xfanout437 _05697_ vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__clkbuf_4
Xfanout448 net451 vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__buf_2
Xfanout459 net462 vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__buf_2
XFILLER_140_381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout387_A net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09754_ net326 _04362_ _04363_ vssd1 vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_107_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12250__A _06168_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06966_ net964 net909 _01795_ vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__and3_2
XFILLER_39_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08705_ net560 _03079_ vssd1 vssd1 vccd1 vccd1 _03541_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_61_Left_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09685_ _04249_ _04432_ net353 vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__mux2_1
XFILLER_67_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06897_ net976 net928 vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_93_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_93_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_87_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_126_Right_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08636_ _01981_ _02003_ vssd1 vssd1 vccd1 vccd1 _03472_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_120_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07998__B net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08567_ datapath.rf.registers\[15\]\[0\] net968 _01825_ vssd1 vssd1 vccd1 vccd1 _03403_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10909__S net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09637__C1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout819_A net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1084_X net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07518_ datapath.rf.registers\[12\]\[20\] net826 net794 datapath.rf.registers\[31\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _02354_ sky130_fd_sc_hd__a22o_1
XANTENNA__07112__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08498_ datapath.rf.registers\[15\]\[1\] net970 _01825_ vssd1 vssd1 vccd1 vccd1 _03334_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12409__B net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07510__C net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07449_ net563 _02284_ vssd1 vssd1 vccd1 vccd1 _02285_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout1251_X net1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout607_X net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10460_ keypad.decode.sticky\[3\] keypad.decode.sticky\[2\] net1022 vssd1 vssd1 vccd1
+ vccd1 keypad.decode.sticky_n\[2\] sky130_fd_sc_hd__mux2_1
XFILLER_6_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_70_Left_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09119_ _02169_ _02217_ net442 vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__mux2_1
XFILLER_108_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10391_ _03263_ _03657_ _04346_ net458 vssd1 vssd1 vccd1 vccd1 _05227_ sky130_fd_sc_hd__o211ai_1
XANTENNA__13020__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12130_ screen.counter.ct\[21\] screen.counter.ct\[22\] _06166_ vssd1 vssd1 vccd1
+ vccd1 _06167_ sky130_fd_sc_hd__and3_2
XFILLER_2_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout976_X net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08341__C net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10970__B2 _01443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12061_ net1011 _06099_ _06101_ net1001 vssd1 vssd1 vccd1 vccd1 _06102_ sky130_fd_sc_hd__a22o_1
Xhold480 datapath.rf.registers\[30\]\[27\] vssd1 vssd1 vccd1 vccd1 net1828 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07179__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold491 datapath.rf.registers\[22\]\[11\] vssd1 vssd1 vccd1 vccd1 net1839 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07718__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11012_ net279 net1920 net540 vssd1 vssd1 vccd1 vccd1 _00074_ sky130_fd_sc_hd__mux2_1
XFILLER_78_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06926__B1 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10722__A1 _02960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11475__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout960 _01708_ vssd1 vssd1 vccd1 vccd1 net960 sky130_fd_sc_hd__buf_4
Xfanout971 _01675_ vssd1 vssd1 vccd1 vccd1 net971 sky130_fd_sc_hd__clkbuf_4
XFILLER_49_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout982 net983 vssd1 vssd1 vccd1 vccd1 net982 sky130_fd_sc_hd__clkbuf_2
XFILLER_92_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout993 _01567_ vssd1 vssd1 vccd1 vccd1 net993 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_51_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12963_ net258 net1555 net481 vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_84_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_clk sky130_fd_sc_hd__clkbuf_8
Xhold1180 datapath.rf.registers\[17\]\[26\] vssd1 vssd1 vccd1 vccd1 net2528 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09340__A1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1191 datapath.mulitply_result\[7\] vssd1 vssd1 vccd1 vccd1 net2539 sky130_fd_sc_hd__dlygate4sd3_1
X_11914_ screen.register.currentYbus\[19\] net162 vssd1 vssd1 vccd1 vccd1 _05973_
+ sky130_fd_sc_hd__nand2_1
X_12894_ net170 net2315 net399 vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__mux2_1
XANTENNA__07351__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14633_ clknet_leaf_62_clk _01338_ net1165 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11845_ _05358_ _05913_ _05919_ _05335_ _05923_ vssd1 vssd1 vccd1 vccd1 _05924_ sky130_fd_sc_hd__a221o_1
XFILLER_61_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14564_ clknet_leaf_22_clk _01269_ net1157 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11776_ columns.count\[5\] columns.count\[4\] _05893_ vssd1 vssd1 vccd1 vccd1 _05894_
+ sky130_fd_sc_hd__nor3_4
XANTENNA__07103__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12319__B _04600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13515_ clknet_leaf_57_clk _00325_ net1161 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_109_Left_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10727_ net2642 _02704_ _05367_ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[13\]
+ sky130_fd_sc_hd__mux2_1
X_14495_ clknet_leaf_12_clk _01200_ net1080 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_13446_ clknet_leaf_23_clk _00256_ net1154 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10658_ _05473_ _05476_ _05462_ vssd1 vssd1 vccd1 vccd1 _05477_ sky130_fd_sc_hd__o21a_1
Xclkload14 clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clkload14/Y sky130_fd_sc_hd__inv_6
Xclkload25 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 clkload25/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_58_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload36 clknet_leaf_138_clk vssd1 vssd1 vccd1 vccd1 clkload36/Y sky130_fd_sc_hd__bufinv_16
Xclkload47 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 clkload47/Y sky130_fd_sc_hd__clkinvlp_4
X_13377_ clknet_leaf_46_clk _00187_ net1171 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10589_ _01855_ _01908_ _01954_ _02002_ vssd1 vssd1 vccd1 vccd1 _05412_ sky130_fd_sc_hd__or4_1
Xclkload58 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 clkload58/Y sky130_fd_sc_hd__clkinv_8
Xclkload69 clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 clkload69/Y sky130_fd_sc_hd__inv_6
XANTENNA__10410__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07957__A2 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12328_ net894 _04084_ _06299_ _06300_ vssd1 vssd1 vccd1 vccd1 _06301_ sky130_fd_sc_hd__o22a_1
XFILLER_5_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12259_ _05205_ net308 _06249_ _06248_ vssd1 vssd1 vccd1 vccd1 _00781_ sky130_fd_sc_hd__o31a_1
XFILLER_141_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_118_Left_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10713__A1 _03262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06987__B _01637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11385__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08382__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06820_ net1002 net1018 _01654_ net1026 datapath.ru.latched_instruction\[16\] vssd1
+ vssd1 vccd1 vccd1 _01656_ sky130_fd_sc_hd__a32o_4
XANTENNA__13166__A datapath.rf.registers\[0\]\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07590__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06751_ _01576_ _01589_ vssd1 vssd1 vccd1 vccd1 MemWrite sky130_fd_sc_hd__nor2_2
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_75_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_92_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08134__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06682_ datapath.ru.latched_instruction\[18\] _01454_ _01498_ datapath.ru.latched_instruction\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__a22o_1
X_09470_ net552 net548 _02912_ vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__a21o_1
XFILLER_63_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08421_ datapath.rf.registers\[11\]\[2\] net884 net843 datapath.rf.registers\[25\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_102_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10729__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13105__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08352_ datapath.rf.registers\[31\]\[3\] net978 net916 vssd1 vssd1 vccd1 vccd1 _03188_
+ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_127_Left_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07303_ datapath.rf.registers\[17\]\[25\] net748 net724 datapath.rf.registers\[18\]\[25\]
+ _02138_ vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__a221o_2
XANTENNA__08842__A0 _03358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08283_ datapath.rf.registers\[26\]\[5\] net779 net727 datapath.rf.registers\[25\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03119_ sky130_fd_sc_hd__a22o_1
XANTENNA__12944__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout135_A _05934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload8 clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clkload8/Y sky130_fd_sc_hd__inv_6
X_07234_ _02069_ vssd1 vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__inv_2
X_07165_ _01986_ _02000_ _01415_ net788 vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__a2bb2o_4
XANTENNA_fanout1044_A _03729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07096_ _01913_ _01915_ _01930_ _01931_ vssd1 vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__or4_1
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_136_Left_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1211_A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout201 net202 vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__clkbuf_2
XFILLER_120_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout212 net213 vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__clkbuf_2
Xfanout223 _04713_ vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout671_A net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10704__A1 _02934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout234 _05623_ vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__buf_1
Xfanout245 net246 vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11295__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout256 net257 vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__buf_1
XANTENNA__06897__B net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09806_ net322 _04638_ _04641_ vssd1 vssd1 vccd1 vccd1 _04642_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_89_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout267 net269 vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__08373__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout278 _05554_ vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__clkbuf_2
XFILLER_28_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07998_ datapath.rf.registers\[6\]\[10\] net952 net935 vssd1 vssd1 vccd1 vccd1 _02834_
+ sky130_fd_sc_hd__and3_1
Xfanout289 _05706_ vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__buf_1
XANTENNA__07074__A _01889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09737_ net377 _04066_ _04572_ vssd1 vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__o21a_1
X_06949_ _01593_ _01784_ vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__nor2_1
XFILLER_55_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout936_A _01725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09322__A1 _02467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_66_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_28_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09668_ net371 _04406_ _04503_ vssd1 vssd1 vccd1 vccd1 _04504_ sky130_fd_sc_hd__a21o_1
XFILLER_91_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08619_ _02311_ _02332_ vssd1 vssd1 vccd1 vccd1 _03455_ sky130_fd_sc_hd__or2_1
X_09599_ net349 _04434_ _04433_ net359 vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__o211a_1
XFILLER_91_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout724_X net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13015__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11630_ _05787_ _05853_ vssd1 vssd1 vccd1 vccd1 _05854_ sky130_fd_sc_hd__nor2_1
XFILLER_42_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10585__D _03170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11561_ _05293_ _05774_ vssd1 vssd1 vccd1 vccd1 _05785_ sky130_fd_sc_hd__or2_2
XANTENNA__12854__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13300_ clknet_leaf_94_clk _00110_ net1211 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10512_ net1280 net1275 net1271 vssd1 vssd1 vccd1 vccd1 _05342_ sky130_fd_sc_hd__nor3_1
XANTENNA__08192__X _03028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14280_ clknet_leaf_64_clk _00985_ net1236 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_11492_ net251 net2439 net510 vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__mux2_1
XFILLER_155_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_133_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13231_ clknet_leaf_30_clk _00041_ net1132 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10443_ _04837_ _04838_ net227 vssd1 vssd1 vccd1 vccd1 _05279_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_150_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13162_ net286 net2136 net544 vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__mux2_1
X_10374_ net222 _04837_ net1292 vssd1 vssd1 vccd1 vccd1 _05210_ sky130_fd_sc_hd__a21oi_1
XFILLER_156_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12113_ screen.counter.currentCt\[21\] screen.counter.currentCt\[20\] screen.counter.currentCt\[22\]
+ _06149_ vssd1 vssd1 vccd1 vccd1 _06150_ sky130_fd_sc_hd__or4_1
X_13093_ net1799 net170 net387 vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12044_ _05782_ _06083_ _06085_ net1011 vssd1 vssd1 vccd1 vccd1 _06086_ sky130_fd_sc_hd__o31a_1
XFILLER_78_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08364__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07255__Y _02091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06600__B _01438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout790 net792 vssd1 vssd1 vccd1 vccd1 net790 sky130_fd_sc_hd__clkbuf_8
XFILLER_93_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13995_ clknet_leaf_112_clk _00772_ net1197 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_57_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_74_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08116__A2 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12946_ net240 net2145 net396 vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__mux2_1
XANTENNA__07324__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08367__X _03203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08808__A net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06678__A2 _01467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12877_ net251 net2284 net399 vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__mux2_1
XANTENNA__08527__B net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14616_ clknet_leaf_6_clk _01321_ net1067 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11828_ net1278 net1279 vssd1 vssd1 vccd1 vccd1 _05907_ sky130_fd_sc_hd__and2_1
XFILLER_61_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14547_ clknet_leaf_34_clk _01252_ net1128 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11759_ net1463 net146 net141 _02439_ vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__a22o_1
XANTENNA__12764__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11888__B net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14478_ clknet_leaf_1_clk _01183_ net1063 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload103 clknet_leaf_123_clk vssd1 vssd1 vccd1 vccd1 clkload103/Y sky130_fd_sc_hd__clkinv_8
Xclkload114 clknet_leaf_109_clk vssd1 vssd1 vccd1 vccd1 clkload114/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__11240__Y _05722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13429_ clknet_leaf_19_clk _00239_ net1116 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload125 clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 clkload125/Y sky130_fd_sc_hd__inv_6
XANTENNA__06850__A2 _01595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload136 clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 clkload136/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload147 clknet_leaf_83_clk vssd1 vssd1 vccd1 vccd1 clkload147/Y sky130_fd_sc_hd__inv_6
XFILLER_142_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08970_ _03803_ _03805_ net448 vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__mux2_1
XANTENNA__06998__A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07921_ datapath.rf.registers\[1\]\[12\] net763 net692 datapath.rf.registers\[13\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__a22o_1
XANTENNA__10147__C1 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08355__A2 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07852_ datapath.rf.registers\[14\]\[13\] net829 net794 datapath.rf.registers\[31\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__a22o_1
X_06803_ _01453_ net1003 net1019 net1026 datapath.ru.latched_instruction\[18\] vssd1
+ vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__a32o_4
Xinput1 ACK_I vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_1
X_07783_ datapath.rf.registers\[12\]\[15\] net755 net684 datapath.rf.registers\[27\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02619_ sky130_fd_sc_hd__a22o_1
XANTENNA__12939__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_48_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_65_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08107__A2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09522_ net354 net458 _03772_ vssd1 vssd1 vccd1 vccd1 _04358_ sky130_fd_sc_hd__or3_1
X_06734_ _01441_ net1005 _01566_ datapath.ru.latched_instruction\[5\] vssd1 vssd1
+ vccd1 vccd1 _01573_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_84_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06669__A2 _01502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09453_ _02751_ _02805_ net442 vssd1 vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__mux2_1
XFILLER_80_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06665_ net1288 net1283 mmio.memload_or_instruction\[26\] vssd1 vssd1 vccd1 vccd1
+ _01504_ sky130_fd_sc_hd__or3b_1
XFILLER_25_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout252_A _05588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08437__B _01797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08404_ datapath.rf.registers\[6\]\[2\] net953 net936 vssd1 vssd1 vccd1 vccd1 _03240_
+ sky130_fd_sc_hd__and3_1
X_09384_ net357 net352 net458 _03772_ vssd1 vssd1 vccd1 vccd1 _04220_ sky130_fd_sc_hd__or4_2
X_06596_ net34 net39 vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__nand2_2
XANTENNA__08815__A0 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08335_ _03150_ _03170_ net613 vssd1 vssd1 vccd1 vccd1 _03171_ sky130_fd_sc_hd__mux2_2
XANTENNA_fanout1161_A net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout517_A _05731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07094__A2 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08266_ _03094_ _03097_ _03098_ _03101_ vssd1 vssd1 vccd1 vccd1 _03102_ sky130_fd_sc_hd__or4_1
XANTENNA__07995__C net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07217_ datapath.rf.registers\[24\]\[26\] net856 net845 datapath.rf.registers\[1\]\[26\]
+ _02052_ vssd1 vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_115_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08197_ _03009_ _03030_ vssd1 vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_144_Left_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08043__A1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07148_ datapath.rf.registers\[2\]\[28\] net744 net685 datapath.rf.registers\[27\]\[28\]
+ _01983_ vssd1 vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__a221o_1
XFILLER_145_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout886_A _01716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10922__S net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07079_ datapath.rf.registers\[11\]\[29\] net883 net836 datapath.rf.registers\[26\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01915_ sky130_fd_sc_hd__a22o_1
XFILLER_105_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10090_ _04921_ _04922_ _04924_ _04925_ net895 vssd1 vssd1 vccd1 vccd1 _04926_ sky130_fd_sc_hd__o221a_1
Xfanout1007 _05756_ vssd1 vssd1 vccd1 vccd1 net1007 sky130_fd_sc_hd__clkbuf_2
Xfanout1018 net1020 vssd1 vssd1 vccd1 vccd1 net1018 sky130_fd_sc_hd__buf_4
XFILLER_102_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1029 net1032 vssd1 vssd1 vccd1 vccd1 net1029 sky130_fd_sc_hd__buf_4
XANTENNA_fanout674_X net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout841_X net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12849__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout939_X net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_39_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_8
X_12800_ net1693 net302 net492 vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_153_Left_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13780_ clknet_leaf_51_clk _00589_ net1181 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10992_ net1610 net203 net435 vssd1 vssd1 vccd1 vccd1 _00057_ sky130_fd_sc_hd__mux2_1
XANTENNA__07306__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08628__A _02170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12731_ net1548 net208 net405 vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__mux2_1
XFILLER_16_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08347__B net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12662_ datapath.mulitply_result\[25\] datapath.multiplication_module.multiplicand_i\[25\]
+ vssd1 vssd1 vccd1 vccd1 _06499_ sky130_fd_sc_hd__nor2_1
X_14401_ clknet_leaf_56_clk _01106_ net1158 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14165__RESET_B net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11613_ net1006 _05762_ vssd1 vssd1 vccd1 vccd1 _05837_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_46_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12593_ datapath.mulitply_result\[14\] datapath.multiplication_module.multiplicand_i\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06441_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_13_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14332_ clknet_leaf_7_clk _01037_ net1071 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11544_ _05292_ net1009 _05763_ vssd1 vssd1 vccd1 vccd1 _05768_ sky130_fd_sc_hd__nor3_4
XANTENNA__07085__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire465 _02238_ vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__buf_4
X_14263_ clknet_leaf_127_clk _00968_ net1210 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11475_ net2362 net168 net406 vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__mux2_1
XFILLER_137_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13214_ clknet_leaf_150_clk _00024_ net1059 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_143_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10426_ net381 _04127_ _05261_ _03614_ vssd1 vssd1 vccd1 vccd1 _05262_ sky130_fd_sc_hd__a211oi_2
X_14194_ clknet_leaf_67_clk datapath.multiplication_module.multiplicand_i_n\[5\] net1239
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08585__A2 _03358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13145_ net2540 net239 net384 vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__mux2_1
X_10357_ _03736_ _05192_ net1039 vssd1 vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__a21oi_1
XFILLER_152_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13076_ net2203 net253 net387 vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__mux2_1
X_10288_ _04846_ _05123_ vssd1 vssd1 vccd1 vccd1 _05124_ sky130_fd_sc_hd__nand2_1
XANTENNA__09534__A1 _02751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12027_ _05759_ _05851_ _05854_ _05846_ vssd1 vssd1 vccd1 vccd1 _06070_ sky130_fd_sc_hd__a211o_1
XFILLER_38_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07545__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12759__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13978_ clknet_leaf_107_clk _00756_ net1223 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[21\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08097__X _02933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06984__C net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12929_ net208 net1657 net397 vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__mux2_1
XFILLER_33_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08825__X _03661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12494__S net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08120_ _02940_ _02953_ _02954_ _02955_ vssd1 vssd1 vccd1 vccd1 _02956_ sky130_fd_sc_hd__or4_1
XANTENNA__09470__B1 _02912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08051_ datapath.rf.registers\[22\]\[9\] net952 net924 vssd1 vssd1 vccd1 vccd1 _02887_
+ sky130_fd_sc_hd__and3_1
XFILLER_116_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12357__B1 _06253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07002_ datapath.rf.registers\[23\]\[31\] net698 net687 datapath.rf.registers\[31\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__a22o_1
XFILLER_131_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10383__A2 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07784__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08953_ _02365_ _02419_ net445 vssd1 vssd1 vccd1 vccd1 _03789_ sky130_fd_sc_hd__mux2_1
XANTENNA__08328__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07904_ net875 _02737_ _02738_ _02739_ vssd1 vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__or4_1
X_08884_ _01613_ _01618_ vssd1 vssd1 vccd1 vccd1 _03720_ sky130_fd_sc_hd__nor2_1
XANTENNA__07536__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07000__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07835_ datapath.rf.registers\[12\]\[14\] net755 net680 datapath.rf.registers\[6\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02671_ sky130_fd_sc_hd__a22o_1
XFILLER_110_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout467_A _01701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07766_ datapath.rf.registers\[18\]\[15\] net792 _02592_ _02600_ _02601_ vssd1 vssd1
+ vccd1 vccd1 _02602_ sky130_fd_sc_hd__a2111o_1
XFILLER_65_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09505_ _03009_ net552 net548 vssd1 vssd1 vccd1 vccd1 _04341_ sky130_fd_sc_hd__and3_1
X_06717_ mmio.memload_or_instruction\[19\] mmio.memload_or_instruction\[21\] mmio.memload_or_instruction\[22\]
+ mmio.memload_or_instruction\[20\] vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__or4bb_1
XFILLER_25_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout634_A net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07697_ datapath.rf.registers\[10\]\[17\] net708 net673 datapath.rf.registers\[7\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__a22o_1
XFILLER_25_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08500__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09436_ net631 _04241_ _04243_ _04271_ vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__a22o_2
X_06648_ datapath.ru.latched_instruction\[4\] _01449_ _01485_ datapath.ru.latched_instruction\[6\]
+ _01483_ vssd1 vssd1 vccd1 vccd1 _01487_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout801_A net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09367_ _03520_ net626 net625 _03521_ net643 vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout422_X net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06579_ screen.register.xFill2 vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__inv_2
XFILLER_138_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11602__A _05773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08318_ datapath.rf.registers\[14\]\[4\] net774 net742 datapath.rf.registers\[2\]\[4\]
+ _03151_ vssd1 vssd1 vccd1 vccd1 _03154_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_10_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07067__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09298_ _04040_ _04133_ net353 vssd1 vssd1 vccd1 vccd1 _04134_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08249_ datapath.rf.registers\[28\]\[5\] net805 net796 datapath.rf.registers\[29\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03085_ sky130_fd_sc_hd__a22o_1
XFILLER_21_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11260_ net237 net2450 net420 vssd1 vssd1 vccd1 vccd1 _00309_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout791_X net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout889_X net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10211_ _04601_ _05046_ _05045_ net230 vssd1 vssd1 vccd1 vccd1 _05047_ sky130_fd_sc_hd__o211a_1
X_11191_ net239 net2555 net424 vssd1 vssd1 vccd1 vccd1 _00243_ sky130_fd_sc_hd__mux2_1
X_10142_ _04611_ _04623_ _01702_ _04609_ vssd1 vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__a211o_1
XANTENNA__08319__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10073_ datapath.PC\[31\] net1292 _04716_ _04908_ vssd1 vssd1 vccd1 vccd1 _04909_
+ sky130_fd_sc_hd__a22o_2
XFILLER_48_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_128_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13901_ clknet_leaf_43_clk net1360 net1150 vssd1 vssd1 vccd1 vccd1 keypad.debounce.debounce\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input28_A DAT_I[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10888__A net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11483__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13832_ clknet_leaf_113_clk _00641_ net1195 vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__dfrtp_1
XFILLER_47_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13763_ clknet_leaf_81_clk _00572_ net1255 vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10975_ net1923 net290 net435 vssd1 vssd1 vccd1 vccd1 _00040_ sky130_fd_sc_hd__mux2_1
XFILLER_71_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12714_ columns.count\[0\] columns.count\[5\] columns.count\[4\] _01433_ vssd1 vssd1
+ vccd1 vccd1 _06538_ sky130_fd_sc_hd__and4_1
XFILLER_16_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13694_ clknet_leaf_150_clk _00504_ net1059 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_12645_ _06477_ _06483_ _06482_ _06481_ vssd1 vssd1 vccd1 vccd1 _06485_ sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_61_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07058__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12576_ datapath.mulitply_result\[11\] datapath.multiplication_module.multiplicand_i\[11\]
+ vssd1 vssd1 vccd1 vccd1 _06427_ sky130_fd_sc_hd__nor2_1
XANTENNA__12327__B _06254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14315_ clknet_leaf_56_clk _01020_ net1173 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11527_ _05749_ _05750_ vssd1 vssd1 vccd1 vccd1 _05751_ sky130_fd_sc_hd__or2_2
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14246_ clknet_leaf_124_clk datapath.multiplication_module.multiplier_i_n\[14\] net1215
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i\[14\] sky130_fd_sc_hd__dfrtp_1
Xhold309 datapath.rf.registers\[3\]\[0\] vssd1 vssd1 vccd1 vccd1 net1657 sky130_fd_sc_hd__dlygate4sd3_1
X_11458_ net2599 _05588_ net407 vssd1 vssd1 vccd1 vccd1 _00496_ sky130_fd_sc_hd__mux2_1
XANTENNA__09755__A1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10409_ net607 _05243_ _05244_ _03604_ net555 vssd1 vssd1 vccd1 vccd1 _05245_ sky130_fd_sc_hd__o221a_1
X_14177_ clknet_leaf_48_clk _00932_ net1177 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11389_ net1936 net265 net411 vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__mux2_1
XFILLER_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08963__C1 _03673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13128_ net2166 net207 net384 vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__mux2_1
XANTENNA__07230__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13059_ net174 net2088 net476 vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__mux2_1
XFILLER_23_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08967__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1009 datapath.rf.registers\[16\]\[1\] vssd1 vssd1 vccd1 vccd1 net2357 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07518__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12511__B1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12489__S net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11393__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06995__B _01637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07620_ datapath.rf.registers\[16\]\[18\] net860 net826 datapath.rf.registers\[12\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07551_ _02365_ _02386_ vssd1 vssd1 vccd1 vccd1 _02387_ sky130_fd_sc_hd__nor2_1
XANTENNA__14016__RESET_B net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07482_ datapath.rf.registers\[19\]\[21\] net730 net683 datapath.rf.registers\[27\]\[21\]
+ _02316_ vssd1 vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__a221o_1
XANTENNA__07297__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09221_ _01706_ _04025_ _04056_ net605 vssd1 vssd1 vccd1 vccd1 _04057_ sky130_fd_sc_hd__o22ai_4
XANTENNA__13113__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09152_ _03985_ _03987_ net375 vssd1 vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__mux2_1
XANTENNA__07049__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12042__A2 _05786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09443__B1 _02804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08103_ datapath.rf.registers\[11\]\[8\] net883 net806 datapath.rf.registers\[28\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__a22o_1
XANTENNA__12952__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09083_ _02025_ _02069_ net442 vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08034_ datapath.rf.registers\[12\]\[10\] net756 net700 datapath.rf.registers\[23\]\[10\]
+ _02867_ vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__a221o_1
XANTENNA__06803__X _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold810 datapath.rf.registers\[24\]\[26\] vssd1 vssd1 vccd1 vccd1 net2158 sky130_fd_sc_hd__dlygate4sd3_1
Xhold821 datapath.rf.registers\[20\]\[15\] vssd1 vssd1 vccd1 vccd1 net2169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold832 datapath.rf.registers\[28\]\[28\] vssd1 vssd1 vccd1 vccd1 net2180 sky130_fd_sc_hd__dlygate4sd3_1
Xhold843 datapath.rf.registers\[21\]\[7\] vssd1 vssd1 vccd1 vccd1 net2191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold854 datapath.rf.registers\[5\]\[22\] vssd1 vssd1 vccd1 vccd1 net2202 sky130_fd_sc_hd__dlygate4sd3_1
Xhold865 datapath.rf.registers\[12\]\[25\] vssd1 vssd1 vccd1 vccd1 net2213 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold876 datapath.rf.registers\[24\]\[17\] vssd1 vssd1 vccd1 vccd1 net2224 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold887 datapath.rf.registers\[10\]\[4\] vssd1 vssd1 vccd1 vccd1 net2235 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06889__C net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_51_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07221__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold898 datapath.rf.registers\[24\]\[20\] vssd1 vssd1 vccd1 vccd1 net2246 sky130_fd_sc_hd__dlygate4sd3_1
X_09985_ _04722_ _04820_ vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__and2b_1
XFILLER_89_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08936_ net566 _01889_ net453 vssd1 vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__mux2_1
X_08867_ _03701_ _03702_ net449 vssd1 vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout751_A _01804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08182__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout849_A _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_66_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07818_ datapath.rf.registers\[2\]\[14\] net888 net837 datapath.rf.registers\[26\]\[14\]
+ _02653_ vssd1 vssd1 vccd1 vccd1 _02654_ sky130_fd_sc_hd__a221o_1
XFILLER_85_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08798_ net328 _03633_ _03623_ vssd1 vssd1 vccd1 vccd1 _03634_ sky130_fd_sc_hd__o21a_1
X_07749_ datapath.rf.registers\[4\]\[16\] net714 net671 datapath.rf.registers\[7\]\[16\]
+ _02583_ vssd1 vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_123_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07513__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10760_ _05524_ _05525_ vssd1 vssd1 vccd1 vccd1 _05526_ sky130_fd_sc_hd__nor2_1
XANTENNA__12281__A2 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09419_ net648 _04254_ net438 vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__a21oi_1
X_10691_ button\[4\] net1022 _05458_ _05465_ vssd1 vssd1 vccd1 vccd1 _05507_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout804_X net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_124_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13023__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12430_ net1429 net131 _06362_ vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_101_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08344__C net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12361_ net637 _04645_ net309 vssd1 vssd1 vccd1 vccd1 _06325_ sky130_fd_sc_hd__a21o_1
XFILLER_148_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14100_ clknet_leaf_111_clk _00866_ net1198 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_126_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11312_ net2456 net304 net416 vssd1 vssd1 vccd1 vccd1 _00357_ sky130_fd_sc_hd__mux2_1
XFILLER_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12292_ net634 _04835_ vssd1 vssd1 vccd1 vccd1 _06275_ sky130_fd_sc_hd__nor2_1
XANTENNA__07460__A2 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_139_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14031_ clknet_leaf_83_clk _00800_ net1260 vssd1 vssd1 vccd1 vccd1 datapath.PC\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_4_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13321__RESET_B net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11478__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11243_ net289 net2361 net421 vssd1 vssd1 vccd1 vccd1 _00292_ sky130_fd_sc_hd__mux2_1
XFILLER_4_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07748__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_19_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11174_ net207 net2018 net425 vssd1 vssd1 vccd1 vccd1 _00226_ sky130_fd_sc_hd__mux2_1
X_10125_ _04603_ _04960_ _04959_ _04957_ net226 vssd1 vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__a2111o_1
XFILLER_95_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10056_ _04885_ _04888_ _04891_ vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__or3b_1
XFILLER_76_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13815_ clknet_leaf_115_clk _00624_ net1187 vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_34_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13746_ clknet_leaf_76_clk net1291 net1247 vssd1 vssd1 vccd1 vccd1 mmio.wishbone.prev_BUSY_O
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07279__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10958_ _05693_ _05694_ vssd1 vssd1 vccd1 vccd1 _05696_ sky130_fd_sc_hd__or2_4
X_13677_ clknet_leaf_123_clk _00487_ net1207 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10889_ datapath.PC\[23\] _05629_ vssd1 vssd1 vccd1 vccd1 _05636_ sky130_fd_sc_hd__and2_1
XFILLER_148_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12628_ net498 _06469_ _06470_ net502 net2615 vssd1 vssd1 vccd1 vccd1 _00929_ sky130_fd_sc_hd__a32o_1
XANTENNA__09274__A1_N _03667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12772__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12559_ _06410_ _06411_ _06412_ vssd1 vssd1 vccd1 vccd1 _06413_ sky130_fd_sc_hd__or3_1
XFILLER_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold106 mmio.key_data\[3\] vssd1 vssd1 vccd1 vccd1 net1454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold117 datapath.multiplication_module.multiplier_i\[13\] vssd1 vssd1 vccd1 vccd1
+ net1465 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold128 net92 vssd1 vssd1 vccd1 vccd1 net1476 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11388__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14229_ clknet_leaf_42_clk _00950_ net1144 vssd1 vssd1 vccd1 vccd1 columns.count\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold139 keypad.decode.sticky_n\[4\] vssd1 vssd1 vccd1 vccd1 net1487 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_153_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_74_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07203__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout608 _03608_ vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__clkbuf_2
Xfanout619 MemRead vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__buf_2
XFILLER_98_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_107_Right_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09770_ _03947_ _03949_ _03978_ _04604_ vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__a211oi_1
X_06982_ net968 net909 net908 vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__and3_1
XFILLER_86_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11299__A0 _05653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08721_ _03555_ _03556_ _03543_ vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__a21o_1
XFILLER_94_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1190 net1204 vssd1 vssd1 vccd1 vccd1 net1190 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13108__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08652_ _02025_ _02047_ vssd1 vssd1 vccd1 vccd1 _03488_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_1_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07911__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07603_ _02438_ vssd1 vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_1_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08583_ net612 _03417_ _03384_ vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__a21o_2
XFILLER_82_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12947__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout165_A _05288_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07534_ datapath.rf.registers\[19\]\[20\] net732 net687 datapath.rf.registers\[31\]\[20\]
+ _02366_ vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__a221o_1
X_07465_ datapath.rf.registers\[13\]\[21\] net810 net807 datapath.rf.registers\[27\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1074_A net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09204_ net454 _03961_ _03962_ _04039_ vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__a31oi_1
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07396_ datapath.rf.registers\[17\]\[23\] net746 net694 datapath.rf.registers\[8\]\[23\]
+ _02231_ vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__a221o_1
XANTENNA__07690__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09135_ net321 _03707_ net323 vssd1 vssd1 vccd1 vccd1 _03971_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_20_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1241_A net1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07978__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09557__A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09066_ net338 _03901_ _03900_ net322 vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__a211o_1
XFILLER_136_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07442__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11298__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout799_A net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08017_ datapath.rf.registers\[10\]\[10\] net881 net838 datapath.rf.registers\[26\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__a22o_1
Xhold640 datapath.rf.registers\[25\]\[7\] vssd1 vssd1 vccd1 vccd1 net1988 sky130_fd_sc_hd__dlygate4sd3_1
Xhold651 datapath.rf.registers\[17\]\[25\] vssd1 vssd1 vccd1 vccd1 net1999 sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 datapath.rf.registers\[0\]\[18\] vssd1 vssd1 vccd1 vccd1 net2010 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold673 datapath.rf.registers\[0\]\[21\] vssd1 vssd1 vccd1 vccd1 net2021 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold684 datapath.rf.registers\[9\]\[12\] vssd1 vssd1 vccd1 vccd1 net2032 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold695 datapath.rf.registers\[13\]\[31\] vssd1 vssd1 vccd1 vccd1 net2043 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout966_A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09968_ _04753_ _04757_ _04801_ _04752_ _04750_ vssd1 vssd1 vccd1 vccd1 _04804_ sky130_fd_sc_hd__a311o_1
XFILLER_77_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08919_ _03732_ _03754_ net637 vssd1 vssd1 vccd1 vccd1 _03755_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_125_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09899_ datapath.PC\[17\] _04727_ _04734_ vssd1 vssd1 vccd1 vccd1 _04735_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout754_X net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08155__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13018__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11930_ _02189_ net658 vssd1 vssd1 vccd1 vccd1 _05984_ sky130_fd_sc_hd__nand2_1
XFILLER_58_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07902__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10588__D _02189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08339__C net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11861_ _03357_ net658 vssd1 vssd1 vccd1 vccd1 _05938_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout921_X net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12857__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13600_ clknet_leaf_136_clk _00410_ net1090 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10812_ net269 net2040 net543 vssd1 vssd1 vccd1 vccd1 _00013_ sky130_fd_sc_hd__mux2_1
X_14580_ clknet_leaf_128_clk _01285_ net1117 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11792_ datapath.ru.ack_mul_reg _05898_ _05899_ _05903_ _05902_ vssd1 vssd1 vccd1
+ vccd1 _05904_ sky130_fd_sc_hd__o221ai_4
XANTENNA__08636__A _01981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10265__A1 _04272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13531_ clknet_leaf_36_clk _00341_ net1136 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10743_ net1521 net569 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[29\]
+ sky130_fd_sc_hd__and2_1
XFILLER_43_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13462_ clknet_leaf_141_clk _00272_ net1096 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10674_ _05429_ _05491_ vssd1 vssd1 vccd1 vccd1 _05492_ sky130_fd_sc_hd__nor2_1
XANTENNA__07681__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12413_ _05970_ net158 vssd1 vssd1 vccd1 vccd1 _06354_ sky130_fd_sc_hd__nor2_1
X_13393_ clknet_leaf_41_clk _00203_ net1141 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07969__B1 _02803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11765__B2 _02145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12344_ _04884_ _05649_ net230 vssd1 vssd1 vccd1 vccd1 _06312_ sky130_fd_sc_hd__mux2_1
XFILLER_138_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07433__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12275_ net639 _04474_ vssd1 vssd1 vccd1 vccd1 _06262_ sky130_fd_sc_hd__nand2_1
XFILLER_154_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10406__A net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14014_ clknet_leaf_87_clk _00783_ net1252 vssd1 vssd1 vccd1 vccd1 datapath.PC\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_11226_ net219 net2297 net526 vssd1 vssd1 vccd1 vccd1 _00276_ sky130_fd_sc_hd__mux2_1
XFILLER_141_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10851__B1_N _05603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11157_ net246 net1787 net530 vssd1 vssd1 vccd1 vccd1 _00210_ sky130_fd_sc_hd__mux2_1
XFILLER_49_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10108_ _04933_ _04943_ vssd1 vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__nand2_1
X_11088_ net247 net2374 net534 vssd1 vssd1 vccd1 vccd1 _00145_ sky130_fd_sc_hd__mux2_1
XFILLER_49_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10039_ datapath.PC\[20\] net596 _04814_ vssd1 vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__a21oi_1
XFILLER_49_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12767__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07450__A net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13729_ clknet_leaf_25_clk _00539_ net1137 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_07250_ datapath.rf.registers\[7\]\[26\] net671 net664 datapath.rf.registers\[15\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__a22o_1
XFILLER_20_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07672__A2 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08833__X _03669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07181_ datapath.rf.registers\[3\]\[27\] net801 net793 datapath.rf.registers\[31\]\[27\]
+ _02006_ vssd1 vssd1 vccd1 vccd1 _02017_ sky130_fd_sc_hd__a221o_1
XANTENNA__11756__B2 _02587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07424__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07609__B net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout405 _06549_ vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08385__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout416 net417 vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_6_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout427 _05716_ vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__buf_4
X_09822_ net321 _04007_ _04657_ net322 vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__a211oi_1
Xfanout438 net439 vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__buf_2
XFILLER_99_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout449 net450 vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__buf_2
XFILLER_87_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06800__Y _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09753_ net381 _04388_ net311 vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__o21bai_1
X_06965_ net914 _01800_ vssd1 vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_107_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08137__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08704_ _03008_ _03030_ vssd1 vssd1 vccd1 vccd1 _03540_ sky130_fd_sc_hd__and2_1
X_09684_ _03566_ _04518_ _03604_ vssd1 vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__a21oi_1
X_06896_ _01629_ _01638_ _01656_ net961 vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__and4_1
X_08635_ _01935_ _01956_ vssd1 vssd1 vccd1 vccd1 _03471_ sky130_fd_sc_hd__nand2_1
XFILLER_55_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07631__Y _02467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08566_ datapath.rf.registers\[3\]\[0\] _01788_ _01797_ vssd1 vssd1 vccd1 vccd1 _03402_
+ sky130_fd_sc_hd__and3_1
XFILLER_70_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07998__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07517_ net872 _02350_ _02351_ _02352_ vssd1 vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__or4_1
XFILLER_22_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08497_ datapath.rf.registers\[13\]\[1\] net970 _01823_ vssd1 vssd1 vccd1 vccd1 _03333_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout714_A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07448_ net612 _02283_ net564 vssd1 vssd1 vccd1 vccd1 _02284_ sky130_fd_sc_hd__a21oi_2
XFILLER_156_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07379_ datapath.rf.registers\[17\]\[23\] net849 net836 datapath.rf.registers\[26\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1244_X net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11747__B2 _03028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09118_ _03587_ _03951_ vssd1 vssd1 vccd1 vccd1 _03954_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_118_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07415__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10390_ net559 net558 net452 vssd1 vssd1 vccd1 vccd1 _05226_ sky130_fd_sc_hd__mux2_1
XFILLER_136_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09049_ net551 net547 _02125_ vssd1 vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__a21o_1
XFILLER_136_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12060_ _06090_ _06091_ _06092_ _06100_ vssd1 vssd1 vccd1 vccd1 _06101_ sky130_fd_sc_hd__or4_1
XFILLER_151_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold470 datapath.rf.registers\[30\]\[1\] vssd1 vssd1 vccd1 vccd1 net1818 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout871_X net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold481 datapath.rf.registers\[13\]\[0\] vssd1 vssd1 vccd1 vccd1 net1829 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout969_X net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08376__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold492 datapath.rf.registers\[14\]\[16\] vssd1 vssd1 vccd1 vccd1 net1840 sky130_fd_sc_hd__dlygate4sd3_1
X_11011_ net282 net2464 net540 vssd1 vssd1 vccd1 vccd1 _00073_ sky130_fd_sc_hd__mux2_1
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout961 net962 vssd1 vssd1 vccd1 vccd1 net961 sky130_fd_sc_hd__clkbuf_2
Xfanout983 net989 vssd1 vssd1 vccd1 vccd1 net983 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08128__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout994 _01567_ vssd1 vssd1 vccd1 vccd1 net994 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_51_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12962_ net207 net2477 net481 vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__mux2_1
Xhold1170 screen.register.currentYbus\[7\] vssd1 vssd1 vccd1 vccd1 net2518 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input10_A DAT_I[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09750__A _04146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1181 datapath.rf.registers\[29\]\[31\] vssd1 vssd1 vccd1 vccd1 net2529 sky130_fd_sc_hd__dlygate4sd3_1
X_11913_ net136 _05972_ _05971_ vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__o21ai_1
XFILLER_45_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1192 datapath.rf.registers\[6\]\[17\] vssd1 vssd1 vccd1 vccd1 net2540 sky130_fd_sc_hd__dlygate4sd3_1
X_12893_ net172 net1834 net398 vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__mux2_1
XFILLER_72_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11491__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11844_ _05344_ _05922_ vssd1 vssd1 vccd1 vccd1 _05923_ sky130_fd_sc_hd__nor2_1
X_14632_ clknet_leaf_63_clk _01337_ net1234 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11435__A0 _05653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14563_ clknet_leaf_119_clk _01268_ net1194 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11775_ _01432_ _05892_ vssd1 vssd1 vccd1 vccd1 _05893_ sky130_fd_sc_hd__or2_2
XFILLER_14_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_155_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13514_ clknet_leaf_60_clk _00324_ net1167 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10726_ net1682 _02750_ net573 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[12\]
+ sky130_fd_sc_hd__mux2_1
X_14494_ clknet_leaf_150_clk _01199_ net1059 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10915__A2_N _05657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13445_ clknet_leaf_117_clk _00255_ net1188 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10657_ _05437_ _05439_ vssd1 vssd1 vccd1 vccd1 _05476_ sky130_fd_sc_hd__or2_1
XANTENNA__10835__S net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload15 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 clkload15/X sky130_fd_sc_hd__clkbuf_8
Xclkload26 clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 clkload26/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload37 clknet_leaf_139_clk vssd1 vssd1 vccd1 vccd1 clkload37/Y sky130_fd_sc_hd__bufinv_16
X_13376_ clknet_leaf_135_clk _00186_ net1104 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_58_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10588_ _02046_ _02090_ _02145_ _02189_ vssd1 vssd1 vccd1 vccd1 _05411_ sky130_fd_sc_hd__or4_1
XFILLER_127_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload48 clknet_leaf_129_clk vssd1 vssd1 vccd1 vccd1 clkload48/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload59 clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 clkload59/Y sky130_fd_sc_hd__inv_8
X_12327_ _05619_ _06254_ vssd1 vssd1 vccd1 vccd1 _06300_ sky130_fd_sc_hd__nor2_1
XANTENNA__10410__A1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12258_ net1269 _05002_ net222 _04837_ vssd1 vssd1 vccd1 vccd1 _06249_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_71_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06901__X _01737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11209_ net260 net1982 net529 vssd1 vssd1 vccd1 vccd1 _00259_ sky130_fd_sc_hd__mux2_1
XANTENNA__10174__B1 _01702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12351__A net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12189_ screen.counter.ct\[21\] _06166_ net601 vssd1 vssd1 vccd1 vccd1 _06204_ sky130_fd_sc_hd__and3_1
XFILLER_96_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06987__C _01647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08119__B1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06750_ _01579_ _01588_ vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__or2_1
XFILLER_36_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06681_ datapath.ru.latched_instruction\[11\] _01475_ _01490_ datapath.ru.latched_instruction\[10\]
+ vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__a22o_1
XANTENNA__11674__B1 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12497__S net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_69_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08547__Y _03383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08420_ _03252_ _03253_ _03254_ _03255_ vssd1 vssd1 vccd1 vccd1 _03256_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_102_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08351_ datapath.rf.registers\[3\]\[3\] net988 net927 vssd1 vssd1 vccd1 vccd1 _03187_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_22_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07302_ datapath.rf.registers\[1\]\[25\] net764 _02137_ net788 vssd1 vssd1 vccd1
+ vccd1 _02138_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_82_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08282_ datapath.rf.registers\[22\]\[5\] net735 net669 datapath.rf.registers\[21\]\[5\]
+ _03117_ vssd1 vssd1 vccd1 vccd1 _03118_ sky130_fd_sc_hd__a221o_1
XFILLER_60_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07645__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08842__A1 _01666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload9 clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clkload9/Y sky130_fd_sc_hd__inv_8
X_07233_ datapath.rf.registers\[0\]\[26\] net866 _02058_ _02068_ vssd1 vssd1 vccd1
+ vccd1 _02069_ sky130_fd_sc_hd__o22a_4
XANTENNA_fanout128_A _06369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13121__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07164_ _01988_ _01991_ _01992_ _01999_ vssd1 vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__or4_1
XFILLER_145_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07095_ datapath.rf.registers\[10\]\[29\] net880 net819 datapath.rf.registers\[5\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__a22o_1
XANTENNA__12960__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06811__X _01647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11692__A2_N _05885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14212__RESET_B net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout202 _05646_ vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__buf_1
XANTENNA_fanout497_A _06550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout213 _05634_ vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__buf_1
Xfanout224 net226 vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12261__A net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1204_A net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout235 _05616_ vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__clkbuf_2
XFILLER_141_691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11901__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout246 _05599_ vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__07355__A _02170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input2_A DAT_I[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout257 _05582_ vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__clkbuf_2
X_09805_ net317 _04267_ _04634_ _04635_ _04640_ vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_89_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout268 net269 vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__clkbuf_2
X_07997_ datapath.rf.registers\[9\]\[10\] net984 net944 vssd1 vssd1 vccd1 vccd1 _02833_
+ sky130_fd_sc_hd__and3_1
Xfanout279 _05554_ vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__buf_1
XANTENNA_fanout664_A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09736_ net329 _04407_ net330 vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__o21a_1
X_06948_ _01703_ _01783_ vssd1 vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__nor2_2
XFILLER_27_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09667_ net362 _04377_ _04404_ net373 vssd1 vssd1 vccd1 vccd1 _04503_ sky130_fd_sc_hd__o211a_1
X_06879_ _01629_ _01639_ _01657_ net961 vssd1 vssd1 vccd1 vccd1 _01715_ sky130_fd_sc_hd__and4_2
XFILLER_54_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08530__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout929_A _01727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08618_ _02441_ _03452_ _02443_ _02333_ _02387_ vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07802__B net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09598_ _04303_ _04307_ net454 vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__mux2_1
XFILLER_70_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07884__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08549_ datapath.rf.registers\[24\]\[0\] net965 net912 net908 vssd1 vssd1 vccd1 vccd1
+ _03385_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout717_X net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11560_ net1007 _05783_ vssd1 vssd1 vccd1 vccd1 _05784_ sky130_fd_sc_hd__nor2_1
XANTENNA__12090__B1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07636__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10511_ _05337_ _05338_ _05339_ _05340_ vssd1 vssd1 vccd1 vccd1 _05341_ sky130_fd_sc_hd__and4_1
X_11491_ net255 net2237 net513 vssd1 vssd1 vccd1 vccd1 _00527_ sky130_fd_sc_hd__mux2_1
XANTENNA__13031__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13230_ clknet_leaf_0_clk _00040_ net1055 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10442_ net891 _05273_ _05277_ net227 vssd1 vssd1 vccd1 vccd1 _05278_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_150_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08352__C net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13161_ net260 net1900 net544 vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__mux2_1
XFILLER_156_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12870__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10373_ _05205_ _05208_ net227 vssd1 vssd1 vccd1 vccd1 _05209_ sky130_fd_sc_hd__o21ai_1
XFILLER_152_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10943__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12112_ screen.counter.currentCt\[17\] screen.counter.currentCt\[16\] screen.counter.currentCt\[19\]
+ screen.counter.currentCt\[18\] vssd1 vssd1 vccd1 vccd1 _06149_ sky130_fd_sc_hd__or4_1
XFILLER_2_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13092_ net1939 net172 net388 vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11486__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12043_ screen.register.currentYbus\[11\] _05776_ net995 screen.register.currentXbus\[3\]
+ _06084_ vssd1 vssd1 vccd1 vccd1 _06085_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_148_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10403__B _03384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout780 _01794_ vssd1 vssd1 vccd1 vccd1 net780 sky130_fd_sc_hd__clkbuf_8
Xfanout791 net792 vssd1 vssd1 vccd1 vccd1 net791 sky130_fd_sc_hd__clkbuf_8
XFILLER_93_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13994_ clknet_leaf_112_clk _00771_ net1197 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12945_ net244 net2479 net394 vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__mux2_1
XANTENNA__07712__B net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12876_ net257 net1832 net399 vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__mux2_1
XANTENNA__07875__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08527__C net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14615_ clknet_leaf_131_clk _01320_ net1114 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11827_ keypad.alpha _05906_ vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09077__A1 _03892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07088__B1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12081__B1 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11758_ net1500 net146 net141 _02487_ vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__a22o_1
XANTENNA__07627__A2 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14546_ clknet_leaf_32_clk _01251_ net1123 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10709_ net1464 _02680_ net571 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i_n\[14\]
+ sky130_fd_sc_hd__mux2_1
X_11689_ _05050_ net153 net148 net1498 vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__a22o_1
X_14477_ clknet_leaf_131_clk _01182_ net1113 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload104 clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 clkload104/X sky130_fd_sc_hd__clkbuf_4
Xclkload115 clknet_leaf_112_clk vssd1 vssd1 vccd1 vccd1 clkload115/Y sky130_fd_sc_hd__clkinv_2
X_13428_ clknet_leaf_128_clk _00238_ net1209 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload126 clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 clkload126/Y sky130_fd_sc_hd__clkinv_4
Xclkload137 clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 clkload137/Y sky130_fd_sc_hd__clkinv_4
Xclkload148 clknet_leaf_84_clk vssd1 vssd1 vccd1 vccd1 clkload148/Y sky130_fd_sc_hd__inv_8
XANTENNA__12780__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13359_ clknet_leaf_26_clk _00169_ net1137 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08830__Y _03666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire465_A _02238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11396__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06998__B _01825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07920_ _02754_ _02755_ vssd1 vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__or2_1
XFILLER_130_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07012__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10698__A1 _03227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07851_ datapath.rf.registers\[17\]\[13\] net852 vssd1 vssd1 vccd1 vccd1 _02687_
+ sky130_fd_sc_hd__and2_1
XFILLER_110_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06802_ _01453_ net1002 net1018 net1027 datapath.ru.latched_instruction\[18\] vssd1
+ vssd1 vccd1 vccd1 _01638_ sky130_fd_sc_hd__a32oi_4
XFILLER_111_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput2 DAT_I[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
X_07782_ _02616_ _02617_ vssd1 vssd1 vccd1 vccd1 _02618_ sky130_fd_sc_hd__nor2_1
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09521_ net360 _04355_ _04356_ net326 vssd1 vssd1 vccd1 vccd1 _04357_ sky130_fd_sc_hd__o211a_1
X_06733_ _01571_ vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__inv_2
XFILLER_80_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13116__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09452_ net364 _04124_ _04196_ net374 vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__a211o_1
X_06664_ mmio.memload_or_instruction\[26\] net1050 vssd1 vssd1 vccd1 vccd1 _01503_
+ sky130_fd_sc_hd__and2_2
XFILLER_92_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08403_ datapath.rf.registers\[5\]\[2\] net948 net936 vssd1 vssd1 vccd1 vccd1 _03239_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08437__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09383_ net352 _04213_ vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__and2_1
X_06595_ keypad.decode.push net1486 net1022 vssd1 vssd1 vccd1 vccd1 keypad.decode.sticky_n\[4\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12955__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07079__B1 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08334_ _03156_ _03165_ _03169_ net782 datapath.rf.registers\[0\]\[4\] vssd1 vssd1
+ vccd1 vccd1 _03170_ sky130_fd_sc_hd__o32a_4
XANTENNA__12072__B1 _06018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07618__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08265_ datapath.rf.registers\[11\]\[5\] net882 _03099_ _03100_ vssd1 vssd1 vccd1
+ vccd1 _03101_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout412_A _05730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12256__A net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1154_A net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07216_ datapath.rf.registers\[8\]\[26\] net876 net796 datapath.rf.registers\[29\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_99_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08196_ _03009_ _03030_ vssd1 vssd1 vccd1 vccd1 _03032_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_115_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07147_ datapath.rf.registers\[10\]\[28\] net708 _01824_ datapath.rf.registers\[13\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01983_ sky130_fd_sc_hd__a22o_1
XANTENNA__08043__A2 _02876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07251__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07078_ datapath.rf.registers\[20\]\[29\] net958 net923 vssd1 vssd1 vccd1 vccd1 _01914_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout781_A _01794_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout879_A net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09528__C1 _01607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1008 net1009 vssd1 vssd1 vccd1 vccd1 net1008 sky130_fd_sc_hd__buf_2
XFILLER_59_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1019 net1020 vssd1 vssd1 vccd1 vccd1 net1019 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout667_X net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09719_ net344 net320 _04018_ _04554_ vssd1 vssd1 vccd1 vccd1 _04555_ sky130_fd_sc_hd__a31o_1
X_10991_ net1552 net212 net435 vssd1 vssd1 vccd1 vccd1 _00056_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout834_X net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13026__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08628__B _02190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09700__C1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ _05696_ _06370_ vssd1 vssd1 vccd1 vccd1 _06549_ sky130_fd_sc_hd__nor2_4
XANTENNA__07857__A2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08347__C net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12661_ datapath.mulitply_result\[25\] datapath.multiplication_module.multiplicand_i\[25\]
+ vssd1 vssd1 vccd1 vccd1 _06498_ sky130_fd_sc_hd__and2_1
XFILLER_31_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12865__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11612_ _05331_ _05830_ _05835_ vssd1 vssd1 vccd1 vccd1 _05836_ sky130_fd_sc_hd__o21ai_1
XFILLER_30_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14400_ clknet_leaf_133_clk _01105_ net1112 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_12592_ datapath.mulitply_result\[14\] datapath.multiplication_module.multiplicand_i\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06440_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_46_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08644__A _01706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11543_ _05766_ vssd1 vssd1 vccd1 vccd1 _05767_ sky130_fd_sc_hd__inv_2
X_14331_ clknet_leaf_38_clk _01036_ net1145 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11810__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08282__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11070__A _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14262_ clknet_leaf_141_clk _00967_ net1095 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_11474_ net1755 net172 net408 vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__mux2_1
XFILLER_137_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13213_ clknet_leaf_144_clk _00023_ net1085 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10425_ net377 _04525_ _05260_ net331 vssd1 vssd1 vccd1 vccd1 _05261_ sky130_fd_sc_hd__o211a_1
XANTENNA__12366__B2 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08034__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14193_ clknet_leaf_90_clk datapath.multiplication_module.multiplicand_i_n\[4\] net1239
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[4\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__07242__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13144_ net1883 net243 net383 vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__mux2_1
XFILLER_3_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10356_ datapath.PC\[8\] _03735_ vssd1 vssd1 vccd1 vccd1 _05192_ sky130_fd_sc_hd__nand2_1
XFILLER_140_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08990__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13075_ net2087 net255 net387 vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__mux2_1
XFILLER_112_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10414__A _03262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10287_ _04844_ _04845_ vssd1 vssd1 vccd1 vccd1 _05123_ sky130_fd_sc_hd__or2_1
X_12026_ net1010 _06063_ _06068_ net1001 _06026_ vssd1 vssd1 vccd1 vccd1 _06069_ sky130_fd_sc_hd__a221o_1
XFILLER_66_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08819__A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13977_ clknet_leaf_107_clk _00755_ net1223 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[20\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_74_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06984__D _01666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12928_ _05695_ _05734_ vssd1 vssd1 vccd1 vccd1 _06555_ sky130_fd_sc_hd__nand2_4
XANTENNA__12775__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12859_ net182 net2190 net487 vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__mux2_1
XFILLER_33_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11899__B net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12054__B1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14529_ clknet_leaf_46_clk _01234_ net1172 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11801__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08273__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08050_ datapath.rf.registers\[31\]\[9\] net977 net915 vssd1 vssd1 vccd1 vccd1 _02886_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07481__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12357__A1 _05002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07001_ datapath.rf.registers\[30\]\[31\] net758 net750 datapath.rf.registers\[28\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__a22o_1
XANTENNA__08025__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13857__RESET_B net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08952_ net341 _03782_ _03787_ net320 vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_110_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07903_ datapath.rf.registers\[19\]\[12\] net854 net791 datapath.rf.registers\[18\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__a22o_1
X_08883_ net566 _03718_ _01856_ vssd1 vssd1 vccd1 vccd1 _03719_ sky130_fd_sc_hd__or3b_1
XANTENNA__09911__A_N _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout195_A _05659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07834_ datapath.rf.registers\[17\]\[14\] net747 net688 datapath.rf.registers\[31\]\[14\]
+ _02667_ vssd1 vssd1 vccd1 vccd1 _02670_ sky130_fd_sc_hd__a221o_1
XFILLER_56_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07765_ datapath.rf.registers\[22\]\[15\] net822 net817 datapath.rf.registers\[7\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02601_ sky130_fd_sc_hd__a22o_1
X_06716_ mmio.memload_or_instruction\[17\] mmio.memload_or_instruction\[18\] mmio.memload_or_instruction\[15\]
+ mmio.memload_or_instruction\[16\] vssd1 vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__or4bb_1
X_09504_ _02912_ _02960_ net452 vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__mux2_1
XANTENNA__12293__B1 _06253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07839__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07696_ datapath.rf.registers\[14\]\[17\] net776 net704 datapath.rf.registers\[9\]\[17\]
+ _02529_ vssd1 vssd1 vccd1 vccd1 _02532_ sky130_fd_sc_hd__a221o_1
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09435_ net607 _04241_ _04270_ net555 vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__o211a_1
X_06647_ mmio.key_data\[6\] net1049 _01484_ vssd1 vssd1 vccd1 vccd1 _01486_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout150_X net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout627_A net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09366_ net574 _04193_ _04194_ _04201_ vssd1 vssd1 vccd1 vccd1 _04202_ sky130_fd_sc_hd__a22o_1
X_06578_ net1 vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__inv_2
XFILLER_24_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08317_ datapath.rf.registers\[21\]\[4\] net668 net665 datapath.rf.registers\[15\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__a22o_1
XANTENNA__08264__A2 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09297_ _04129_ _04132_ vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__nor2_1
XANTENNA__09461__A1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout415_X net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07472__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08248_ datapath.rf.registers\[10\]\[5\] net983 net937 vssd1 vssd1 vccd1 vccd1 _03084_
+ sky130_fd_sc_hd__and3_1
XFILLER_107_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08016__A2 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08179_ _03013_ _03014_ vssd1 vssd1 vccd1 vccd1 _03015_ sky130_fd_sc_hd__or2_1
X_10210_ _04586_ _04600_ net894 vssd1 vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__a21o_1
XFILLER_137_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07224__B1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11190_ net244 net2045 net422 vssd1 vssd1 vccd1 vccd1 _00242_ sky130_fd_sc_hd__mux2_1
Xteam_04_1296 vssd1 vssd1 vccd1 vccd1 team_04_1296/HI gpio_oeb[1] sky130_fd_sc_hd__conb_1
XANTENNA__10505__Y _05335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout784_X net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10141_ net1265 net1260 _04974_ _04976_ vssd1 vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__o22a_1
XFILLER_121_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10072_ net224 _04907_ net1292 vssd1 vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__a21oi_1
XFILLER_102_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13900_ clknet_leaf_43_clk net1358 net1149 vssd1 vssd1 vccd1 vccd1 keypad.debounce.debounce\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_145_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10888__B _03978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13831_ clknet_leaf_116_clk _00640_ net1187 vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__dfrtp_1
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13762_ clknet_leaf_76_clk _00571_ net1248 vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__dfrtp_1
X_10974_ net1679 net295 net434 vssd1 vssd1 vccd1 vccd1 _00039_ sky130_fd_sc_hd__mux2_1
XFILLER_90_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10295__C1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12713_ net1916 _06537_ vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13693_ clknet_leaf_145_clk _00503_ net1088 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_12644_ _06481_ _06482_ _06483_ _06477_ vssd1 vssd1 vccd1 vccd1 _06484_ sky130_fd_sc_hd__a211o_1
XFILLER_31_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12575_ datapath.mulitply_result\[11\] datapath.multiplication_module.multiplicand_i\[11\]
+ vssd1 vssd1 vccd1 vccd1 _06426_ sky130_fd_sc_hd__and2_1
XANTENNA__08255__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11004__S net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14314_ clknet_leaf_58_clk _01019_ net1167 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11526_ screen.counter.ct\[1\] screen.counter.ct\[0\] vssd1 vssd1 vccd1 vccd1 _05750_
+ sky130_fd_sc_hd__or2_1
XFILLER_7_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14245_ clknet_leaf_124_clk datapath.multiplication_module.multiplier_i_n\[13\] net1215
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i\[13\] sky130_fd_sc_hd__dfrtp_1
X_11457_ datapath.rf.registers\[14\]\[13\] _05582_ net407 vssd1 vssd1 vccd1 vccd1
+ _00495_ sky130_fd_sc_hd__mux2_1
XANTENNA__08007__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07215__B1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10408_ _03547_ _03548_ vssd1 vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__xor2_1
X_14176_ clknet_leaf_47_clk _00931_ net1172 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11388_ net2001 net266 net412 vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__mux2_1
XFILLER_140_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10339_ _04860_ _04861_ vssd1 vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13950__RESET_B net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13127_ _05696_ _05713_ vssd1 vssd1 vccd1 vccd1 _06562_ sky130_fd_sc_hd__nor2_1
XANTENNA__09492__X _04328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13058_ net183 net2240 net474 vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__mux2_1
XFILLER_112_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12511__A1 datapath.multiplication_module.multiplier_i\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12009_ screen.register.currentXbus\[25\] _05772_ _05837_ screen.register.currentYbus\[17\]
+ vssd1 vssd1 vccd1 vccd1 _06053_ sky130_fd_sc_hd__a22o_1
XFILLER_94_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06995__C net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07550_ net613 _02385_ net564 vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_37_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07481_ datapath.rf.registers\[26\]\[21\] net778 net766 datapath.rf.registers\[24\]\[21\]
+ _02313_ vssd1 vssd1 vccd1 vccd1 _02317_ sky130_fd_sc_hd__a221o_1
XFILLER_34_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09220_ _03607_ _04025_ _04026_ _04027_ _04055_ vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__a221o_1
X_09151_ _03920_ _03986_ net368 vssd1 vssd1 vccd1 vccd1 _03987_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_8_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08102_ datapath.rf.registers\[16\]\[8\] _01707_ net930 vssd1 vssd1 vccd1 vccd1 _02938_
+ sky130_fd_sc_hd__and3_1
XFILLER_148_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09082_ _03589_ _03917_ net578 vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__o21ai_1
XFILLER_108_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08033_ datapath.rf.registers\[11\]\[10\] net712 net693 datapath.rf.registers\[13\]\[10\]
+ _02858_ vssd1 vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__a221o_1
Xhold800 screen.counter.currentCt\[10\] vssd1 vssd1 vccd1 vccd1 net2148 sky130_fd_sc_hd__dlygate4sd3_1
Xhold811 datapath.rf.registers\[25\]\[19\] vssd1 vssd1 vccd1 vccd1 net2159 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07206__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold822 datapath.rf.registers\[4\]\[12\] vssd1 vssd1 vccd1 vccd1 net2170 sky130_fd_sc_hd__dlygate4sd3_1
Xhold833 datapath.rf.registers\[23\]\[17\] vssd1 vssd1 vccd1 vccd1 net2181 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold844 datapath.rf.registers\[25\]\[16\] vssd1 vssd1 vccd1 vccd1 net2192 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold855 datapath.rf.registers\[5\]\[14\] vssd1 vssd1 vccd1 vccd1 net2203 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold866 datapath.rf.registers\[29\]\[9\] vssd1 vssd1 vccd1 vccd1 net2214 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold877 datapath.rf.registers\[9\]\[15\] vssd1 vssd1 vccd1 vccd1 net2225 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap585 net586 vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__clkbuf_1
Xhold888 datapath.rf.registers\[29\]\[19\] vssd1 vssd1 vccd1 vccd1 net2236 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09984_ _04816_ _04818_ _04819_ _04725_ vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__a31o_1
Xhold899 datapath.rf.registers\[2\]\[15\] vssd1 vssd1 vccd1 vccd1 net2247 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07797__A2_N net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07915__X _02751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09843__A _01859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08935_ net648 _03642_ _03641_ vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__a21o_1
XFILLER_29_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08866_ _02705_ _02751_ net444 vssd1 vssd1 vccd1 vccd1 _03702_ sky130_fd_sc_hd__mux2_1
X_07817_ datapath.rf.registers\[17\]\[14\] net850 net808 datapath.rf.registers\[27\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02653_ sky130_fd_sc_hd__a22o_1
X_08797_ net370 _03632_ _03627_ vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__o21ba_1
XFILLER_72_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout744_A net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07748_ datapath.rf.registers\[6\]\[16\] net679 net660 datapath.rf.registers\[5\]\[16\]
+ _02577_ vssd1 vssd1 vccd1 vccd1 _02584_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_123_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07679_ datapath.rf.registers\[30\]\[17\] net834 net802 datapath.rf.registers\[3\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02515_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout532_X net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12018__B1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09418_ _04252_ _04253_ net325 _04251_ vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__o2bb2a_1
X_10690_ _05458_ _05503_ _05504_ _05506_ vssd1 vssd1 vccd1 vccd1 keypad.decode.button_n\[3\]
+ sky130_fd_sc_hd__a211o_1
XANTENNA__07693__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08237__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09349_ _02567_ net553 net549 vssd1 vssd1 vccd1 vccd1 _04185_ sky130_fd_sc_hd__or3_1
XFILLER_8_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07445__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12360_ net229 _04898_ _06323_ net893 vssd1 vssd1 vccd1 vccd1 _06324_ sky130_fd_sc_hd__o211a_1
XFILLER_20_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout999_X net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11311_ net2491 net286 net417 vssd1 vssd1 vccd1 vccd1 _00356_ sky130_fd_sc_hd__mux2_1
XFILLER_138_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12291_ net634 _04562_ vssd1 vssd1 vccd1 vccd1 _06274_ sky130_fd_sc_hd__nand2_1
X_14030_ clknet_leaf_80_clk _00799_ net1257 vssd1 vssd1 vccd1 vccd1 datapath.PC\[20\]
+ sky130_fd_sc_hd__dfrtp_4
X_11242_ net260 net1836 net421 vssd1 vssd1 vccd1 vccd1 _00291_ sky130_fd_sc_hd__mux2_1
XFILLER_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08945__A0 _02264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11173_ _05695_ _05717_ vssd1 vssd1 vccd1 vccd1 _05719_ sky130_fd_sc_hd__nand2_1
XFILLER_122_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10124_ net640 _04057_ vssd1 vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__and2_1
XFILLER_122_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11494__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10055_ _04824_ _04890_ vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__xnor2_1
XFILLER_76_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13814_ clknet_leaf_113_clk _00623_ net1197 vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_3_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10268__C1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13745_ clknet_leaf_50_clk _00555_ net1181 vssd1 vssd1 vccd1 vccd1 mmio.key_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10838__S net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08476__A2 _01753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09673__A1 _02961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10957_ _05693_ _05694_ vssd1 vssd1 vccd1 vccd1 _05695_ sky130_fd_sc_hd__nor2_4
XFILLER_31_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13676_ clknet_leaf_17_clk _00486_ net1106 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10888_ net902 _03978_ vssd1 vssd1 vccd1 vccd1 _05635_ sky130_fd_sc_hd__or2_2
XFILLER_31_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12627_ _06461_ _06465_ _06468_ vssd1 vssd1 vccd1 vccd1 _06470_ sky130_fd_sc_hd__nand3_1
XANTENNA__08228__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07436__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06904__X _01740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12558_ _06406_ _06408_ _06405_ vssd1 vssd1 vccd1 vccd1 _06412_ sky130_fd_sc_hd__o21ba_1
XFILLER_145_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11509_ net168 net2423 net511 vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__mux2_1
XFILLER_156_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold107 net42 vssd1 vssd1 vccd1 vccd1 net1455 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08551__B _01800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12489_ net266 net2358 net507 vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__mux2_1
Xhold118 net76 vssd1 vssd1 vccd1 vccd1 net1466 sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 datapath.multiplication_module.multiplier_i\[3\] vssd1 vssd1 vccd1 vccd1
+ net1477 sky130_fd_sc_hd__dlygate4sd3_1
X_14228_ clknet_leaf_42_clk _00949_ net1144 vssd1 vssd1 vccd1 vccd1 columns.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13449__RESET_B net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08936__A0 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14159_ clknet_leaf_67_clk _00914_ net1239 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout609 _03607_ vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__clkbuf_4
X_06981_ net971 _01816_ vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__and2_1
X_08720_ _03173_ _03174_ vssd1 vssd1 vccd1 vccd1 _03556_ sky130_fd_sc_hd__or2_2
Xfanout1180 net1185 vssd1 vssd1 vccd1 vccd1 net1180 sky130_fd_sc_hd__clkbuf_4
Xfanout1191 net1194 vssd1 vssd1 vccd1 vccd1 net1191 sky130_fd_sc_hd__clkbuf_4
XFILLER_94_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08651_ _02004_ _03472_ vssd1 vssd1 vccd1 vccd1 _03487_ sky130_fd_sc_hd__nand2b_2
XFILLER_82_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07602_ datapath.rf.registers\[0\]\[19\] net783 net590 net562 vssd1 vssd1 vccd1 vccd1
+ _02438_ sky130_fd_sc_hd__a2bb2o_2
XTAP_TAPCELL_ROW_1_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08582_ net612 _03417_ _03384_ vssd1 vssd1 vccd1 vccd1 _03418_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_105_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09113__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07533_ datapath.rf.registers\[16\]\[20\] net738 net722 datapath.rf.registers\[18\]\[20\]
+ _02368_ vssd1 vssd1 vccd1 vccd1 _02369_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_105_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13124__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout158_A net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07464_ datapath.rf.registers\[29\]\[21\] net796 _02295_ _02299_ vssd1 vssd1 vccd1
+ vccd1 _02300_ sky130_fd_sc_hd__a211oi_1
X_09203_ net459 _04037_ _04038_ vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__and3_1
XANTENNA__08219__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07395_ datapath.rf.registers\[10\]\[23\] net706 net691 datapath.rf.registers\[13\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__a22o_1
XANTENNA__12963__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09134_ _03667_ _03968_ _03969_ _03959_ vssd1 vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__o22a_1
XFILLER_148_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09065_ _03893_ _03894_ net342 vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__mux2_1
XFILLER_135_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1234_A net1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08016_ datapath.rf.registers\[8\]\[10\] net878 net854 datapath.rf.registers\[19\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__a22o_1
XANTENNA__06650__A1 datapath.ru.latched_instruction\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold630 datapath.rf.registers\[3\]\[4\] vssd1 vssd1 vccd1 vccd1 net1978 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold641 datapath.rf.registers\[22\]\[6\] vssd1 vssd1 vccd1 vccd1 net1989 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout694_A net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold652 datapath.rf.registers\[18\]\[21\] vssd1 vssd1 vccd1 vccd1 net2000 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold663 datapath.rf.registers\[30\]\[26\] vssd1 vssd1 vccd1 vccd1 net2011 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07077__B net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold674 datapath.rf.registers\[26\]\[13\] vssd1 vssd1 vccd1 vccd1 net2022 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold685 datapath.rf.registers\[22\]\[31\] vssd1 vssd1 vccd1 vccd1 net2033 sky130_fd_sc_hd__dlygate4sd3_1
Xhold696 datapath.rf.registers\[15\]\[3\] vssd1 vssd1 vccd1 vccd1 net2044 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09967_ _04753_ _04757_ _04801_ _04752_ vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout861_A net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout482_X net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout959_A net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07805__B net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08918_ datapath.PC\[31\] _03752_ _03753_ vssd1 vssd1 vccd1 vccd1 _03754_ sky130_fd_sc_hd__o21ai_1
X_09898_ _01585_ net900 _01630_ vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__and3_1
X_08849_ _01935_ _01981_ net445 vssd1 vssd1 vccd1 vccd1 _03685_ sky130_fd_sc_hd__mux2_1
XFILLER_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout747_X net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11860_ net2273 net163 vssd1 vssd1 vccd1 vccd1 _05937_ sky130_fd_sc_hd__nand2_1
X_10811_ _01474_ net655 _05568_ _05569_ vssd1 vssd1 vccd1 vccd1 _05570_ sky130_fd_sc_hd__o22a_2
X_11791_ datapath.ru.ack_mul_reg2 net1016 _01590_ datapath.ru.ack_mul_reg vssd1 vssd1
+ vccd1 vccd1 _05903_ sky130_fd_sc_hd__or4bb_1
XANTENNA_fanout914_X net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13034__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13530_ clknet_leaf_146_clk _00340_ net1065 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10742_ net1519 net569 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[28\]
+ sky130_fd_sc_hd__and2_1
XFILLER_41_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07130__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10673_ net1013 _05489_ _05437_ vssd1 vssd1 vccd1 vccd1 _05491_ sky130_fd_sc_hd__o21ba_1
XFILLER_9_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13461_ clknet_leaf_19_clk _00271_ net1116 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12873__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08923__Y _03759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07418__B1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12412_ net1433 net131 _06353_ vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__a21o_1
XANTENNA__09748__A _04207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13392_ clknet_leaf_25_clk _00202_ net1158 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08652__A _02025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11489__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12343_ _06310_ _06311_ net1264 net310 vssd1 vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08091__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12274_ net2651 net309 _06261_ vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__a21o_1
XFILLER_5_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11225_ net241 net2074 net528 vssd1 vssd1 vccd1 vccd1 _00275_ sky130_fd_sc_hd__mux2_1
X_14013_ clknet_4_14_0_clk _00782_ net1252 vssd1 vssd1 vccd1 vccd1 datapath.PC\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_56_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07197__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11156_ net249 net2503 net531 vssd1 vssd1 vccd1 vccd1 _00209_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10107_ net229 _04938_ _04940_ _04942_ net1293 vssd1 vssd1 vccd1 vccd1 _04943_ sky130_fd_sc_hd__a311o_1
XFILLER_67_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11087_ net253 net2093 net534 vssd1 vssd1 vccd1 vccd1 _00144_ sky130_fd_sc_hd__mux2_1
XFILLER_49_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10038_ _04873_ _04834_ vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__and2b_1
XFILLER_91_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08449__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11989_ screen.register.currentXbus\[0\] _05755_ _06018_ screen.register.currentYbus\[0\]
+ _06033_ vssd1 vssd1 vccd1 vccd1 _06034_ sky130_fd_sc_hd__a221o_1
XFILLER_17_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07450__B _02284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13728_ clknet_leaf_137_clk _00538_ net1090 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_50_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13659_ clknet_leaf_38_clk _00469_ net1146 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12783__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_140_Right_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07180_ datapath.rf.registers\[4\]\[27\] net864 _02015_ net873 vssd1 vssd1 vccd1
+ vccd1 _02016_ sky130_fd_sc_hd__a211o_1
XANTENNA__11399__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08082__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_65_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07609__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout406 _05733_ vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__clkbuf_8
X_09821_ net341 _04655_ _04656_ net338 vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__o211a_1
Xfanout417 _05726_ vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__clkbuf_4
Xfanout428 net429 vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__clkbuf_8
Xfanout439 _03771_ vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkload12_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13119__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_123_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09752_ _03513_ _03580_ vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__xor2_1
X_06964_ net991 net972 vssd1 vssd1 vccd1 vccd1 _01800_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_107_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09334__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08703_ _02961_ _02983_ vssd1 vssd1 vccd1 vccd1 _03539_ sky130_fd_sc_hd__nor2_1
X_06895_ datapath.rf.registers\[9\]\[31\] net885 net856 datapath.rf.registers\[24\]\[31\]
+ _01729_ vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__a221o_1
XANTENNA__12958__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09683_ _03566_ _04518_ vssd1 vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__or2_1
XFILLER_82_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07896__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08634_ _02048_ _03469_ _02049_ vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_87_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_138_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08565_ _03388_ _03392_ _03396_ _03400_ vssd1 vssd1 vccd1 vccd1 _03401_ sky130_fd_sc_hd__or4_1
XANTENNA__09637__A1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout442_A net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09637__B2 _03607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1184_A net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08456__B net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07648__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07360__B net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07516_ datapath.rf.registers\[14\]\[20\] net830 _02334_ _02339_ _02340_ vssd1 vssd1
+ vccd1 vccd1 _02352_ sky130_fd_sc_hd__a2111o_1
XANTENNA_clkbuf_leaf_18_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08496_ datapath.rf.registers\[25\]\[1\] net729 _03329_ _03330_ _03331_ vssd1 vssd1
+ vccd1 vccd1 _03332_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07112__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07447_ _02270_ _02274_ _02282_ net782 datapath.rf.registers\[0\]\[22\] vssd1 vssd1
+ vccd1 vccd1 _02283_ sky130_fd_sc_hd__o32a_4
XANTENNA_fanout230_X net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout707_A net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07378_ datapath.rf.registers\[25\]\[23\] net841 net826 datapath.rf.registers\[12\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__a22o_1
XFILLER_148_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09117_ _03587_ _03951_ vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_118_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08073__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06704__B datapath.ru.latched_instruction\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11102__S net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09048_ _02069_ net553 net549 vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__or3_1
XANTENNA__07820__B1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout697_X net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold460 datapath.rf.registers\[16\]\[23\] vssd1 vssd1 vccd1 vccd1 net1808 sky130_fd_sc_hd__dlygate4sd3_1
Xhold471 datapath.rf.registers\[22\]\[29\] vssd1 vssd1 vccd1 vccd1 net1819 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold482 datapath.rf.registers\[28\]\[27\] vssd1 vssd1 vccd1 vccd1 net1830 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07179__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11010_ net292 net1857 net538 vssd1 vssd1 vccd1 vccd1 _00072_ sky130_fd_sc_hd__mux2_1
Xhold493 datapath.rf.registers\[3\]\[27\] vssd1 vssd1 vccd1 vccd1 net1841 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06720__A _01441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout864_X net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout940 _01717_ vssd1 vssd1 vccd1 vccd1 net940 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06926__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13029__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout962 _01678_ vssd1 vssd1 vccd1 vccd1 net962 sky130_fd_sc_hd__buf_1
Xfanout973 net974 vssd1 vssd1 vccd1 vccd1 net973 sky130_fd_sc_hd__buf_2
Xfanout984 net987 vssd1 vssd1 vccd1 vccd1 net984 sky130_fd_sc_hd__clkbuf_2
Xfanout995 _05792_ vssd1 vssd1 vccd1 vccd1 net995 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_51_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12961_ _05518_ _05729_ vssd1 vssd1 vccd1 vccd1 _06556_ sky130_fd_sc_hd__or2_4
XANTENNA__09876__A1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12868__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1160 datapath.rf.registers\[30\]\[8\] vssd1 vssd1 vccd1 vccd1 net2508 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1171 datapath.rf.registers\[28\]\[20\] vssd1 vssd1 vccd1 vccd1 net2519 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1182 datapath.rf.registers\[14\]\[3\] vssd1 vssd1 vccd1 vccd1 net2530 sky130_fd_sc_hd__dlygate4sd3_1
X_11912_ _02487_ net657 vssd1 vssd1 vccd1 vccd1 _05972_ sky130_fd_sc_hd__nand2_1
Xhold1193 mmio.memload_or_instruction\[8\] vssd1 vssd1 vccd1 vccd1 net2541 sky130_fd_sc_hd__dlygate4sd3_1
X_12892_ net181 net2298 net399 vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__mux2_1
XANTENNA__08647__A _01935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07351__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07551__A _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14631_ clknet_leaf_145_clk _01336_ net1089 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11843_ _05819_ _05921_ vssd1 vssd1 vccd1 vccd1 _05922_ sky130_fd_sc_hd__nand2_1
XFILLER_72_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07639__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07270__B net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14562_ clknet_leaf_152_clk _01267_ net1054 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11774_ columns.count\[0\] _01433_ vssd1 vssd1 vccd1 vccd1 _05892_ sky130_fd_sc_hd__nand2_1
XANTENNA__07103__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13513_ clknet_leaf_91_clk _00323_ net1241 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10725_ net1778 _02804_ net572 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[11\]
+ sky130_fd_sc_hd__mux2_1
X_14493_ clknet_leaf_149_clk _01198_ net1060 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13444_ clknet_leaf_19_clk _00254_ net1119 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10656_ _05443_ _05450_ _05471_ _05447_ vssd1 vssd1 vccd1 vccd1 _05475_ sky130_fd_sc_hd__a31o_1
XANTENNA__06862__B2 datapath.ru.latched_instruction\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_155_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload16 clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 clkload16/Y sky130_fd_sc_hd__clkinv_2
X_10587_ _05406_ _05407_ _05408_ _05409_ vssd1 vssd1 vccd1 vccd1 _05410_ sky130_fd_sc_hd__or4_1
Xclkload27 clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 clkload27/Y sky130_fd_sc_hd__clkinv_2
X_13375_ clknet_leaf_13_clk _00185_ net1079 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload38 clknet_leaf_140_clk vssd1 vssd1 vccd1 vccd1 clkload38/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload49 clknet_leaf_130_clk vssd1 vssd1 vccd1 vccd1 clkload49/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__11012__S net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12326_ net894 _04834_ net191 vssd1 vssd1 vccd1 vccd1 _06299_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07811__B1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10136__B _04023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12257_ _01416_ net308 vssd1 vssd1 vccd1 vccd1 _06248_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_71_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11208_ net207 net2322 net529 vssd1 vssd1 vccd1 vccd1 _00258_ sky130_fd_sc_hd__mux2_1
X_12188_ screen.counter.ct\[21\] _06201_ _06203_ vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__a21o_1
XANTENNA__10174__A1 _03947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06987__D net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11139_ _05707_ _05712_ vssd1 vssd1 vccd1 vccd1 _05717_ sky130_fd_sc_hd__nor2_1
XANTENNA__09316__A0 _02523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07590__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12778__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07732__Y _02568_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06680_ _01512_ _01516_ _01517_ _01518_ vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__or4_1
XANTENNA__11674__A1 _05281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire1045_X net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07342__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08350_ datapath.rf.registers\[12\]\[3\] net956 _01744_ vssd1 vssd1 vccd1 vccd1 _03186_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_22_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07301_ datapath.rf.registers\[25\]\[25\] net728 net704 datapath.rf.registers\[9\]\[25\]
+ _02136_ vssd1 vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__a221o_1
XFILLER_149_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08281_ datapath.rf.registers\[19\]\[5\] net731 _03115_ _03116_ net787 vssd1 vssd1
+ vccd1 vccd1 _03117_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_82_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_152_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_152_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_82_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07232_ _02060_ _02063_ _02065_ _02067_ vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__or4_1
XFILLER_149_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_4_Left_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08292__A net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11729__A2 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07163_ _01994_ _01996_ _01998_ vssd1 vssd1 vccd1 vccd1 _01999_ sky130_fd_sc_hd__or3_1
XFILLER_145_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07094_ datapath.rf.registers\[16\]\[29\] net860 net808 datapath.rf.registers\[27\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__a22o_1
XFILLER_117_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10761__S net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout203 _05641_ vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__clkbuf_2
XFILLER_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_130_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout214 net215 vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__clkbuf_2
Xfanout225 net226 vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__buf_2
XANTENNA_fanout392_A net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout236 _05616_ vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__clkbuf_1
Xfanout247 net250 vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__clkbuf_2
X_09804_ net905 _04628_ _04639_ vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__a21oi_1
Xfanout258 net261 vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07355__B _02190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout269 _05570_ vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_89_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07996_ datapath.rf.registers\[16\]\[10\] _01707_ net929 vssd1 vssd1 vccd1 vccd1
+ _02832_ sky130_fd_sc_hd__and3_1
XFILLER_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09735_ net647 _04570_ _03770_ vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__o21ai_1
X_06947_ _01591_ net897 vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__nand2_1
XFILLER_39_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09666_ net648 _04501_ net438 vssd1 vssd1 vccd1 vccd1 _04502_ sky130_fd_sc_hd__a21o_1
XFILLER_82_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06878_ _01657_ net961 vssd1 vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__and2_1
XANTENNA__07333__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08617_ _02441_ _03452_ _02443_ vssd1 vssd1 vccd1 vccd1 _03453_ sky130_fd_sc_hd__a21o_1
XFILLER_27_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07802__C net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout824_A net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09597_ net455 _04280_ _04431_ net353 vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__a211o_1
XFILLER_43_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08818__C1 _03384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08548_ MemWrite _01644_ _01780_ net992 vssd1 vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__a22o_4
XTAP_TAPCELL_ROW_137_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08294__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_143_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_143_clk
+ sky130_fd_sc_hd__clkbuf_8
X_08479_ datapath.rf.registers\[24\]\[1\] net858 _03299_ _03300_ _03303_ vssd1 vssd1
+ vccd1 vccd1 _03315_ sky130_fd_sc_hd__a2111o_1
X_10510_ screen.counter.ct\[0\] screen.counter.ct\[3\] screen.counter.ct\[22\] vssd1
+ vssd1 vccd1 vccd1 _05340_ sky130_fd_sc_hd__nor3_1
X_11490_ net264 net2083 net513 vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__mux2_1
XFILLER_137_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10441_ net1044 _05276_ _05275_ net636 vssd1 vssd1 vccd1 vccd1 _05277_ sky130_fd_sc_hd__a211o_1
XANTENNA__09243__C1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10928__B1 _05668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13160_ net209 net2343 net544 vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__mux2_1
X_10372_ net1269 net1039 _05207_ net891 vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout981_X net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12111_ screen.counter.currentCt\[9\] screen.counter.currentCt\[8\] screen.counter.currentCt\[11\]
+ _06147_ vssd1 vssd1 vccd1 vccd1 _06148_ sky130_fd_sc_hd__or4_1
X_13091_ net1636 net183 net387 vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__mux2_1
XANTENNA__09745__B _04580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12042_ screen.register.currentYbus\[27\] _05786_ net996 screen.register.currentXbus\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06084_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_53_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10156__A1 _04084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold290 datapath.rf.registers\[19\]\[11\] vssd1 vssd1 vccd1 vccd1 net1638 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07265__B net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_148_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout770 net773 vssd1 vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__buf_4
XFILLER_1_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07572__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout781 _01794_ vssd1 vssd1 vccd1 vccd1 net781 sky130_fd_sc_hd__buf_2
Xfanout792 _01776_ vssd1 vssd1 vccd1 vccd1 net792 sky130_fd_sc_hd__clkbuf_8
X_13993_ clknet_leaf_112_clk _00770_ net1198 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12944_ net247 net2501 net394 vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__mux2_1
XFILLER_34_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07324__A2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07712__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12875_ net265 net2121 net400 vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__mux2_1
XANTENNA__11007__S net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06626__D_N mmio.memload_or_instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14614_ clknet_leaf_138_clk _01319_ net1100 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_11826_ _01427_ _05895_ button\[4\] _05874_ vssd1 vssd1 vccd1 vccd1 _05906_ sky130_fd_sc_hd__or4b_1
XANTENNA__08285__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14545_ clknet_leaf_40_clk _01250_ net1140 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11757_ net1478 net143 net138 _02542_ vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__a22o_1
XANTENNA__10846__S net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_134_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_134_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_64_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10708_ net1458 _02725_ net571 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i_n\[13\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14476_ clknet_leaf_16_clk _01181_ net1108 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11688_ _05031_ net153 net148 net1437 vssd1 vssd1 vccd1 vccd1 _00573_ sky130_fd_sc_hd__a22o_1
XFILLER_146_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload105 clknet_leaf_125_clk vssd1 vssd1 vccd1 vccd1 clkload105/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__08037__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13427_ clknet_leaf_34_clk _00237_ net1127 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10639_ _05448_ _05450_ vssd1 vssd1 vccd1 vccd1 _05459_ sky130_fd_sc_hd__nand2_1
Xclkload116 clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 clkload116/Y sky130_fd_sc_hd__bufinv_16
Xclkload127 clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 clkload127/Y sky130_fd_sc_hd__inv_6
XANTENNA__12384__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload138 clknet_leaf_85_clk vssd1 vssd1 vccd1 vccd1 clkload138/X sky130_fd_sc_hd__clkbuf_8
X_13358_ clknet_leaf_0_clk _00168_ net1057 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_12309_ net228 _04863_ vssd1 vssd1 vccd1 vccd1 _06287_ sky130_fd_sc_hd__nor2_1
XANTENNA__10434__X _05270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13289_ clknet_leaf_91_clk _00099_ net1233 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07850_ datapath.rf.registers\[21\]\[13\] net946 net923 vssd1 vssd1 vccd1 vccd1 _02686_
+ sky130_fd_sc_hd__and3_1
XFILLER_111_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06801_ net1004 net1020 _01634_ _01633_ vssd1 vssd1 vccd1 vccd1 _01637_ sky130_fd_sc_hd__a31o_4
X_07781_ datapath.rf.registers\[3\]\[15\] net771 net763 datapath.rf.registers\[1\]\[15\]
+ _02614_ vssd1 vssd1 vccd1 vccd1 _02617_ sky130_fd_sc_hd__a221o_1
Xinput3 DAT_I[10] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
X_09520_ net351 _04344_ _04348_ net358 vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__a211o_1
XANTENNA__13193__A datapath.rf.registers\[0\]\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06732_ net1002 net1018 _01569_ _01570_ vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__a31oi_4
XTAP_TAPCELL_ROW_84_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06663_ mmio.key_data\[1\] mmio.memload_or_instruction\[1\] net1048 vssd1 vssd1 vccd1
+ vccd1 _01502_ sky130_fd_sc_hd__mux2_4
XFILLER_25_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09451_ net327 _04094_ vssd1 vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__nand2_1
XFILLER_80_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08402_ datapath.rf.registers\[23\]\[2\] net942 net926 vssd1 vssd1 vccd1 vccd1 _03238_
+ sky130_fd_sc_hd__and3_1
XFILLER_52_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06594_ columns.count\[0\] _01432_ _01433_ _01434_ vssd1 vssd1 vccd1 vccd1 _01435_
+ sky130_fd_sc_hd__or4bb_2
X_09382_ net458 _04161_ _04216_ net352 vssd1 vssd1 vccd1 vccd1 _04218_ sky130_fd_sc_hd__a211oi_1
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08333_ _03158_ _03161_ _03167_ _03168_ vssd1 vssd1 vccd1 vccd1 _03169_ sky130_fd_sc_hd__or4_1
Xclkbuf_leaf_125_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_125_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08276__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_49_Left_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout140_A net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13132__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout238_A _05616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08264_ datapath.rf.registers\[2\]\[5\] net888 net837 datapath.rf.registers\[26\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03100_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_15_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07215_ datapath.rf.registers\[14\]\[26\] net829 net793 datapath.rf.registers\[31\]\[26\]
+ _02050_ vssd1 vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__a221o_1
XANTENNA__08028__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08195_ _03009_ _03030_ vssd1 vssd1 vccd1 vccd1 _03031_ sky130_fd_sc_hd__and2_1
XANTENNA__12971__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout405_A _06549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09776__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07146_ datapath.rf.registers\[20\]\[28\] net721 net700 datapath.rf.registers\[23\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__a22o_1
XFILLER_106_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07077_ datapath.rf.registers\[1\]\[29\] net845 vssd1 vssd1 vccd1 vccd1 _01913_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_58_Left_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1009 _05748_ vssd1 vssd1 vccd1 vccd1 net1009 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout774_A _01796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout395_X net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07979_ datapath.rf.registers\[3\]\[11\] net772 net666 datapath.rf.registers\[15\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout941_A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12835__A0 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09718_ net337 _04553_ vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__and2_1
XANTENNA__10520__A _05335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10990_ net1615 net217 net434 vssd1 vssd1 vccd1 vccd1 _00055_ sky130_fd_sc_hd__mux2_1
XANTENNA__08197__A _03009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07306__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_143_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09649_ net331 _03958_ _04484_ _03613_ vssd1 vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout827_X net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12660_ _06492_ _06495_ _06491_ vssd1 vssd1 vccd1 vccd1 _06497_ sky130_fd_sc_hd__a21boi_1
XANTENNA__13386__RESET_B net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_67_Left_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11611_ net999 _05832_ _05833_ _05834_ vssd1 vssd1 vccd1 vccd1 _05835_ sky130_fd_sc_hd__or4_1
Xclkbuf_leaf_116_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_116_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12591_ net2379 net504 net500 _06439_ vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_46_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13042__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14330_ clknet_leaf_14_clk _01035_ net1078 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_129_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11542_ _05302_ _05765_ vssd1 vssd1 vccd1 vccd1 _05766_ sky130_fd_sc_hd__or2_1
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11070__B _01663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14261_ clknet_leaf_19_clk _00966_ net1119 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12881__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11473_ net2571 net181 net407 vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__mux2_1
XFILLER_143_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13212_ clknet_leaf_7_clk _00022_ net1073 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07227__D1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10424_ net329 _05256_ _05259_ vssd1 vssd1 vccd1 vccd1 _05260_ sky130_fd_sc_hd__or3_1
XFILLER_125_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08660__A _02169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14192_ clknet_leaf_90_clk datapath.multiplication_module.multiplicand_i_n\[3\] net1239
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[3\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11497__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13143_ net1856 net248 net382 vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_76_Left_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10355_ datapath.PC\[8\] _04515_ net466 vssd1 vssd1 vccd1 vccd1 _05191_ sky130_fd_sc_hd__mux2_1
XFILLER_152_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07793__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13074_ net1626 net262 net387 vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__mux2_1
X_10286_ net892 _04496_ _05117_ _05121_ vssd1 vssd1 vccd1 vccd1 _05122_ sky130_fd_sc_hd__o31a_1
XFILLER_140_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12025_ _06058_ _06065_ _06067_ vssd1 vssd1 vccd1 vccd1 _06068_ sky130_fd_sc_hd__or3_1
XANTENNA__11877__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07545__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13976_ clknet_leaf_105_clk _00754_ net1223 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12927_ net2324 net168 net482 vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__mux2_1
XFILLER_34_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_698 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_85_Left_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08173__A2_N net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12858_ net176 net2086 net489 vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__mux2_1
XFILLER_34_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08835__A _01609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06907__X _01743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11809_ _01510_ net1015 net314 net334 datapath.ru.latched_instruction\[15\] vssd1
+ vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__a32o_1
XANTENNA__08258__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_107_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_107_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12789_ net196 net1752 net496 vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__mux2_1
XFILLER_14_381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08554__B net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14528_ clknet_leaf_134_clk _01233_ net1112 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_32_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12791__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14459_ clknet_leaf_36_clk _01164_ net1135 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_07000_ datapath.rf.registers\[26\]\[31\] net778 net719 datapath.rf.registers\[20\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12357__A2 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_94_Left_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11200__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07784__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08951_ net341 _03786_ vssd1 vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_94_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07902_ datapath.rf.registers\[26\]\[12\] net838 net809 datapath.rf.registers\[27\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__a22o_1
XFILLER_97_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08882_ _01610_ _03716_ vssd1 vssd1 vccd1 vccd1 _03718_ sky130_fd_sc_hd__or2_2
XFILLER_111_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07536__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_4_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07833_ datapath.rf.registers\[2\]\[14\] net743 net684 datapath.rf.registers\[27\]\[14\]
+ _02668_ vssd1 vssd1 vccd1 vccd1 _02669_ sky130_fd_sc_hd__a221o_1
XFILLER_57_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout188_A _05664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07764_ datapath.rf.registers\[20\]\[15\] net839 net816 datapath.rf.registers\[21\]\[15\]
+ _02591_ vssd1 vssd1 vccd1 vccd1 _02600_ sky130_fd_sc_hd__a221o_1
XFILLER_37_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09503_ _03422_ _03550_ vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__xor2_1
XFILLER_112_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06715_ mmio.memload_or_instruction\[8\] _01553_ mmio.memload_or_instruction\[10\]
+ _01552_ vssd1 vssd1 vccd1 vccd1 _01554_ sky130_fd_sc_hd__or4b_1
XFILLER_112_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12966__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07695_ datapath.rf.registers\[8\]\[17\] net696 net666 datapath.rf.registers\[15\]\[17\]
+ _02530_ vssd1 vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__a221o_1
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09434_ _04264_ _04265_ _04268_ _04269_ vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__or4_1
X_06646_ mmio.key_data\[6\] net1049 _01484_ vssd1 vssd1 vccd1 vccd1 _01485_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10843__A2 _04177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08249__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09365_ _03613_ _04200_ vssd1 vssd1 vccd1 vccd1 _04201_ sky130_fd_sc_hd__nand2_1
XFILLER_40_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout522_A _05723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12267__A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06577_ datapath.PC\[30\] vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__inv_2
XANTENNA__08464__B net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08316_ datapath.rf.registers\[17\]\[4\] _01800_ net907 vssd1 vssd1 vccd1 vccd1 _03152_
+ sky130_fd_sc_hd__and3_1
XANTENNA__11602__C _05778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09296_ net459 _04130_ _04131_ vssd1 vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_10_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout310_X net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08247_ datapath.rf.registers\[3\]\[5\] net983 net927 vssd1 vssd1 vccd1 vccd1 _03083_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout408_X net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12348__A2 _06254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08178_ datapath.rf.registers\[3\]\[7\] net772 net764 datapath.rf.registers\[1\]\[7\]
+ _03011_ vssd1 vssd1 vccd1 vccd1 _03014_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout891_A net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07129_ datapath.rf.registers\[1\]\[28\] net847 net838 datapath.rf.registers\[26\]\[28\]
+ _01959_ vssd1 vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__a221o_1
XANTENNA__08421__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11110__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10140_ net226 _04975_ net1295 vssd1 vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__a21o_1
XANTENNA__07775__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_04_1297 vssd1 vssd1 vccd1 vccd1 team_04_1297/HI gpio_oeb[2] sky130_fd_sc_hd__conb_1
XANTENNA_fanout777_X net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10071_ _04903_ _04906_ vssd1 vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__xnor2_1
XFILLER_102_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout944_X net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13037__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13830_ clknet_leaf_113_clk _00639_ net1197 vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__dfrtp_1
X_13761_ clknet_leaf_76_clk _00570_ net1248 vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07262__C net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10973_ net1671 net298 net434 vssd1 vssd1 vccd1 vccd1 _00038_ sky130_fd_sc_hd__mux2_1
XANTENNA__12876__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11780__S _05894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12712_ _05894_ _06536_ _06537_ vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__and3b_1
X_13692_ clknet_leaf_10_clk _00502_ net1073 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07160__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12643_ _06476_ _06478_ vssd1 vssd1 vccd1 vccd1 _06483_ sky130_fd_sc_hd__nor2_1
XANTENNA__10249__X _05085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12574_ _06422_ _06423_ _06420_ vssd1 vssd1 vccd1 vccd1 _06425_ sky130_fd_sc_hd__o21a_1
X_14313_ clknet_leaf_20_clk _01018_ net1165 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11525_ screen.counter.ct\[3\] screen.counter.ct\[2\] vssd1 vssd1 vccd1 vccd1 _05749_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_129_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14244_ clknet_leaf_123_clk datapath.multiplication_module.multiplier_i_n\[12\] net1215
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_7_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11456_ net2409 net265 net409 vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__mux2_1
XANTENNA__06903__A _01630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10407_ _03420_ _03548_ vssd1 vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__xor2_1
X_14175_ clknet_leaf_47_clk _00930_ net1174 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08412__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11387_ net2104 net273 net412 vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__mux2_1
XANTENNA__11020__S net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07766__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13126_ net169 net2652 net473 vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__mux2_1
X_10338_ _05172_ _05173_ net228 _05171_ vssd1 vssd1 vccd1 vccd1 _05174_ sky130_fd_sc_hd__o211a_1
X_13057_ net176 net1624 net474 vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__mux2_1
X_10269_ net228 _05100_ _05104_ net1294 vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__a31o_1
XANTENNA__07518__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12008_ screen.register.currentXbus\[1\] _05755_ _05757_ screen.register.currentYbus\[25\]
+ _06051_ vssd1 vssd1 vccd1 vccd1 _06052_ sky130_fd_sc_hd__a221o_1
XFILLER_94_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07923__C1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08549__B net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07453__B net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06995__D net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12786__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13959_ clknet_leaf_109_clk _00737_ net1221 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_47_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07480_ datapath.rf.registers\[22\]\[21\] net734 net668 datapath.rf.registers\[21\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__a22o_1
XANTENNA__10825__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07151__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09150_ _02217_ net563 net442 vssd1 vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__mux2_1
X_08101_ _02913_ _02936_ vssd1 vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__nor2_1
X_09081_ _03499_ _03588_ _03497_ vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_79_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08032_ datapath.rf.registers\[6\]\[10\] net681 net662 datapath.rf.registers\[5\]\[10\]
+ _02866_ vssd1 vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_96_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold801 datapath.rf.registers\[27\]\[20\] vssd1 vssd1 vccd1 vccd1 net2149 sky130_fd_sc_hd__dlygate4sd3_1
Xhold812 datapath.rf.registers\[25\]\[13\] vssd1 vssd1 vccd1 vccd1 net2160 sky130_fd_sc_hd__dlygate4sd3_1
Xhold823 datapath.rf.registers\[8\]\[22\] vssd1 vssd1 vccd1 vccd1 net2171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold834 datapath.rf.registers\[22\]\[4\] vssd1 vssd1 vccd1 vccd1 net2182 sky130_fd_sc_hd__dlygate4sd3_1
Xhold845 datapath.rf.registers\[10\]\[22\] vssd1 vssd1 vccd1 vccd1 net2193 sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 datapath.rf.registers\[16\]\[0\] vssd1 vssd1 vccd1 vccd1 net2204 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold867 datapath.rf.registers\[17\]\[6\] vssd1 vssd1 vccd1 vccd1 net2215 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold878 datapath.rf.registers\[31\]\[8\] vssd1 vssd1 vccd1 vccd1 net2226 sky130_fd_sc_hd__dlygate4sd3_1
X_09983_ datapath.PC\[23\] net595 vssd1 vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__xor2_1
Xhold889 datapath.rf.registers\[19\]\[13\] vssd1 vssd1 vccd1 vccd1 net2237 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08934_ net649 _03642_ _03641_ vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__a21oi_4
X_08865_ _02613_ _02661_ net444 vssd1 vssd1 vccd1 vccd1 _03701_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout472_A net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08459__B _03294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08182__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07816_ datapath.rf.registers\[8\]\[14\] net877 net873 _02643_ _02651_ vssd1 vssd1
+ vccd1 vccd1 _02652_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07363__B net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08796_ _03617_ _03631_ net368 vssd1 vssd1 vccd1 vccd1 _03632_ sky130_fd_sc_hd__mux2_1
XANTENNA__07390__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07747_ datapath.rf.registers\[10\]\[16\] net706 net691 datapath.rf.registers\[13\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_154_Right_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_140_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10816__A2 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07142__B1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07678_ datapath.rf.registers\[11\]\[17\] net883 net843 datapath.rf.registers\[25\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13362__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09417_ net359 _04244_ _04250_ net345 vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__a31oi_1
X_06629_ net1287 net1282 datapath.ru.latched_instruction\[8\] mmio.memload_or_instruction\[8\]
+ vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__or4b_1
XFILLER_80_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout904_A _01620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08890__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout525_X net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09348_ net349 _04102_ _04103_ vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_43_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09279_ net905 _04085_ _04114_ vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__a21oi_1
X_11310_ net2090 net260 net417 vssd1 vssd1 vccd1 vccd1 _00355_ sky130_fd_sc_hd__mux2_1
X_12290_ _06272_ _06273_ net2617 net308 vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_107_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11241_ _05700_ net1621 net421 vssd1 vssd1 vccd1 vccd1 _00290_ sky130_fd_sc_hd__mux2_1
XFILLER_134_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12163__C net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07748__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08945__A1 _02311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11172_ net171 net2144 net531 vssd1 vssd1 vccd1 vccd1 _00225_ sky130_fd_sc_hd__mux2_1
X_10123_ _03729_ _04958_ _04956_ vssd1 vssd1 vccd1 vccd1 _04959_ sky130_fd_sc_hd__o21ba_1
XFILLER_79_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07825__Y _02661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13748__RESET_B net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input33_A DAT_I[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10054_ _04826_ _04887_ _04720_ vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__o21a_1
XANTENNA__11701__B1 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07273__B net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13813_ clknet_leaf_98_clk _00622_ net1230 vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__dfrtp_1
XFILLER_29_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_121_Right_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13744_ clknet_leaf_50_clk _00554_ net1181 vssd1 vssd1 vccd1 vccd1 mmio.key_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10956_ _01641_ _05516_ vssd1 vssd1 vccd1 vccd1 _05694_ sky130_fd_sc_hd__or2_2
XFILLER_44_774 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07133__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13675_ clknet_leaf_47_clk _00485_ net1171 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10887_ net211 net2447 net542 vssd1 vssd1 vccd1 vccd1 _00024_ sky130_fd_sc_hd__mux2_1
XFILLER_43_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11015__S net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12626_ _06461_ _06465_ _06468_ vssd1 vssd1 vccd1 vccd1 _06469_ sky130_fd_sc_hd__a21o_1
XFILLER_156_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12557_ datapath.mulitply_result\[8\] datapath.multiplication_module.multiplicand_i\[8\]
+ vssd1 vssd1 vccd1 vccd1 _06411_ sky130_fd_sc_hd__nor2_1
XANTENNA__08391__Y _03227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07288__X _02124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11508_ net175 net2283 net512 vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__mux2_1
X_12488_ net272 net1706 net507 vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__mux2_1
Xhold108 net44 vssd1 vssd1 vccd1 vccd1 net1456 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_156_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08551__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14227_ clknet_leaf_42_clk _00948_ net1144 vssd1 vssd1 vccd1 vccd1 columns.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold119 datapath.multiplication_module.multiplier_i\[7\] vssd1 vssd1 vccd1 vccd1
+ net1467 sky130_fd_sc_hd__dlygate4sd3_1
X_11439_ net182 net2296 net515 vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__mux2_1
XFILLER_125_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07739__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08936__A1 _01889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14158_ clknet_leaf_67_clk _00913_ net1239 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06920__X _01756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13109_ net251 net2517 net470 vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__mux2_1
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14089_ clknet_leaf_97_clk _00855_ net1226 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_06980_ net992 _01636_ _01647_ _01666_ vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__and4_2
XANTENNA__12370__A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1170 net1186 vssd1 vssd1 vccd1 vccd1 net1170 sky130_fd_sc_hd__clkbuf_2
Xfanout1181 net1182 vssd1 vssd1 vccd1 vccd1 net1181 sky130_fd_sc_hd__clkbuf_4
X_08650_ _01980_ _02003_ vssd1 vssd1 vccd1 vccd1 _03486_ sky130_fd_sc_hd__or2_1
Xfanout1192 net1194 vssd1 vssd1 vccd1 vccd1 net1192 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07372__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07751__X _02587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07911__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07601_ _02434_ _02435_ _02436_ vssd1 vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__nor3_1
XFILLER_19_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08581_ datapath.rf.registers\[0\]\[0\] net783 _03401_ _03416_ vssd1 vssd1 vccd1
+ vccd1 _03417_ sky130_fd_sc_hd__o22a_4
XANTENNA__09649__C1 _03613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_105_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07532_ datapath.rf.registers\[26\]\[20\] net778 net675 datapath.rf.registers\[29\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_105_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07463_ net872 _02296_ _02297_ _02298_ vssd1 vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__or4_1
XANTENNA__08872__A0 _03009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09202_ net551 net547 _02311_ vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_22_Left_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07394_ datapath.rf.registers\[22\]\[23\] net734 net718 datapath.rf.registers\[20\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__a22o_1
X_09133_ net647 _03968_ _03770_ vssd1 vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__o21a_1
XANTENNA__10764__S net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13140__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07978__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09064_ net338 _03899_ vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__nor2_1
XANTENNA__12264__B net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08015_ datapath.rf.registers\[24\]\[10\] net858 net851 datapath.rf.registers\[17\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__a22o_1
Xhold620 datapath.rf.registers\[0\]\[4\] vssd1 vssd1 vccd1 vccd1 net1968 sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 datapath.rf.registers\[20\]\[5\] vssd1 vssd1 vccd1 vccd1 net1979 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold642 datapath.rf.registers\[6\]\[19\] vssd1 vssd1 vccd1 vccd1 net1990 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1227_A net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08927__A1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold653 datapath.rf.registers\[13\]\[11\] vssd1 vssd1 vccd1 vccd1 net2001 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold664 datapath.rf.registers\[9\]\[29\] vssd1 vssd1 vccd1 vccd1 net2012 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06830__X _01666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06938__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold675 datapath.rf.registers\[28\]\[17\] vssd1 vssd1 vccd1 vccd1 net2023 sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 datapath.rf.registers\[31\]\[24\] vssd1 vssd1 vccd1 vccd1 net2034 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold697 datapath.rf.registers\[10\]\[16\] vssd1 vssd1 vccd1 vccd1 net2045 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout687_A net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09966_ _04757_ _04801_ vssd1 vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_31_Left_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08917_ datapath.PC\[31\] _03752_ net1038 vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11608__B _05786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09897_ datapath.PC\[18\] _04731_ vssd1 vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__xor2_2
XANTENNA__07805__C net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_96_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_96_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout475_X net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout854_A net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08155__A2 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08848_ _03229_ _01647_ _03671_ vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__mux2_1
XANTENNA__07902__A2 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08779_ net648 net555 _03613_ vssd1 vssd1 vccd1 vccd1 _03615_ sky130_fd_sc_hd__and3_2
XANTENNA_fanout642_X net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10810_ datapath.mulitply_result\[11\] net598 net620 vssd1 vssd1 vccd1 vccd1 _05569_
+ sky130_fd_sc_hd__a21o_1
X_11790_ _01670_ _05901_ _05899_ vssd1 vssd1 vccd1 vccd1 _05902_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07115__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10741_ net1504 net568 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[27\]
+ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_40_Left_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout907_X net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13460_ clknet_leaf_93_clk _00270_ net1210 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10672_ button\[2\] net1022 vssd1 vssd1 vccd1 vccd1 _05490_ sky130_fd_sc_hd__nand2_1
X_12411_ _05968_ net158 vssd1 vssd1 vccd1 vccd1 _06353_ sky130_fd_sc_hd__nor2_1
X_13391_ clknet_leaf_23_clk _00201_ net1134 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_138_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13050__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_20_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_8
X_12342_ net641 _03950_ net309 vssd1 vssd1 vccd1 vccd1 _06311_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_153_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12273_ net892 _04454_ _06259_ _06260_ vssd1 vssd1 vccd1 vccd1 _06261_ sky130_fd_sc_hd__o22a_1
XANTENNA__07268__B net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_12_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14012_ clknet_leaf_68_clk _00781_ net1249 vssd1 vssd1 vccd1 vccd1 datapath.PC\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11224_ net245 net2410 net526 vssd1 vssd1 vccd1 vccd1 _00274_ sky130_fd_sc_hd__mux2_1
XANTENNA__06740__X _01579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10725__A1 _02804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11155_ net253 net2156 net531 vssd1 vssd1 vccd1 vccd1 _00208_ sky130_fd_sc_hd__mux2_1
XFILLER_122_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10106_ _04892_ _04941_ net229 vssd1 vssd1 vccd1 vccd1 _04942_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11086_ net254 net1804 net534 vssd1 vssd1 vccd1 vccd1 _00143_ sky130_fd_sc_hd__mux2_1
XFILLER_76_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_87_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08099__B _01784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10037_ _04868_ _04869_ _04871_ vssd1 vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__or3b_1
XFILLER_64_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07354__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07290__Y _02126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07106__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11988_ screen.register.currentXbus\[16\] _05769_ _05837_ screen.register.currentYbus\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06033_ sky130_fd_sc_hd__a22o_1
XANTENNA__11989__B1 _06018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09004__A _01888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13727_ clknet_leaf_12_clk _00537_ net1082 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08854__A0 _02419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10939_ datapath.PC\[30\] _05671_ vssd1 vssd1 vccd1 vccd1 _05679_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_27_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13658_ clknet_leaf_2_clk _00468_ net1065 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12609_ _06446_ _06453_ _06452_ _06451_ vssd1 vssd1 vccd1 vccd1 _06455_ sky130_fd_sc_hd__o211ai_1
X_13589_ clknet_leaf_19_clk _00399_ net1116 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_145_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_11_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08562__B net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10716__A1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout407 _05733_ vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__buf_4
X_09820_ net341 _04616_ vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__nand2_1
XANTENNA__08385__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout418 _05722_ vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__clkbuf_8
XFILLER_113_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout429 _05716_ vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__buf_4
XANTENNA__07593__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09751_ _03451_ _03513_ vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__xnor2_1
X_06963_ net965 net911 net908 vssd1 vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_78_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09334__A1 _02567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08137__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08702_ _02912_ _02936_ vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_107_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10900__X _05646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09682_ _03537_ _03538_ vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__and2_1
XANTENNA__07345__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06894_ _01712_ net929 vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__and2_1
X_08633_ _02094_ _03462_ _03463_ _03465_ _02093_ vssd1 vssd1 vccd1 vccd1 _03469_ sky130_fd_sc_hd__a41o_1
XANTENNA__06699__A2 _01502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13135__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout268_A net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08564_ datapath.rf.registers\[26\]\[0\] net781 _03397_ _03398_ _03399_ vssd1 vssd1
+ vccd1 vccd1 _03400_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_120_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07515_ datapath.rf.registers\[24\]\[20\] net856 _02337_ _02348_ _02349_ vssd1 vssd1
+ vccd1 vccd1 _02351_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07360__C net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08845__A0 _02126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12974__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08495_ datapath.rf.registers\[8\]\[1\] net970 net912 _01793_ vssd1 vssd1 vccd1 vccd1
+ _03331_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout435_A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1177_A net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07446_ _02276_ _02278_ _02280_ _02281_ vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__or4_1
XANTENNA__09849__A net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07377_ datapath.rf.registers\[11\]\[23\] net882 net832 datapath.rf.registers\[30\]\[23\]
+ _02212_ vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__a221o_1
XANTENNA__12275__A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09116_ _03460_ _03951_ vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_135_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06704__C datapath.ru.latched_instruction\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09047_ _03881_ _03882_ vssd1 vssd1 vccd1 vccd1 _03883_ sky130_fd_sc_hd__nor2_1
XFILLER_117_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold450 datapath.rf.registers\[22\]\[10\] vssd1 vssd1 vccd1 vccd1 net1798 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10707__A1 _02771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold461 datapath.rf.registers\[13\]\[4\] vssd1 vssd1 vccd1 vccd1 net1809 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold472 datapath.rf.registers\[11\]\[5\] vssd1 vssd1 vccd1 vccd1 net1820 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08376__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold483 datapath.rf.registers\[8\]\[1\] vssd1 vssd1 vccd1 vccd1 net1831 sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 datapath.rf.registers\[1\]\[6\] vssd1 vssd1 vccd1 vccd1 net1842 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_78 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06720__B _01443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07584__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout930 _01727_ vssd1 vssd1 vccd1 vccd1 net930 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout941 net942 vssd1 vssd1 vccd1 vccd1 net941 sky130_fd_sc_hd__clkbuf_4
X_09949_ _01416_ _03265_ vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__nand2_1
Xfanout952 net953 vssd1 vssd1 vccd1 vccd1 net952 sky130_fd_sc_hd__buf_2
Xfanout963 net965 vssd1 vssd1 vccd1 vccd1 net963 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout857_X net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_69_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_58_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09325__A1 _02522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout974 net975 vssd1 vssd1 vccd1 vccd1 net974 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08128__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout985 net986 vssd1 vssd1 vccd1 vccd1 net985 sky130_fd_sc_hd__clkbuf_2
Xfanout996 _05790_ vssd1 vssd1 vccd1 vccd1 net996 sky130_fd_sc_hd__buf_2
X_12960_ net168 net2641 net395 vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_51_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1150 datapath.rf.registers\[12\]\[9\] vssd1 vssd1 vccd1 vccd1 net2498 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07336__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09876__A2 _04710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1161 datapath.mulitply_result\[17\] vssd1 vssd1 vccd1 vccd1 net2509 sky130_fd_sc_hd__dlygate4sd3_1
X_11911_ screen.register.currentYbus\[18\] net162 vssd1 vssd1 vccd1 vccd1 _05971_
+ sky130_fd_sc_hd__nand2_1
XFILLER_100_782 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1172 datapath.rf.registers\[0\]\[20\] vssd1 vssd1 vccd1 vccd1 net2520 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1183 datapath.mulitply_result\[18\] vssd1 vssd1 vccd1 vccd1 net2531 sky130_fd_sc_hd__dlygate4sd3_1
X_12891_ net176 net1897 net401 vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__mux2_1
Xhold1194 datapath.mulitply_result\[2\] vssd1 vssd1 vccd1 vccd1 net2542 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13045__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14630_ clknet_leaf_11_clk _01335_ net1083 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11842_ _05760_ _05804_ _05909_ _05920_ vssd1 vssd1 vccd1 vccd1 _05921_ sky130_fd_sc_hd__or4_1
XANTENNA__09089__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14561_ clknet_leaf_37_clk _01266_ net1147 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12884__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11773_ net1391 net144 net139 vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__a21o_1
XANTENNA__07270__C net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08934__Y _03770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08300__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13512_ clknet_leaf_91_clk _00322_ net1233 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10724_ net1963 _02856_ net572 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[10\]
+ sky130_fd_sc_hd__mux2_1
X_14492_ clknet_leaf_9_clk _01197_ net1074 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08663__A _02217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09111__X _03947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13443_ clknet_leaf_119_clk _00253_ net1191 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10655_ _05437_ _05472_ _05466_ vssd1 vssd1 vccd1 vccd1 _05474_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06862__A2 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13374_ clknet_leaf_148_clk _00184_ net1062 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload17 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 clkload17/Y sky130_fd_sc_hd__clkinv_4
XFILLER_139_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10586_ _03227_ _03292_ _03357_ _03417_ vssd1 vssd1 vccd1 vccd1 _05409_ sky130_fd_sc_hd__or4_1
Xclkload28 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 clkload28/X sky130_fd_sc_hd__clkbuf_8
Xclkload39 clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 clkload39/X sky130_fd_sc_hd__clkbuf_4
X_12325_ datapath.PC\[19\] _06298_ net306 vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__mux2_1
XFILLER_154_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09494__A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12256_ net310 vssd1 vssd1 vccd1 vccd1 _06247_ sky130_fd_sc_hd__inv_2
XANTENNA__09013__B1 _03770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11207_ _05517_ _05720_ vssd1 vssd1 vccd1 vccd1 _05721_ sky130_fd_sc_hd__nand2_4
X_12187_ screen.counter.ct\[21\] _06152_ _06166_ vssd1 vssd1 vccd1 vccd1 _06203_ sky130_fd_sc_hd__and3b_1
XANTENNA__07575__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11138_ net169 net2189 net426 vssd1 vssd1 vccd1 vccd1 _00193_ sky130_fd_sc_hd__mux2_1
XFILLER_122_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09316__A1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08119__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11069_ net169 net2546 net430 vssd1 vssd1 vccd1 vccd1 _00129_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_0_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07327__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08838__A _03669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08827__A0 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12794__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14759_ screen.screenLogic.currentWrx vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__clkbuf_1
X_07300_ datapath.rf.registers\[10\]\[25\] net708 net693 datapath.rf.registers\[13\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_22_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08280_ datapath.rf.registers\[9\]\[5\] net703 net684 datapath.rf.registers\[27\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_82_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07231_ datapath.rf.registers\[16\]\[26\] net860 net853 datapath.rf.registers\[19\]\[26\]
+ _02066_ vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__a221o_1
XANTENNA__11203__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07162_ datapath.rf.registers\[6\]\[28\] net682 net667 datapath.rf.registers\[15\]\[28\]
+ _01997_ vssd1 vssd1 vccd1 vccd1 _01998_ sky130_fd_sc_hd__a221o_1
XFILLER_118_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07093_ datapath.rf.registers\[30\]\[29\] net833 _01927_ _01928_ vssd1 vssd1 vccd1
+ vccd1 _01929_ sky130_fd_sc_hd__a211o_1
XANTENNA__08358__A2 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_130_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout204 _05641_ vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_130_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout215 net217 vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__clkbuf_2
Xfanout226 _04713_ vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__buf_2
Xfanout237 _05616_ vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__clkbuf_2
X_09803_ _03483_ net628 net624 _03484_ net645 vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__a221o_1
Xfanout248 net250 vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__clkbuf_2
Xfanout259 net261 vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12969__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07995_ datapath.rf.registers\[12\]\[10\] net955 net920 vssd1 vssd1 vccd1 vccd1 _02831_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09307__A1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09734_ net326 _03776_ _04568_ _04569_ vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__a2bb2o_1
XPHY_EDGE_ROW_105_Left_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06946_ MemWrite _01780_ vssd1 vssd1 vccd1 vccd1 _01782_ sky130_fd_sc_hd__or2_1
XANTENNA__07318__B1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12311__B1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09665_ _04499_ _04500_ net325 _03932_ vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_28_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06877_ net985 net949 vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__and2_2
XANTENNA_fanout1294_A _01436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08467__B net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14292__RESET_B net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08616_ _02491_ _02545_ _03449_ _03450_ _02489_ vssd1 vssd1 vccd1 vccd1 _03452_ sky130_fd_sc_hd__a41o_1
XANTENNA__08530__A2 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10873__B1 _05621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09596_ net455 _04280_ _04431_ vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__a21o_1
XFILLER_70_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08547_ datapath.rf.registers\[0\]\[0\] net869 _03369_ _03382_ vssd1 vssd1 vccd1
+ vccd1 _03383_ sky130_fd_sc_hd__o22ai_4
XANTENNA_fanout817_A net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12090__A2 _05786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08478_ datapath.rf.registers\[4\]\[1\] net865 net823 datapath.rf.registers\[22\]\[1\]
+ _03301_ vssd1 vssd1 vccd1 vccd1 _03314_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_137_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07429_ datapath.rf.registers\[25\]\[22\] net726 net668 datapath.rf.registers\[21\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_114_Left_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout605_X net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11113__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_922 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10440_ net1269 datapath.PC\[3\] vssd1 vssd1 vccd1 vccd1 _05276_ sky130_fd_sc_hd__xor2_1
XANTENNA__10928__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10237__B _05052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10371_ net466 _04395_ _05206_ net1044 vssd1 vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__a211o_1
XFILLER_152_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12110_ screen.counter.currentCt\[13\] screen.counter.currentCt\[12\] screen.counter.currentCt\[15\]
+ screen.counter.currentCt\[14\] vssd1 vssd1 vccd1 vccd1 _06147_ sky130_fd_sc_hd__or4_1
XFILLER_2_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13090_ net2107 net176 net388 vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__mux2_1
XFILLER_6_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout974_X net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12041_ screen.register.currentYbus\[19\] _05773_ net997 screen.register.currentXbus\[19\]
+ _06082_ vssd1 vssd1 vccd1 vccd1 _06083_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_53_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold280 datapath.rf.registers\[31\]\[30\] vssd1 vssd1 vccd1 vccd1 net1628 sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 datapath.rf.registers\[9\]\[20\] vssd1 vssd1 vccd1 vccd1 net1639 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_120_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_123_Left_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12879__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07265__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout760 _01802_ vssd1 vssd1 vccd1 vccd1 net760 sky130_fd_sc_hd__buf_4
Xfanout771 net773 vssd1 vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_148_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout782 net785 vssd1 vssd1 vccd1 vccd1 net782 sky130_fd_sc_hd__buf_6
XANTENNA__10540__X _05368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13992_ clknet_leaf_112_clk _00769_ net1218 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout793 net795 vssd1 vssd1 vccd1 vccd1 net793 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07309__B1 _02139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08658__A _02126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12943_ net251 net2606 net394 vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__mux2_1
XANTENNA__08521__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_64_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12874_ net269 datapath.rf.registers\[2\]\[11\] net400 vssd1 vssd1 vccd1 vccd1 _01124_
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11825_ _01477_ net1017 net315 net335 datapath.ru.latched_instruction\[31\] vssd1
+ vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__a32o_1
X_14613_ clknet_leaf_18_clk _01318_ net1108 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_14544_ clknet_leaf_23_clk _01249_ net1155 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07088__A2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11756_ net1507 net143 net138 _02587_ vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__a22o_1
XANTENNA__12081__A2 _05778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08393__A _03228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_79_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10707_ net1465 _02771_ net571 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i_n\[12\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14475_ clknet_leaf_55_clk _01180_ net1173 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11687_ _05008_ net152 net148 net1422 vssd1 vssd1 vccd1 vccd1 _00572_ sky130_fd_sc_hd__a22o_1
XANTENNA__11023__S net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_122_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap1000 _05755_ vssd1 vssd1 vccd1 vccd1 net1000 sky130_fd_sc_hd__clkbuf_2
X_13426_ clknet_leaf_30_clk _00236_ net1124 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10638_ _05449_ _05451_ vssd1 vssd1 vccd1 vccd1 _05458_ sky130_fd_sc_hd__nor2_1
Xclkload106 clknet_leaf_126_clk vssd1 vssd1 vccd1 vccd1 clkload106/Y sky130_fd_sc_hd__inv_8
Xclkload117 clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 clkload117/Y sky130_fd_sc_hd__inv_6
Xclkload128 clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 clkload128/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__09785__A1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08588__A2 _03423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload139 clknet_leaf_86_clk vssd1 vssd1 vccd1 vccd1 clkload139/Y sky130_fd_sc_hd__clkinv_4
X_13357_ clknet_leaf_132_clk _00167_ net1100 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10569_ _05389_ _05390_ _05392_ vssd1 vssd1 vccd1 vccd1 _05393_ sky130_fd_sc_hd__or3_1
X_12308_ datapath.PC\[14\] _06246_ _06286_ vssd1 vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__a21o_1
XFILLER_5_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13288_ clknet_leaf_91_clk _00098_ net1232 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_137_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07456__B _01717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12239_ net1511 _06233_ _06235_ vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__a21oi_1
XFILLER_69_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_17_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07012__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12789__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06800_ net1004 net1020 _01634_ _01633_ vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__a31oi_4
XFILLER_96_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07780_ datapath.rf.registers\[16\]\[15\] net739 net723 datapath.rf.registers\[18\]\[15\]
+ _02615_ vssd1 vssd1 vccd1 vccd1 _02616_ sky130_fd_sc_hd__a221o_1
Xinput4 DAT_I[11] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
X_06731_ datapath.ru.latched_instruction\[4\] net1026 vssd1 vssd1 vccd1 vccd1 _01570_
+ sky130_fd_sc_hd__and2_1
XANTENNA__11706__B net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10304__C1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09450_ net648 _04285_ net438 vssd1 vssd1 vccd1 vccd1 _04286_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_84_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06662_ _01408_ _01500_ vssd1 vssd1 vccd1 vccd1 _01501_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_84_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09715__A2_N net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07720__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08401_ datapath.rf.registers\[7\]\[2\] net942 net936 vssd1 vssd1 vccd1 vccd1 _03237_
+ sky130_fd_sc_hd__and3_1
X_09381_ net458 _04161_ _04216_ vssd1 vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__a21o_1
X_06593_ columns.count\[5\] columns.count\[4\] vssd1 vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__nor2_1
XANTENNA__12377__X _06335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08332_ datapath.rf.registers\[16\]\[4\] net738 net672 datapath.rf.registers\[7\]\[4\]
+ _03157_ vssd1 vssd1 vccd1 vccd1 _03168_ sky130_fd_sc_hd__a221o_1
XANTENNA__07079__A2 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08263_ datapath.rf.registers\[1\]\[5\] net846 net817 datapath.rf.registers\[7\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03099_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_4_0_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07214_ datapath.rf.registers\[17\]\[26\] net849 net826 datapath.rf.registers\[12\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02050_ sky130_fd_sc_hd__a22o_1
X_08194_ _03028_ _03029_ net611 vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08579__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07145_ _01970_ _01979_ _01415_ net874 vssd1 vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__a2bb2o_4
XFILLER_134_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10772__S net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07787__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07251__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07076_ _01911_ vssd1 vssd1 vccd1 vccd1 _01912_ sky130_fd_sc_hd__inv_2
XANTENNA__08242__S net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12272__B _06254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09528__A1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07539__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout767_A net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout388_X net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14473__RESET_B net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07978_ datapath.rf.registers\[17\]\[11\] net748 net677 datapath.rf.registers\[29\]\[11\]
+ _02813_ vssd1 vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__a221o_1
XFILLER_74_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07382__A _02217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09717_ _04010_ _04016_ net340 vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__mux2_1
X_06929_ net981 net917 vssd1 vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__and2_2
XANTENNA_fanout555_X net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout934_A net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11108__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09648_ net327 _04198_ _04482_ _04483_ net379 vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__a221o_1
XFILLER_83_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08765__X _03601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10310__A2 net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout722_X net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09579_ _04162_ _04413_ net354 vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__mux2_1
XANTENNA__10947__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08484__Y _03320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11610_ net1010 _05794_ vssd1 vssd1 vccd1 vccd1 _05834_ sky130_fd_sc_hd__nand2_1
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12590_ _06435_ _06438_ vssd1 vssd1 vccd1 vccd1 _06439_ sky130_fd_sc_hd__xor2_1
XFILLER_143_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11541_ _05293_ _05753_ vssd1 vssd1 vccd1 vccd1 _05765_ sky130_fd_sc_hd__or2_1
XANTENNA__06817__A2 _01575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14260_ clknet_leaf_127_clk _00965_ net1209 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11472_ net1957 net176 net408 vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__mux2_1
XANTENNA__08941__A net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11778__S _05894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13211_ clknet_leaf_37_clk _00021_ net1138 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10423_ net366 _04323_ _05258_ vssd1 vssd1 vccd1 vccd1 _05259_ sky130_fd_sc_hd__o21a_1
X_14191_ clknet_leaf_90_clk datapath.multiplication_module.multiplicand_i_n\[2\] net1241
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__06732__Y _01571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07778__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08660__B _02190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13142_ net2178 _05588_ net382 vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__mux2_1
XANTENNA__07242__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10354_ _05189_ net891 _04517_ vssd1 vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__or3b_1
XFILLER_136_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12182__B net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13073_ net2129 net266 net388 vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__mux2_1
XFILLER_112_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10285_ net1038 _05118_ _05120_ net639 vssd1 vssd1 vccd1 vccd1 _05121_ sky130_fd_sc_hd__a211o_1
XFILLER_111_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07844__X _02680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12024_ screen.register.currentXbus\[26\] _05772_ _05837_ screen.register.currentYbus\[18\]
+ _06066_ vssd1 vssd1 vccd1 vccd1 _06067_ sky130_fd_sc_hd__a221o_1
XFILLER_78_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10711__A net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13975_ clknet_leaf_105_clk _00753_ net1224 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[18\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__11018__S net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10837__B1 _05590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload9_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12926_ net1775 net173 net484 vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07702__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12857_ net185 net1828 net487 vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__mux2_1
XFILLER_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08835__B net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11808_ net2360 net1051 net315 net335 datapath.ru.latched_instruction\[14\] vssd1
+ vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__a32o_1
XANTENNA__12054__A2 _05786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12788_ net199 net2036 net495 vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__mux2_1
X_11739_ datapath.ru.n_memwrite _05289_ _05291_ vssd1 vssd1 vccd1 vccd1 _05891_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_32_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14527_ clknet_leaf_13_clk _01232_ net1076 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11801__A2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07481__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14458_ clknet_leaf_3_clk _01163_ net1076 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_13409_ clknet_leaf_45_clk _00219_ net1147 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_14389_ clknet_leaf_130_clk _01094_ net1111 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10445__X _05281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07769__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07233__A2 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08950_ _03783_ _03784_ net450 vssd1 vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__mux2_1
XFILLER_142_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07901_ datapath.rf.registers\[17\]\[12\] net852 _02728_ _02729_ _02730_ vssd1 vssd1
+ vccd1 vccd1 _02737_ sky130_fd_sc_hd__a2111o_1
X_08881_ _01610_ _03716_ vssd1 vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_135_Right_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08194__A0 _03028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07832_ datapath.rf.registers\[19\]\[14\] net731 net727 datapath.rf.registers\[25\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__a22o_1
XFILLER_111_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06744__A1 _01502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07763_ _02595_ _02596_ _02598_ vssd1 vssd1 vccd1 vccd1 _02599_ sky130_fd_sc_hd__or3_1
X_09502_ _04333_ _04335_ _04337_ _04302_ vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__o31a_2
X_06714_ mmio.memload_or_instruction\[7\] mmio.memload_or_instruction\[9\] vssd1 vssd1
+ vccd1 vccd1 _01553_ sky130_fd_sc_hd__nand2_1
XFILLER_65_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07694_ datapath.rf.registers\[19\]\[17\] net732 net712 datapath.rf.registers\[11\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__a22o_1
X_09433_ _03526_ net626 net625 _03525_ net643 vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__a221o_1
X_06645_ net1290 net1285 mmio.memload_or_instruction\[6\] vssd1 vssd1 vccd1 vccd1
+ _01484_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout250_A _05592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13866__RESET_B net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13143__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09364_ _03634_ _04199_ net331 vssd1 vssd1 vccd1 vccd1 _04200_ sky130_fd_sc_hd__mux2_1
X_06576_ datapath.PC\[4\] vssd1 vssd1 vccd1 vccd1 _01417_ sky130_fd_sc_hd__inv_2
X_08315_ datapath.rf.registers\[30\]\[4\] net758 net750 datapath.rf.registers\[28\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__a22o_1
XANTENNA__08464__C net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09295_ net551 net547 _02522_ vssd1 vssd1 vccd1 vccd1 _04131_ sky130_fd_sc_hd__a21o_1
XANTENNA__12982__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout515_A _05731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1257_A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08246_ datapath.rf.registers\[0\]\[5\] net871 vssd1 vssd1 vccd1 vccd1 _03082_ sky130_fd_sc_hd__or2_1
XFILLER_21_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07472__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08177_ datapath.rf.registers\[2\]\[7\] net744 net666 datapath.rf.registers\[15\]\[7\]
+ _03012_ vssd1 vssd1 vccd1 vccd1 _03013_ sky130_fd_sc_hd__a221o_1
XFILLER_119_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12283__A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07128_ _01962_ _01963_ vssd1 vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__or2_1
XFILLER_137_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07224__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout884_A _01719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xteam_04_1298 vssd1 vssd1 vccd1 vccd1 team_04_1298/HI gpio_oeb[3] sky130_fd_sc_hd__conb_1
X_07059_ datapath.rf.registers\[2\]\[30\] net744 net685 datapath.rf.registers\[27\]\[30\]
+ _01894_ vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__a221o_1
XFILLER_88_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10070_ _04904_ _04905_ vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__xnor2_1
XFILLER_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout672_X net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_102_Right_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08185__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06735__A1 _01441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07932__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout937_X net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13760_ clknet_leaf_76_clk _00569_ net1248 vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__dfrtp_1
XFILLER_44_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10972_ net1705 net302 net436 vssd1 vssd1 vccd1 vccd1 _00037_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12711_ _01404_ _05892_ _01432_ vssd1 vssd1 vccd1 vccd1 _06537_ sky130_fd_sc_hd__or3b_1
X_13691_ clknet_leaf_45_clk _00501_ net1146 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13053__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08655__B _02091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12642_ datapath.mulitply_result\[22\] datapath.multiplication_module.multiplicand_i\[22\]
+ vssd1 vssd1 vccd1 vccd1 _06482_ sky130_fd_sc_hd__or2_1
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12177__B net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12892__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12573_ net2430 net504 net500 _06424_ vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__a22o_1
XFILLER_7_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09767__A _04084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11795__B2 _01502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11524_ net1280 screen.counter.ct\[5\] _05301_ vssd1 vssd1 vccd1 vccd1 _05748_ sky130_fd_sc_hd__or3_1
XFILLER_7_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14312_ clknet_leaf_61_clk _01017_ net1166 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_14243_ clknet_leaf_124_clk datapath.multiplication_module.multiplier_i_n\[11\] net1215
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_144_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11455_ net1692 net268 net408 vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__mux2_1
XFILLER_125_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11301__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10406_ net222 _05241_ vssd1 vssd1 vccd1 vccd1 _05242_ sky130_fd_sc_hd__and2_1
X_14174_ clknet_leaf_47_clk _00929_ net1174 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07215__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11386_ net2155 net274 net412 vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__mux2_1
XFILLER_152_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13125_ net173 net2039 net471 vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__mux2_1
X_10337_ net636 _04583_ vssd1 vssd1 vccd1 vccd1 _05173_ sky130_fd_sc_hd__nand2_1
XFILLER_125_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13056_ net185 net2205 net474 vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__mux2_1
X_10268_ net1043 _03739_ _05103_ _05102_ net899 vssd1 vssd1 vccd1 vccd1 _05104_ sky130_fd_sc_hd__a311o_1
XANTENNA__08176__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12007_ screen.register.currentXbus\[9\] _05768_ _06018_ screen.register.currentYbus\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06051_ sky130_fd_sc_hd__a22o_1
XFILLER_78_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10199_ net1265 _03746_ datapath.PC\[23\] vssd1 vssd1 vccd1 vccd1 _05035_ sky130_fd_sc_hd__o21a_1
XANTENNA__09007__A _01980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07453__C net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13958_ clknet_leaf_107_clk _00736_ net1223 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_17_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12909_ net2056 net254 net483 vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__mux2_1
XFILLER_62_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13889_ clknet_leaf_49_clk keypad.decode.button_n\[0\] net1176 vssd1 vssd1 vccd1
+ vccd1 button\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12368__A net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08100__A0 _02934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08100_ _02934_ _02935_ net611 vssd1 vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__mux2_1
X_09080_ _03868_ _03914_ vssd1 vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_79_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08031_ datapath.rf.registers\[30\]\[10\] net760 net752 datapath.rf.registers\[28\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__a22o_1
XFILLER_135_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold802 datapath.rf.registers\[28\]\[4\] vssd1 vssd1 vccd1 vccd1 net2150 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11211__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07206__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold813 datapath.mulitply_result\[15\] vssd1 vssd1 vccd1 vccd1 net2161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold824 datapath.rf.registers\[23\]\[20\] vssd1 vssd1 vccd1 vccd1 net2172 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09600__B1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold835 datapath.rf.registers\[24\]\[30\] vssd1 vssd1 vccd1 vccd1 net2183 sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 datapath.rf.registers\[18\]\[14\] vssd1 vssd1 vccd1 vccd1 net2194 sky130_fd_sc_hd__dlygate4sd3_1
Xhold857 datapath.rf.registers\[21\]\[27\] vssd1 vssd1 vccd1 vccd1 net2205 sky130_fd_sc_hd__dlygate4sd3_1
X_09982_ _04724_ _04817_ vssd1 vssd1 vccd1 vccd1 _04818_ sky130_fd_sc_hd__nor2_1
Xhold868 datapath.rf.registers\[7\]\[12\] vssd1 vssd1 vccd1 vccd1 net2216 sky130_fd_sc_hd__dlygate4sd3_1
Xhold879 datapath.rf.registers\[10\]\[27\] vssd1 vssd1 vccd1 vccd1 net2227 sky130_fd_sc_hd__dlygate4sd3_1
X_08933_ net330 _03768_ net311 vssd1 vssd1 vccd1 vccd1 _03769_ sky130_fd_sc_hd__a21o_1
XANTENNA__13138__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08864_ net317 vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_127_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07815_ _02642_ _02648_ _02649_ _02650_ vssd1 vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__or4_1
XANTENNA__12977__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07363__C net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08795_ _03419_ _03615_ _01779_ vssd1 vssd1 vccd1 vccd1 _03631_ sky130_fd_sc_hd__a21oi_1
X_07746_ _02580_ _02581_ vssd1 vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__or2_1
XFILLER_26_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12266__A2 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07677_ net874 _02510_ _02511_ _02512_ vssd1 vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout632_A net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09416_ _04041_ _04042_ net356 vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__o21ai_1
X_06628_ net1287 net1282 mmio.memload_or_instruction\[8\] vssd1 vssd1 vccd1 vccd1
+ _01467_ sky130_fd_sc_hd__or3b_2
XFILLER_53_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07693__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09347_ net607 _04180_ vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout420_X net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1162_X net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout518_X net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13657__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07445__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09278_ _03509_ net627 net624 _03508_ net644 vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__a221o_1
XFILLER_21_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08229_ datapath.rf.registers\[24\]\[6\] net766 _03064_ net786 vssd1 vssd1 vccd1
+ vccd1 _03065_ sky130_fd_sc_hd__a211o_1
XFILLER_153_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11121__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11240_ _05695_ _05708_ vssd1 vssd1 vccd1 vccd1 _05722_ sky130_fd_sc_hd__nand2_4
XANTENNA_fanout887_X net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11171_ net172 net1773 net531 vssd1 vssd1 vccd1 vccd1 _00224_ sky130_fd_sc_hd__mux2_1
XANTENNA__10960__S net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10122_ datapath.PC\[21\] _04057_ net469 vssd1 vssd1 vccd1 vccd1 _04958_ sky130_fd_sc_hd__mux2_1
XANTENNA__11690__A2_N _05885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08158__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13048__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10053_ _04885_ _04888_ vssd1 vssd1 vccd1 vccd1 _04889_ sky130_fd_sc_hd__or2_1
XFILLER_88_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input26_A DAT_I[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12887__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07273__C net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13788__RESET_B net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07381__B2 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13812_ clknet_leaf_98_clk _00621_ net1230 vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_3_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10268__A1 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13743_ clknet_leaf_49_clk _00553_ net1176 vssd1 vssd1 vccd1 vccd1 mmio.key_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10955_ _05513_ _05692_ vssd1 vssd1 vccd1 vccd1 _05693_ sky130_fd_sc_hd__nor2_1
XANTENNA__08330__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10886_ net1047 net652 _05632_ _05633_ vssd1 vssd1 vccd1 vccd1 _05634_ sky130_fd_sc_hd__o22a_4
X_13674_ clknet_leaf_59_clk _00484_ net1170 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_12625_ _06466_ _06467_ vssd1 vssd1 vccd1 vccd1 _06468_ sky130_fd_sc_hd__or2_1
XANTENNA__07436__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12556_ datapath.mulitply_result\[8\] datapath.multiplication_module.multiplicand_i\[8\]
+ vssd1 vssd1 vccd1 vccd1 _06410_ sky130_fd_sc_hd__and2_1
XFILLER_156_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11507_ net182 net2341 net511 vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__mux2_1
XANTENNA__10436__A _04338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12487_ net274 net1926 net507 vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__mux2_1
XANTENNA__11031__S net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold109 mmio.memload_or_instruction\[0\] vssd1 vssd1 vccd1 vccd1 net1457 sky130_fd_sc_hd__dlygate4sd3_1
X_14226_ clknet_leaf_42_clk _00947_ net1144 vssd1 vssd1 vccd1 vccd1 columns.count\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_11438_ net179 net1826 net517 vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__mux2_1
X_14157_ clknet_leaf_68_clk _00912_ net1239 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11369_ net195 net1574 net519 vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__mux2_1
XFILLER_98_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13108_ net255 net1969 net472 vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__mux2_1
XFILLER_140_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14088_ clknet_leaf_96_clk _00854_ net1227 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_140_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13039_ net270 net1917 net476 vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__mux2_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1160 net1162 vssd1 vssd1 vccd1 vccd1 net1160 sky130_fd_sc_hd__clkbuf_4
Xfanout1171 net1178 vssd1 vssd1 vccd1 vccd1 net1171 sky130_fd_sc_hd__clkbuf_4
XFILLER_94_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1182 net1185 vssd1 vssd1 vccd1 vccd1 net1182 sky130_fd_sc_hd__clkbuf_4
XFILLER_82_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12797__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1193 net1194 vssd1 vssd1 vccd1 vccd1 net1193 sky130_fd_sc_hd__clkbuf_2
X_07600_ datapath.rf.registers\[23\]\[19\] net700 net689 datapath.rf.registers\[31\]\[19\]
+ _02425_ vssd1 vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__a221o_1
XFILLER_94_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08580_ _03405_ _03407_ _03411_ _03415_ vssd1 vssd1 vccd1 vccd1 _03416_ sky130_fd_sc_hd__or4_1
X_07531_ datapath.rf.registers\[22\]\[20\] net734 net668 datapath.rf.registers\[21\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__a22o_1
XANTENNA__11273__Y _05723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08321__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07462_ datapath.rf.registers\[18\]\[21\] net790 _02288_ _02289_ _02294_ vssd1 vssd1
+ vccd1 vccd1 _02298_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07675__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08872__A1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09201_ net563 net553 net549 vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__or3_1
X_07393_ datapath.rf.registers\[25\]\[23\] net726 net722 datapath.rf.registers\[18\]\[23\]
+ _02226_ vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__a221o_1
XANTENNA__10447__C_N _05211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08582__Y _03418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11759__B2 _02439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09132_ net325 _03967_ vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__and2_1
XANTENNA_wire590_X net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10431__A1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09063_ _03896_ _03898_ net341 vssd1 vssd1 vccd1 vccd1 _03899_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout213_A _05634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08014_ _02840_ _02847_ _02848_ _02849_ vssd1 vssd1 vccd1 vccd1 _02850_ sky130_fd_sc_hd__or4_1
Xhold610 datapath.rf.registers\[31\]\[7\] vssd1 vssd1 vccd1 vccd1 net1958 sky130_fd_sc_hd__dlygate4sd3_1
Xhold621 datapath.rf.registers\[28\]\[13\] vssd1 vssd1 vccd1 vccd1 net1969 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold632 datapath.rf.registers\[12\]\[11\] vssd1 vssd1 vccd1 vccd1 net1980 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08388__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold643 datapath.rf.registers\[26\]\[11\] vssd1 vssd1 vccd1 vccd1 net1991 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold654 datapath.rf.registers\[27\]\[15\] vssd1 vssd1 vccd1 vccd1 net2002 sky130_fd_sc_hd__dlygate4sd3_1
Xhold665 datapath.rf.registers\[26\]\[18\] vssd1 vssd1 vccd1 vccd1 net2013 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold676 datapath.rf.registers\[18\]\[6\] vssd1 vssd1 vccd1 vccd1 net2024 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold687 datapath.rf.registers\[17\]\[24\] vssd1 vssd1 vccd1 vccd1 net2035 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07060__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold698 datapath.rf.registers\[8\]\[23\] vssd1 vssd1 vccd1 vccd1 net2046 sky130_fd_sc_hd__dlygate4sd3_1
X_09965_ _04762_ _04763_ _04798_ _04759_ _04756_ vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__a311o_1
XFILLER_58_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09337__C1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08916_ datapath.PC\[30\] _03751_ vssd1 vssd1 vccd1 vccd1 _03752_ sky130_fd_sc_hd__nor2_1
X_09896_ datapath.PC\[18\] _04731_ vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__and2_1
XFILLER_58_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08847_ _03228_ _01646_ _03671_ vssd1 vssd1 vccd1 vccd1 _03683_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout847_A _01737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12500__S net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08778_ _03601_ _03612_ vssd1 vssd1 vccd1 vccd1 _03614_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_0_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07729_ datapath.rf.registers\[17\]\[16\] net849 net807 datapath.rf.registers\[27\]\[16\]
+ _02564_ vssd1 vssd1 vccd1 vccd1 _02565_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout635_X net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11116__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10740_ net1517 net569 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[26\]
+ sky130_fd_sc_hd__and2_1
XFILLER_81_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10671_ button\[2\] net1022 vssd1 vssd1 vccd1 vccd1 _05489_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout802_X net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12410_ net1384 net130 _06352_ vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__a21o_1
XFILLER_138_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13390_ clknet_leaf_0_clk _00200_ net1056 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07418__A2 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12341_ net225 _05642_ _06309_ net895 vssd1 vssd1 vccd1 vccd1 _06310_ sky130_fd_sc_hd__o211a_1
XFILLER_139_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09110__A _03935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08091__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12272_ _05532_ _06254_ vssd1 vssd1 vccd1 vccd1 _06260_ sky130_fd_sc_hd__nor2_1
XANTENNA__07268__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14011_ clknet_leaf_75_clk _00002_ net1247 vssd1 vssd1 vccd1 vccd1 mmio.wishbone.curr_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08379__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11223_ net248 net2608 net527 vssd1 vssd1 vccd1 vccd1 _00273_ sky130_fd_sc_hd__mux2_1
XFILLER_153_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11154_ net254 net2022 net531 vssd1 vssd1 vccd1 vccd1 _00207_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10105_ _04891_ _04889_ vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__nand2b_1
X_11085_ net263 net2307 net537 vssd1 vssd1 vccd1 vccd1 _00142_ sky130_fd_sc_hd__mux2_1
XFILLER_0_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10036_ _04871_ vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__inv_2
XFILLER_76_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13803__Q mmio.memload_or_instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11987_ screen.register.currentYbus\[24\] _05757_ _06019_ screen.register.currentYbus\[8\]
+ _06031_ vssd1 vssd1 vccd1 vccd1 _06032_ sky130_fd_sc_hd__a221o_1
XANTENNA__08303__B1 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11026__S net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13726_ clknet_leaf_147_clk _00536_ net1064 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_27_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08854__A1 _02467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10938_ datapath.PC\[30\] _05671_ vssd1 vssd1 vccd1 vccd1 _05678_ sky130_fd_sc_hd__nand2_1
XFILLER_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10869_ _05617_ _05618_ vssd1 vssd1 vccd1 vccd1 _05619_ sky130_fd_sc_hd__or2_1
X_13657_ clknet_leaf_30_clk _00467_ net1124 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09939__B _03150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12608_ _06451_ _06452_ _06453_ _06446_ vssd1 vssd1 vccd1 vccd1 _06454_ sky130_fd_sc_hd__a211o_1
XANTENNA__08335__S net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13588_ clknet_leaf_129_clk _00398_ net1209 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09803__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08562__C _01816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10166__A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12539_ datapath.mulitply_result\[5\] datapath.multiplication_module.multiplicand_i\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06396_ sky130_fd_sc_hd__nor2_1
XANTENNA__08082__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13202__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07290__B1 _02124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09567__C1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14209_ clknet_leaf_47_clk datapath.multiplication_module.multiplicand_i_n\[20\]
+ net1172 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10453__X _05288_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10716__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07042__B1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout408 _05733_ vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__clkbuf_8
Xfanout419 _05722_ vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__buf_4
XFILLER_141_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09750_ _04146_ _04585_ vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__nand2_1
X_06962_ net914 _01797_ vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__and2_1
X_08701_ _02912_ _02936_ vssd1 vssd1 vccd1 vccd1 _03537_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_107_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11677__B1 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09681_ _04496_ _04516_ vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__nand2_1
X_06893_ datapath.rf.registers\[4\]\[31\] net864 net860 datapath.rf.registers\[16\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__a22o_1
XANTENNA__08542__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08632_ _03466_ _03462_ vssd1 vssd1 vccd1 vccd1 _03468_ sky130_fd_sc_hd__nand2b_1
XFILLER_55_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07896__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08563_ datapath.rf.registers\[21\]\[0\] net966 _01831_ vssd1 vssd1 vccd1 vccd1 _03399_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12451__A1_N net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09098__A1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout163_A _05933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07514_ datapath.rf.registers\[13\]\[20\] net810 net807 datapath.rf.registers\[27\]\[20\]
+ _02338_ vssd1 vssd1 vccd1 vccd1 _02350_ sky130_fd_sc_hd__a221o_1
XANTENNA__10101__B1 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07648__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08494_ datapath.rf.registers\[23\]\[1\] net965 _01820_ vssd1 vssd1 vccd1 vccd1 _03330_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08845__A1 _02170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07445_ datapath.rf.registers\[2\]\[22\] net742 net683 datapath.rf.registers\[27\]\[22\]
+ _02279_ vssd1 vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout428_A net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13151__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07376_ datapath.rf.registers\[24\]\[23\] net856 net807 datapath.rf.registers\[27\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__a22o_1
X_09115_ _03498_ _03499_ vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__nand2b_2
XFILLER_109_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12990__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1278_A mmio.memload_or_instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08073__A2 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09046_ net462 _03840_ _03841_ vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__and3_1
XFILLER_124_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07820__A2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout797_A net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold440 datapath.rf.registers\[6\]\[23\] vssd1 vssd1 vccd1 vccd1 net1788 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10363__X _05199_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12291__A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold451 datapath.rf.registers\[5\]\[31\] vssd1 vssd1 vccd1 vccd1 net1799 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold462 datapath.rf.registers\[20\]\[13\] vssd1 vssd1 vccd1 vccd1 net1810 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold473 datapath.rf.registers\[12\]\[31\] vssd1 vssd1 vccd1 vccd1 net1821 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold484 datapath.rf.registers\[2\]\[13\] vssd1 vssd1 vccd1 vccd1 net1832 sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 datapath.rf.registers\[18\]\[29\] vssd1 vssd1 vccd1 vccd1 net1843 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout964_A net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06720__C _01502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout920 _01744_ vssd1 vssd1 vccd1 vccd1 net920 sky130_fd_sc_hd__buf_2
Xfanout931 net933 vssd1 vssd1 vccd1 vccd1 net931 sky130_fd_sc_hd__buf_2
XFILLER_132_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_5_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout942 _01717_ vssd1 vssd1 vccd1 vccd1 net942 sky130_fd_sc_hd__buf_2
X_09948_ datapath.PC\[0\] _03384_ _04782_ _04780_ vssd1 vssd1 vccd1 vccd1 _04784_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__08768__X _03604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout953 net954 vssd1 vssd1 vccd1 vccd1 net953 sky130_fd_sc_hd__clkbuf_2
Xfanout964 net965 vssd1 vssd1 vccd1 vccd1 net964 sky130_fd_sc_hd__buf_1
Xfanout975 net980 vssd1 vssd1 vccd1 vccd1 net975 sky130_fd_sc_hd__buf_2
Xfanout986 net987 vssd1 vssd1 vccd1 vccd1 net986 sky130_fd_sc_hd__clkbuf_2
Xfanout997 _05789_ vssd1 vssd1 vccd1 vccd1 net997 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_51_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout752_X net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09879_ _03728_ _04714_ vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_51_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1140 datapath.rf.registers\[31\]\[13\] vssd1 vssd1 vccd1 vccd1 net2488 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1151 datapath.rf.registers\[28\]\[21\] vssd1 vssd1 vccd1 vccd1 net2499 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1162 datapath.rf.registers\[29\]\[14\] vssd1 vssd1 vccd1 vccd1 net2510 sky130_fd_sc_hd__dlygate4sd3_1
X_11910_ net136 _05970_ _05969_ vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__o21ai_1
XFILLER_58_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1173 datapath.rf.registers\[2\]\[25\] vssd1 vssd1 vccd1 vccd1 net2521 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10340__B1 net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12890_ net186 net2076 net399 vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__mux2_1
Xhold1184 datapath.rf.registers\[17\]\[21\] vssd1 vssd1 vccd1 vccd1 net2532 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06729__A net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1195 screen.register.currentYbus\[24\] vssd1 vssd1 vccd1 vccd1 net2543 sky130_fd_sc_hd__dlygate4sd3_1
X_11841_ net1280 _01425_ _05296_ _05817_ vssd1 vssd1 vccd1 vccd1 _05920_ sky130_fd_sc_hd__or4b_1
XFILLER_14_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11772_ net1291 net151 net152 vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__a21o_1
X_14560_ clknet_leaf_136_clk _01265_ net1090 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07639__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08836__A1 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11675__A1_N _05085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13511_ clknet_leaf_137_clk _00321_ net1089 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10723_ net1600 _02912_ net572 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[9\]
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_24_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14491_ clknet_leaf_36_clk _01196_ net1136 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08663__B _02240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10654_ _05472_ vssd1 vssd1 vccd1 vccd1 _05473_ sky130_fd_sc_hd__inv_2
X_13442_ clknet_leaf_151_clk _00252_ net1052 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_41_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14168__RESET_B net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13373_ clknet_leaf_147_clk _00183_ net1064 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10585_ _03028_ _03076_ _03123_ _03170_ vssd1 vssd1 vccd1 vccd1 _05408_ sky130_fd_sc_hd__or4_1
XANTENNA__08064__A2 _01749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload18 clknet_leaf_146_clk vssd1 vssd1 vccd1 vccd1 clkload18/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload29 clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 clkload29/X sky130_fd_sc_hd__clkbuf_8
XFILLER_154_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12324_ _04118_ _06297_ net894 vssd1 vssd1 vccd1 vccd1 _06298_ sky130_fd_sc_hd__mux2_1
XANTENNA__07811__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12255_ datapath.multiplication_module.zero_multi _06245_ _01407_ datapath.pc_module.i_ack2
+ vssd1 vssd1 vccd1 vccd1 _06246_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_108_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09013__A1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11206_ _05513_ _05712_ vssd1 vssd1 vccd1 vccd1 _05720_ sky130_fd_sc_hd__nor2_1
XFILLER_141_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12186_ _06201_ _06202_ vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_71_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11137_ net174 net2038 net428 vssd1 vssd1 vccd1 vccd1 _00192_ sky130_fd_sc_hd__mux2_1
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07582__X _02418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11068_ net174 net1608 net432 vssd1 vssd1 vccd1 vccd1 _00128_ sky130_fd_sc_hd__mux2_1
X_10019_ _04835_ _04851_ _04854_ vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__nor3_1
XFILLER_37_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14758_ screen.dcx vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__clkbuf_1
X_13709_ clknet_leaf_132_clk _00519_ net1112 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_149_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14689_ clknet_leaf_45_clk _01394_ net1148 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_07230_ datapath.rf.registers\[30\]\[26\] net832 net799 datapath.rf.registers\[15\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__a22o_1
XFILLER_146_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07161_ datapath.rf.registers\[14\]\[28\] net776 net757 datapath.rf.registers\[12\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01997_ sky130_fd_sc_hd__a22o_1
XFILLER_9_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06661__X _01500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07092_ datapath.rf.registers\[2\]\[29\] net888 net853 datapath.rf.registers\[19\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__a22o_1
XFILLER_145_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07476__Y _02312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07015__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout205 _05641_ vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10343__B net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout216 net217 vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08763__B1 _01859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout227 _04712_ vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__clkbuf_4
X_09802_ _04047_ _04637_ net339 vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__mux2_1
Xfanout238 _05616_ vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__buf_1
Xfanout249 net250 vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__dlymetal6s2s_1
X_07994_ datapath.rf.registers\[25\]\[10\] net843 net791 datapath.rf.registers\[18\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__a22o_1
XFILLER_101_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09733_ net360 _04415_ net346 vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__a21oi_1
X_06945_ MemWrite _01780_ vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout280_A _05554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12311__A1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13146__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09664_ net358 _04498_ net325 vssd1 vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__o21a_1
X_06876_ _01630_ _01638_ vssd1 vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__nor2_4
XFILLER_131_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08467__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08615_ _02545_ _03448_ _02544_ vssd1 vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__a21oi_1
XANTENNA__14188__D net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12985__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09595_ _04305_ _04306_ net457 vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__a21oi_1
XFILLER_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08546_ _03371_ _03373_ _03377_ _03381_ vssd1 vssd1 vccd1 vccd1 _03382_ sky130_fd_sc_hd__or4b_2
XFILLER_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11902__B net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_862 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08477_ datapath.rf.registers\[20\]\[1\] net840 net820 datapath.rf.registers\[5\]\[1\]
+ _03312_ vssd1 vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__a221o_1
XANTENNA__11822__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout333_X net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08294__A2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout712_A net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1075_X net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07428_ datapath.rf.registers\[0\]\[22\] net866 _02255_ _02263_ vssd1 vssd1 vccd1
+ vccd1 _02264_ sky130_fd_sc_hd__o22a_4
XFILLER_155_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07359_ datapath.rf.registers\[23\]\[23\] net940 net921 vssd1 vssd1 vccd1 vccd1 _02195_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout500_X net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10389__B1 _01607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_149_Right_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10370_ net1269 net466 vssd1 vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__nor2_1
XFILLER_152_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09029_ _03830_ _03864_ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__nand2_1
XFILLER_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07006__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12040_ screen.register.currentYbus\[3\] _05778_ net999 screen.register.currentXbus\[11\]
+ vssd1 vssd1 vccd1 vccd1 _06082_ sky130_fd_sc_hd__a22o_1
Xhold270 datapath.rf.registers\[7\]\[16\] vssd1 vssd1 vccd1 vccd1 net1618 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_53_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold281 datapath.rf.registers\[4\]\[19\] vssd1 vssd1 vccd1 vccd1 net1629 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout967_X net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold292 datapath.rf.registers\[9\]\[3\] vssd1 vssd1 vccd1 vccd1 net1640 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout750 _01804_ vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_148_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout761 _01802_ vssd1 vssd1 vccd1 vccd1 net761 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_148_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout772 net773 vssd1 vssd1 vccd1 vccd1 net772 sky130_fd_sc_hd__buf_4
X_13991_ clknet_leaf_108_clk _00768_ net1218 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout783 net784 vssd1 vssd1 vccd1 vccd1 net783 sky130_fd_sc_hd__clkbuf_8
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07309__B2 _02144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout794 net795 vssd1 vssd1 vccd1 vccd1 net794 sky130_fd_sc_hd__clkbuf_8
XANTENNA__13056__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07562__B net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12942_ net257 net1925 net395 vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__mux2_1
XFILLER_86_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12873_ net272 net2268 net400 vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__mux2_1
X_14612_ clknet_leaf_129_clk _01317_ net1209 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11824_ net2230 net1050 net315 net335 datapath.ru.latched_instruction\[30\] vssd1
+ vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__a32o_1
XANTENNA__06746__X _01585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08674__A _02466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11813__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14543_ clknet_leaf_28_clk _01248_ net1155 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11755_ net1474 net145 net140 _02634_ vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__a22o_1
XANTENNA__08285__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09482__A1 _02857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11304__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07493__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10706_ net1451 _02824_ net571 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i_n\[11\]
+ sky130_fd_sc_hd__mux2_1
X_14474_ clknet_leaf_60_clk _01179_ net1169 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11686_ _05167_ net152 net151 net1426 vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__a22o_1
Xmax_cap1012 _06152_ vssd1 vssd1 vccd1 vccd1 net1012 sky130_fd_sc_hd__clkbuf_2
X_13425_ clknet_leaf_40_clk _00235_ net1140 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10637_ _05435_ _05437_ _05430_ vssd1 vssd1 vccd1 vccd1 _05457_ sky130_fd_sc_hd__o21a_1
XANTENNA__08037__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload107 clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 clkload107/Y sky130_fd_sc_hd__inv_8
Xclkload118 clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 clkload118/Y sky130_fd_sc_hd__inv_6
Xclkload129 clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 clkload129/Y sky130_fd_sc_hd__clkinv_8
X_10568_ screen.register.currentXbus\[13\] screen.register.currentXbus\[12\] screen.register.currentXbus\[15\]
+ screen.register.currentXbus\[14\] vssd1 vssd1 vccd1 vccd1 _05392_ sky130_fd_sc_hd__or4_1
X_13356_ clknet_leaf_15_clk _00166_ net1105 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_116_Right_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06922__A net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_926 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12307_ _06284_ _06285_ net890 _04239_ vssd1 vssd1 vccd1 vccd1 _06286_ sky130_fd_sc_hd__o2bb2a_1
X_13287_ clknet_leaf_145_clk _00097_ net1089 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10499_ _05323_ _05324_ _05328_ vssd1 vssd1 vccd1 vccd1 _05329_ sky130_fd_sc_hd__or3b_1
X_12238_ screen.counter.currentCt\[17\] _06233_ net602 vssd1 vssd1 vccd1 vccd1 _06235_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__07456__C net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12169_ _06157_ _06172_ vssd1 vssd1 vccd1 vccd1 _06192_ sky130_fd_sc_hd__and2_1
XFILLER_111_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07753__A net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput5 DAT_I[12] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
X_06730_ _01450_ net1014 vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__and2_1
X_06661_ mmio.key_data\[0\] mmio.memload_or_instruction\[0\] net1048 vssd1 vssd1 vccd1
+ vccd1 _01500_ sky130_fd_sc_hd__mux2_4
XFILLER_37_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_84_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08400_ datapath.rf.registers\[20\]\[2\] net960 net926 vssd1 vssd1 vccd1 vccd1 _03236_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12057__B1 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09380_ net460 _04214_ _04215_ vssd1 vssd1 vccd1 vccd1 _04216_ sky130_fd_sc_hd__and3_1
X_06592_ columns.count\[1\] columns.count\[3\] columns.count\[2\] vssd1 vssd1 vccd1
+ vccd1 _01433_ sky130_fd_sc_hd__and3_1
XANTENNA__08584__A net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08331_ datapath.rf.registers\[26\]\[4\] net778 net694 datapath.rf.registers\[8\]\[4\]
+ _03166_ vssd1 vssd1 vccd1 vccd1 _03167_ sky130_fd_sc_hd__a221o_1
XANTENNA__14019__RESET_B net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08276__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11214__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07484__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08262_ datapath.rf.registers\[12\]\[5\] net827 net808 datapath.rf.registers\[27\]\[5\]
+ _03084_ vssd1 vssd1 vccd1 vccd1 _03098_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_15_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07213_ _02026_ _02047_ vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__nand2_1
XANTENNA__08028__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08193_ _01598_ _01784_ vssd1 vssd1 vccd1 vccd1 _03029_ sky130_fd_sc_hd__nor2_1
XANTENNA__10906__X _05651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout126_A net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07236__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07144_ datapath.rf.registers\[0\]\[28\] _01724_ _01970_ _01979_ vssd1 vssd1 vccd1
+ vccd1 _01980_ sky130_fd_sc_hd__o22a_4
XTAP_TAPCELL_ROW_115_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07075_ _01889_ _01909_ vssd1 vssd1 vccd1 vccd1 _01911_ sky130_fd_sc_hd__or2_1
XFILLER_145_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07366__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout495_A _06550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout662_A net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07977_ datapath.rf.registers\[20\]\[11\] net720 net700 datapath.rf.registers\[23\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__a22o_1
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09716_ _03534_ net629 _04551_ net646 vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__a211o_1
XFILLER_28_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06928_ _01630_ _01639_ _01657_ net961 vssd1 vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__and4_2
XFILLER_28_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09647_ net373 _04318_ _04320_ net327 vssd1 vssd1 vccd1 vccd1 _04483_ sky130_fd_sc_hd__a31oi_1
X_06859_ datapath.ru.latched_instruction\[4\] _01571_ _01638_ datapath.ru.latched_instruction\[18\]
+ vssd1 vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout927_A _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09578_ net460 _04351_ _04412_ vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__a21o_1
XFILLER_82_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08529_ datapath.rf.registers\[11\]\[0\] net884 net809 datapath.rf.registers\[27\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03365_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout715_X net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11124__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11540_ _05753_ _05763_ vssd1 vssd1 vccd1 vccd1 _05764_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_46_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11810__A3 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11471_ net2420 net186 net407 vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__mux2_1
XANTENNA__10963__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14035__SET_B net1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13210_ clknet_leaf_2_clk _00020_ net1063 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10422_ net366 _05257_ net371 vssd1 vssd1 vccd1 vccd1 _05258_ sky130_fd_sc_hd__a21oi_1
XFILLER_137_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14190_ clknet_leaf_91_clk datapath.multiplication_module.multiplicand_i_n\[1\] net1241
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_152_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10535__Y screen.counter.ack vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13141_ net1631 net254 net383 vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__mux2_1
X_10353_ _04496_ _04516_ vssd1 vssd1 vccd1 vccd1 _05189_ sky130_fd_sc_hd__nor2_1
XANTENNA__07557__B net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13072_ net1791 net271 net388 vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__mux2_1
X_10284_ _03735_ _05119_ net1038 vssd1 vssd1 vccd1 vccd1 _05120_ sky130_fd_sc_hd__a21oi_1
XFILLER_152_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12023_ screen.register.currentXbus\[2\] _05755_ _05768_ screen.register.currentXbus\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06066_ sky130_fd_sc_hd__a22o_1
XANTENNA__08669__A _02364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10711__B _05368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout580 _03605_ vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__buf_2
XFILLER_120_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13974_ clknet_leaf_105_clk _00752_ net1224 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12925_ net2580 net181 net483 vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12856_ net195 net2011 net486 vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__mux2_1
XFILLER_73_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06917__A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08835__C _03669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11807_ _01446_ net1017 net315 net335 datapath.ru.latched_instruction\[13\] vssd1
+ vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__a32o_1
XANTENNA__08258__A2 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12787_ net204 net1645 net494 vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__mux2_1
XANTENNA__11034__S net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07466__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14526_ clknet_leaf_150_clk _01231_ net1059 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08554__D _01800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11738_ net26 net1034 net1024 net2249 vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_12_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14457_ clknet_leaf_9_clk _01162_ net1074 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_11669_ _01405_ _05291_ _05883_ vssd1 vssd1 vccd1 vccd1 _05885_ sky130_fd_sc_hd__a21o_2
XFILLER_128_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13408_ clknet_leaf_138_clk _00218_ net1098 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_14388_ clknet_leaf_93_clk _01093_ net1210 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08966__A0 _03800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10222__C1 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13339_ clknet_leaf_39_clk _00149_ net1145 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07900_ datapath.rf.registers\[2\]\[12\] net889 net830 datapath.rf.registers\[14\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02736_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_110_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08880_ _01614_ _01618_ vssd1 vssd1 vccd1 vccd1 _03716_ sky130_fd_sc_hd__or2_1
XFILLER_97_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07831_ datapath.rf.registers\[23\]\[14\] net699 net672 datapath.rf.registers\[7\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__a22o_1
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06744__A2 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11209__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07762_ datapath.rf.registers\[10\]\[15\] net880 net873 _02597_ vssd1 vssd1 vccd1
+ vccd1 _02598_ sky130_fd_sc_hd__a211o_1
X_09501_ net607 _04301_ _04336_ _03604_ net555 vssd1 vssd1 vccd1 vccd1 _04337_ sky130_fd_sc_hd__o221ai_1
X_06713_ mmio.memload_or_instruction\[14\] mmio.memload_or_instruction\[13\] mmio.memload_or_instruction\[12\]
+ mmio.memload_or_instruction\[11\] vssd1 vssd1 vccd1 vccd1 _01552_ sky130_fd_sc_hd__and4b_1
XPHY_EDGE_ROW_142_Left_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07693_ datapath.rf.registers\[26\]\[17\] net780 net689 datapath.rf.registers\[31\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02529_ sky130_fd_sc_hd__a22o_1
XFILLER_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09694__B2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06644_ datapath.ru.latched_instruction\[27\] _01479_ _01482_ _01476_ _01478_ vssd1
+ vssd1 vccd1 vccd1 _01483_ sky130_fd_sc_hd__o2111a_1
XFILLER_80_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09432_ net323 _04267_ vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__nor2_1
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09363_ _03957_ _04198_ net376 vssd1 vssd1 vccd1 vccd1 _04199_ sky130_fd_sc_hd__mux2_1
X_06575_ net1269 vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__inv_2
XANTENNA__08249__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07457__B1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08314_ _01641_ _01703_ _01783_ net967 vssd1 vssd1 vccd1 vccd1 _03150_ sky130_fd_sc_hd__a22o_1
XANTENNA__12450__B1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09294_ _02466_ net553 net549 vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__or3_1
XANTENNA_10 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08245_ net560 _03078_ vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__nand2_1
XFILLER_21_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout410_A _05730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1152_A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout508_A net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08176_ datapath.rf.registers\[26\]\[7\] net780 net760 datapath.rf.registers\[30\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03012_ sky130_fd_sc_hd__a22o_1
X_07127_ datapath.rf.registers\[2\]\[28\] _01713_ _01721_ datapath.rf.registers\[10\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__a22o_1
XFILLER_119_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_63_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08421__A2 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07058_ datapath.rf.registers\[15\]\[30\] net666 net662 datapath.rf.registers\[5\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__a22o_1
Xteam_04_1299 vssd1 vssd1 vccd1 vccd1 team_04_1299/HI gpio_oeb[4] sky130_fd_sc_hd__conb_1
XANTENNA_fanout877_A net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12503__S net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09084__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_78_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_145_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_145_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout665_X net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11119__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_121_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12269__B1 _06253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08001__B net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout832_X net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10971_ net1545 net288 net436 vssd1 vssd1 vccd1 vccd1 _00036_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12710_ _05892_ _06530_ _01404_ vssd1 vssd1 vccd1 vccd1 _06536_ sky130_fd_sc_hd__o21ai_1
XFILLER_44_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07696__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13690_ clknet_leaf_135_clk _00500_ net1102 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06737__A _01571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07160__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_136_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12641_ datapath.mulitply_result\[22\] datapath.multiplication_module.multiplicand_i\[22\]
+ vssd1 vssd1 vccd1 vccd1 _06481_ sky130_fd_sc_hd__nand2_1
XFILLER_62_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_16_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07448__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12572_ _06422_ _06423_ vssd1 vssd1 vccd1 vccd1 _06424_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_61_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14311_ clknet_leaf_140_clk _01016_ net1097 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[31\]
+ sky130_fd_sc_hd__dfrtp_2
X_11523_ datapath.i_ack _05747_ WEN vssd1 vssd1 vccd1 vccd1 _00547_ sky130_fd_sc_hd__a21o_1
XFILLER_11_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09767__B _04118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14242_ clknet_leaf_124_clk datapath.multiplication_module.multiplier_i_n\[10\] net1215
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_156_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11454_ net2163 net273 net408 vssd1 vssd1 vccd1 vccd1 _00492_ sky130_fd_sc_hd__mux2_1
XFILLER_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06903__C net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10405_ datapath.PC\[0\] _03384_ _04783_ vssd1 vssd1 vccd1 vccd1 _05241_ sky130_fd_sc_hd__a21o_1
X_14173_ clknet_leaf_47_clk _00928_ net1174 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_11385_ net2066 net278 net412 vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__mux2_1
XANTENNA__08412__A2 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13124_ net181 net2451 net473 vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__mux2_1
X_10336_ _04272_ _04582_ _04239_ vssd1 vssd1 vccd1 vccd1 _05172_ sky130_fd_sc_hd__o21a_1
XANTENNA__07620__B1 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_9_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_9_0_clk sky130_fd_sc_hd__clkbuf_8
X_10267_ net1266 _03738_ datapath.PC\[13\] vssd1 vssd1 vccd1 vccd1 _05103_ sky130_fd_sc_hd__o21ai_1
X_13055_ net194 net2289 net475 vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__mux2_1
XFILLER_87_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12006_ _06047_ _06049_ net1011 vssd1 vssd1 vccd1 vccd1 _06050_ sky130_fd_sc_hd__o21a_1
X_10198_ datapath.PC\[23\] _03978_ net469 vssd1 vssd1 vccd1 vccd1 _05034_ sky130_fd_sc_hd__mux2_1
XFILLER_94_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11029__S net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13957_ clknet_leaf_107_clk _00735_ net1220 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09676__A1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08479__A2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12908_ net2493 net264 net485 vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__mux2_1
XANTENNA__07687__B1 _02521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13888_ clknet_leaf_49_clk _00692_ net1176 vssd1 vssd1 vccd1 vccd1 keypad.alpha sky130_fd_sc_hd__dfrtp_4
XFILLER_50_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07151__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12839_ net274 net2064 net488 vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__mux2_1
XANTENNA__10169__A net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07439__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14509_ clknet_leaf_125_clk _01214_ net1205 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_08030_ datapath.rf.registers\[10\]\[10\] net708 net704 datapath.rf.registers\[9\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02866_ sky130_fd_sc_hd__a22o_1
Xinput30 DAT_I[6] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_96_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold803 datapath.rf.registers\[18\]\[19\] vssd1 vssd1 vccd1 vccd1 net2151 sky130_fd_sc_hd__dlygate4sd3_1
Xhold814 datapath.rf.registers\[0\]\[19\] vssd1 vssd1 vccd1 vccd1 net2162 sky130_fd_sc_hd__dlygate4sd3_1
Xhold825 datapath.rf.registers\[5\]\[26\] vssd1 vssd1 vccd1 vccd1 net2173 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold836 datapath.rf.registers\[11\]\[6\] vssd1 vssd1 vccd1 vccd1 net2184 sky130_fd_sc_hd__dlygate4sd3_1
Xhold847 datapath.mulitply_result\[12\] vssd1 vssd1 vccd1 vccd1 net2195 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10210__A2 _04600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07611__B1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold858 datapath.rf.registers\[12\]\[12\] vssd1 vssd1 vccd1 vccd1 net2206 sky130_fd_sc_hd__dlygate4sd3_1
X_09981_ datapath.PC\[22\] net595 vssd1 vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__nor2_1
Xhold869 datapath.rf.registers\[9\]\[16\] vssd1 vssd1 vccd1 vccd1 net2217 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08932_ net329 _03767_ _03623_ vssd1 vssd1 vccd1 vccd1 _03768_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12323__S net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08863_ _03669_ _03672_ vssd1 vssd1 vccd1 vccd1 _03699_ sky130_fd_sc_hd__nand2b_1
XFILLER_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout193_A _05659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11710__A2 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_150_Left_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07814_ datapath.rf.registers\[3\]\[14\] net802 net796 datapath.rf.registers\[29\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02650_ sky130_fd_sc_hd__a22o_1
X_08794_ _03617_ net367 vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__or2_1
XANTENNA__07390__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10778__S net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07745_ datapath.rf.registers\[3\]\[16\] net770 net762 datapath.rf.registers\[1\]\[16\]
+ _02578_ vssd1 vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__a221o_1
XANTENNA__13154__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_140_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07678__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07676_ datapath.rf.registers\[17\]\[17\] net851 _02494_ _02496_ _02505_ vssd1 vssd1
+ vccd1 vccd1 _02512_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07142__A2 _01716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09415_ net356 net350 _03883_ vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__or3_2
X_06627_ net1288 net1283 mmio.memload_or_instruction\[30\] vssd1 vssd1 vccd1 vccd1
+ _01466_ sky130_fd_sc_hd__or3b_4
XFILLER_13_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12993__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout625_A _03721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08890__A2 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09346_ _03575_ _04179_ net580 vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__o21a_1
XANTENNA__08772__A net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09277_ net319 _03858_ vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout413_X net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08491__B net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11402__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08228_ datapath.rf.registers\[8\]\[6\] net694 net683 datapath.rf.registers\[27\]\[6\]
+ _03063_ vssd1 vssd1 vccd1 vccd1 _03064_ sky130_fd_sc_hd__a221o_1
XFILLER_148_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09874__Y _04710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08159_ datapath.rf.registers\[28\]\[7\] net806 net794 datapath.rf.registers\[31\]\[7\]
+ _02994_ vssd1 vssd1 vccd1 vccd1 _02995_ sky130_fd_sc_hd__a221o_1
XFILLER_134_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11170_ net183 net2201 net531 vssd1 vssd1 vccd1 vccd1 _00223_ sky130_fd_sc_hd__mux2_1
XANTENNA__07602__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout782_X net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10121_ net895 _04057_ _04603_ vssd1 vssd1 vccd1 vccd1 _04957_ sky130_fd_sc_hd__nor3_1
XFILLER_122_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10052_ _04826_ _04887_ vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__xor2_1
XFILLER_76_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07554__C net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13811_ clknet_leaf_141_clk _00620_ net1095 vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__dfrtp_1
XANTENNA_input19_A DAT_I[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13064__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13742_ clknet_leaf_50_clk _00552_ net1181 vssd1 vssd1 vccd1 vccd1 mmio.key_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10954_ _01644_ _01663_ vssd1 vssd1 vccd1 vccd1 _05692_ sky130_fd_sc_hd__or2_1
XANTENNA__07133__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13673_ clknet_leaf_91_clk _00483_ net1232 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13757__RESET_B net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10885_ datapath.mulitply_result\[22\] net597 net617 vssd1 vssd1 vccd1 vccd1 _05633_
+ sky130_fd_sc_hd__a21o_1
XFILLER_31_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12624_ datapath.mulitply_result\[19\] datapath.multiplication_module.multiplicand_i\[19\]
+ vssd1 vssd1 vccd1 vccd1 _06467_ sky130_fd_sc_hd__nor2_1
X_12555_ net2539 net505 net501 _06409_ vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__a22o_1
XANTENNA__11312__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11506_ net177 net2354 net512 vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__mux2_1
XFILLER_156_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07841__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12486_ net278 net2226 net508 vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__mux2_1
X_14225_ clknet_leaf_42_clk _00946_ net1144 vssd1 vssd1 vccd1 vccd1 columns.count\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11437_ net187 net2407 net515 vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__mux2_1
XFILLER_99_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14156_ clknet_leaf_67_clk _00911_ net1239 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06930__A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11368_ net197 net1885 net520 vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__mux2_1
XFILLER_153_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13107_ net262 net2627 net472 vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10319_ _04844_ _05154_ vssd1 vssd1 vccd1 vccd1 _05155_ sky130_fd_sc_hd__or2_1
X_14087_ clknet_leaf_108_clk _00853_ net1218 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_140_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11299_ _05653_ net1672 net524 vssd1 vssd1 vccd1 vccd1 _00347_ sky130_fd_sc_hd__mux2_1
XANTENNA__13142__A1 _05588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09346__B1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13038_ net274 net2004 net476 vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__mux2_1
XFILLER_67_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1150 net1151 vssd1 vssd1 vccd1 vccd1 net1150 sky130_fd_sc_hd__buf_2
XFILLER_67_857 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1161 net1162 vssd1 vssd1 vccd1 vccd1 net1161 sky130_fd_sc_hd__clkbuf_2
Xfanout1172 net1178 vssd1 vssd1 vccd1 vccd1 net1172 sky130_fd_sc_hd__buf_2
XFILLER_14_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1183 net1185 vssd1 vssd1 vccd1 vccd1 net1183 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10900__B1 _05644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06929__X _01765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1194 net1204 vssd1 vssd1 vccd1 vccd1 net1194 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07372__A2 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11554__Y _05778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08576__B net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10259__A2 net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07530_ datapath.rf.registers\[30\]\[20\] net760 net710 datapath.rf.registers\[11\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_105_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07461_ datapath.rf.registers\[10\]\[21\] net879 net832 datapath.rf.registers\[30\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__a22o_1
X_09200_ _03881_ _03882_ net356 net353 vssd1 vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__o211ai_1
XFILLER_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07392_ datapath.rf.registers\[24\]\[23\] net766 net730 datapath.rf.registers\[19\]\[23\]
+ _02227_ vssd1 vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__a221o_1
XANTENNA__06664__X _01503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09131_ net361 _03965_ _03966_ _03960_ vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__a31o_1
XANTENNA__08085__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11222__S net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09062_ net449 _03704_ _03897_ vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__a21oi_1
XFILLER_148_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07832__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08013_ datapath.rf.registers\[23\]\[10\] net814 _02828_ _02836_ _02837_ vssd1 vssd1
+ vccd1 vccd1 _02849_ sky130_fd_sc_hd__a2111o_1
Xhold600 datapath.rf.registers\[23\]\[15\] vssd1 vssd1 vccd1 vccd1 net1948 sky130_fd_sc_hd__dlygate4sd3_1
Xhold611 datapath.rf.registers\[18\]\[5\] vssd1 vssd1 vccd1 vccd1 net1959 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout206_A _05641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold622 datapath.rf.registers\[21\]\[4\] vssd1 vssd1 vccd1 vccd1 net1970 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07495__X _02331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold633 datapath.rf.registers\[4\]\[1\] vssd1 vssd1 vccd1 vccd1 net1981 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold644 datapath.rf.registers\[22\]\[17\] vssd1 vssd1 vccd1 vccd1 net1992 sky130_fd_sc_hd__dlygate4sd3_1
Xhold655 datapath.rf.registers\[2\]\[20\] vssd1 vssd1 vccd1 vccd1 net2003 sky130_fd_sc_hd__dlygate4sd3_1
Xhold666 datapath.rf.registers\[22\]\[26\] vssd1 vssd1 vccd1 vccd1 net2014 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06938__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13149__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold677 datapath.rf.registers\[6\]\[22\] vssd1 vssd1 vccd1 vccd1 net2025 sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 datapath.rf.registers\[23\]\[24\] vssd1 vssd1 vccd1 vccd1 net2036 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold699 datapath.rf.registers\[10\]\[30\] vssd1 vssd1 vccd1 vccd1 net2047 sky130_fd_sc_hd__dlygate4sd3_1
X_09964_ _04760_ _04763_ _04798_ _04759_ vssd1 vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__a31oi_1
XFILLER_134_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1115_A net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08915_ datapath.PC\[29\] _03750_ vssd1 vssd1 vccd1 vccd1 _03751_ sky130_fd_sc_hd__or2_1
XFILLER_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09895_ _01639_ _03670_ net604 vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__a21o_1
XANTENNA__12988__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1300 screen.register.currentXbus\[7\] vssd1 vssd1 vccd1 vccd1 net2648 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout575_A _03666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08846_ _03680_ _03681_ net449 vssd1 vssd1 vccd1 vccd1 _03682_ sky130_fd_sc_hd__mux2_1
XFILLER_85_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout742_A net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08777_ _03601_ _03612_ vssd1 vssd1 vccd1 vccd1 _03613_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_0_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07728_ datapath.rf.registers\[1\]\[16\] net845 net804 datapath.rf.registers\[28\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02564_ sky130_fd_sc_hd__a22o_1
XANTENNA__10104__D1 _01586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07115__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout530_X net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07659_ datapath.rf.registers\[27\]\[17\] net973 net939 vssd1 vssd1 vccd1 vccd1 _02495_
+ sky130_fd_sc_hd__and3_1
XFILLER_81_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11921__A _02331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10670_ _01430_ _05481_ _05485_ _05488_ vssd1 vssd1 vccd1 vccd1 keypad.decode.button_n\[1\]
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_43_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09329_ net346 _04164_ vssd1 vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__or2_1
XANTENNA__08076__B1 _02911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11132__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12340_ net225 _04831_ vssd1 vssd1 vccd1 vccd1 _06309_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_153_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout997_X net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10971__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12271_ net892 _04842_ net190 vssd1 vssd1 vccd1 vccd1 _06259_ sky130_fd_sc_hd__a21oi_1
XFILLER_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14010_ clknet_leaf_75_clk _00001_ net1247 vssd1 vssd1 vccd1 vccd1 mmio.wishbone.curr_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11222_ net252 net2194 net527 vssd1 vssd1 vccd1 vccd1 _00272_ sky130_fd_sc_hd__mux2_1
XANTENNA__07846__A _02661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10186__A1 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06750__A _01579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13059__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11153_ net263 net2352 net532 vssd1 vssd1 vccd1 vccd1 _00206_ sky130_fd_sc_hd__mux2_1
XANTENNA__10272__A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10104_ _03865_ _04625_ _04939_ net901 _01586_ vssd1 vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__o2111ai_1
XFILLER_1_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11084_ net266 net1839 net536 vssd1 vssd1 vccd1 vccd1 _00141_ sky130_fd_sc_hd__mux2_1
XANTENNA__12898__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10035_ _04812_ _04870_ vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07354__A2 _02189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08396__B net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06909__B _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11986_ screen.register.currentXbus\[8\] _05768_ _05772_ screen.register.currentXbus\[24\]
+ vssd1 vssd1 vccd1 vccd1 _06031_ sky130_fd_sc_hd__a22o_1
XANTENNA__08964__X _03800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07106__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13725_ clknet_leaf_148_clk _00535_ net1060 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10937_ net182 net2576 net545 vssd1 vssd1 vccd1 vccd1 _00031_ sky130_fd_sc_hd__mux2_1
XFILLER_44_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13656_ clknet_leaf_3_clk _00466_ net1077 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10868_ datapath.PC\[20\] _05611_ vssd1 vssd1 vccd1 vccd1 _05618_ sky130_fd_sc_hd__nor2_1
XFILLER_31_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08067__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12607_ _06440_ _06444_ _06447_ vssd1 vssd1 vccd1 vccd1 _06453_ sky130_fd_sc_hd__a21oi_1
X_13587_ clknet_leaf_34_clk _00397_ net1127 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10447__A _05240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11042__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10799_ net1267 datapath.PC\[10\] _05548_ vssd1 vssd1 vccd1 vccd1 _05559_ sky130_fd_sc_hd__and3_1
XFILLER_8_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07814__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12538_ _06391_ _06392_ _06390_ vssd1 vssd1 vccd1 vccd1 _06395_ sky130_fd_sc_hd__o21ba_1
XFILLER_129_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10166__B _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12469_ net166 _05986_ net128 screen.register.currentXbus\[25\] vssd1 vssd1 vccd1
+ vccd1 _00871_ sky130_fd_sc_hd__a2bb2o_1
X_14208_ clknet_leaf_47_clk datapath.multiplication_module.multiplicand_i_n\[19\]
+ net1173 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_99_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11549__Y _05773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_810 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12381__B net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14139_ clknet_leaf_2_clk _00896_ net1065 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout409 _05733_ vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08790__A1 _03296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07593__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06961_ net991 _01666_ vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__and2_2
X_08700_ _03534_ _03535_ vssd1 vssd1 vccd1 vccd1 _03536_ sky130_fd_sc_hd__nor2_2
XANTENNA__12874__A0 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09680_ net633 _04513_ _04514_ _03824_ vssd1 vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__o22ai_2
X_06892_ _01707_ net929 vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__and2_1
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07345__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08631_ _03461_ _03464_ _02191_ vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__o21ba_1
XFILLER_39_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11217__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08562_ datapath.rf.registers\[27\]\[0\] net966 _01816_ vssd1 vssd1 vccd1 vccd1 _03398_
+ sky130_fd_sc_hd__and3_1
X_07513_ datapath.rf.registers\[11\]\[20\] net982 net939 vssd1 vssd1 vccd1 vccd1 _02349_
+ sky130_fd_sc_hd__and3_1
XFILLER_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08493_ datapath.rf.registers\[22\]\[1\] net964 net909 _01809_ vssd1 vssd1 vccd1
+ vccd1 _03329_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout156_A net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07444_ datapath.rf.registers\[9\]\[22\] net702 net679 datapath.rf.registers\[6\]\[22\]
+ _02275_ vssd1 vssd1 vccd1 vccd1 _02280_ sky130_fd_sc_hd__a221o_1
XFILLER_149_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07375_ _02194_ _02208_ _02209_ _02210_ vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__or4_1
XFILLER_129_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09114_ _03947_ _03949_ vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__nand2_2
XANTENNA__12448__A2_N _05944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09045_ net462 _03659_ vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout1232_A net1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12157__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold430 datapath.multiplication_module.multiplicand_i\[10\] vssd1 vssd1 vccd1 vccd1
+ net1778 sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 datapath.rf.registers\[31\]\[1\] vssd1 vssd1 vccd1 vccd1 net1789 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold452 datapath.rf.registers\[15\]\[26\] vssd1 vssd1 vccd1 vccd1 net1800 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout692_A _01824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold463 datapath.rf.registers\[15\]\[6\] vssd1 vssd1 vccd1 vccd1 net1811 sky130_fd_sc_hd__dlygate4sd3_1
Xhold474 datapath.rf.registers\[1\]\[21\] vssd1 vssd1 vccd1 vccd1 net1822 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08230__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold485 datapath.rf.registers\[19\]\[5\] vssd1 vssd1 vccd1 vccd1 net1833 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold496 datapath.rf.registers\[15\]\[30\] vssd1 vssd1 vccd1 vccd1 net1844 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout910 _01792_ vssd1 vssd1 vccd1 vccd1 net910 sky130_fd_sc_hd__buf_1
XANTENNA__07584__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout921 net923 vssd1 vssd1 vccd1 vccd1 net921 sky130_fd_sc_hd__clkbuf_4
Xfanout932 net933 vssd1 vssd1 vccd1 vccd1 net932 sky130_fd_sc_hd__buf_2
X_09947_ _04780_ _04782_ vssd1 vssd1 vccd1 vccd1 _04783_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout480_X net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout943 _01715_ vssd1 vssd1 vccd1 vccd1 net943 sky130_fd_sc_hd__buf_4
Xfanout954 _01710_ vssd1 vssd1 vccd1 vccd1 net954 sky130_fd_sc_hd__buf_4
XANTENNA_fanout957_A net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout578_X net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout965 net966 vssd1 vssd1 vccd1 vccd1 net965 sky130_fd_sc_hd__buf_2
Xfanout976 net979 vssd1 vssd1 vccd1 vccd1 net976 sky130_fd_sc_hd__buf_2
X_09878_ _04626_ _04645_ _04664_ net637 vssd1 vssd1 vccd1 vccd1 _04714_ sky130_fd_sc_hd__o31a_1
Xfanout987 net989 vssd1 vssd1 vccd1 vccd1 net987 sky130_fd_sc_hd__buf_2
Xhold1130 datapath.rf.registers\[17\]\[18\] vssd1 vssd1 vccd1 vccd1 net2478 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout998 _05789_ vssd1 vssd1 vccd1 vccd1 net998 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_51_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07336__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1141 datapath.rf.registers\[7\]\[20\] vssd1 vssd1 vccd1 vccd1 net2489 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1152 datapath.rf.registers\[9\]\[14\] vssd1 vssd1 vccd1 vccd1 net2500 sky130_fd_sc_hd__dlygate4sd3_1
X_08829_ net311 _03635_ _03641_ _03664_ vssd1 vssd1 vccd1 vccd1 _03665_ sky130_fd_sc_hd__o22a_1
Xhold1163 datapath.rf.registers\[30\]\[14\] vssd1 vssd1 vccd1 vccd1 net2511 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1174 datapath.rf.registers\[29\]\[17\] vssd1 vssd1 vccd1 vccd1 net2522 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout745_X net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11127__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1185 datapath.rf.registers\[9\]\[28\] vssd1 vssd1 vccd1 vccd1 net2533 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06729__B net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1196 datapath.rf.registers\[11\]\[8\] vssd1 vssd1 vccd1 vccd1 net2544 sky130_fd_sc_hd__dlygate4sd3_1
X_11840_ _05295_ _05760_ _05918_ _05819_ vssd1 vssd1 vccd1 vccd1 _05919_ sky130_fd_sc_hd__o31a_1
XFILLER_14_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08297__B1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_146_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_146_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11771_ net1526 net145 net140 _01855_ vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__a22o_1
X_13510_ clknet_leaf_23_clk _00320_ net1154 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_24_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10722_ net1680 _02960_ net572 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[8\]
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_24_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14490_ clknet_leaf_14_clk _01195_ net1102 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06847__B2 datapath.ru.latched_instruction\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_41_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13441_ clknet_leaf_46_clk _00251_ net1171 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10653_ net1013 _05471_ vssd1 vssd1 vccd1 vccd1 _05472_ sky130_fd_sc_hd__nand2b_1
XANTENNA__09797__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13372_ clknet_leaf_10_clk _00182_ net1073 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10584_ _02824_ _02876_ _02934_ _02980_ vssd1 vssd1 vccd1 vccd1 _05407_ sky130_fd_sc_hd__or4_1
Xclkload19 clknet_leaf_147_clk vssd1 vssd1 vccd1 vccd1 clkload19/X sky130_fd_sc_hd__clkbuf_8
X_12323_ _04872_ _05613_ net230 vssd1 vssd1 vccd1 vccd1 _06297_ sky130_fd_sc_hd__mux2_1
XFILLER_6_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12254_ net599 _06244_ _05898_ vssd1 vssd1 vccd1 vccd1 _06245_ sky130_fd_sc_hd__o21a_1
XFILLER_154_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11205_ net170 net2137 net423 vssd1 vssd1 vccd1 vccd1 _00257_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10206__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12185_ screen.counter.ct\[19\] _06165_ _06172_ screen.counter.ct\[20\] vssd1 vssd1
+ vccd1 vccd1 _06202_ sky130_fd_sc_hd__a31o_1
XANTENNA__07575__A2 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11136_ net182 net2012 net427 vssd1 vssd1 vccd1 vccd1 _00191_ sky130_fd_sc_hd__mux2_1
XANTENNA__11108__A0 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11067_ net182 net2153 net431 vssd1 vssd1 vccd1 vccd1 _00127_ sky130_fd_sc_hd__mux2_1
XFILLER_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07327__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10018_ _04800_ _04853_ vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__xnor2_1
XFILLER_76_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12928__Y _06555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14757_ screen.csx vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__clkbuf_1
X_11969_ screen.dcx _06010_ _06014_ vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_137_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_137_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13708_ clknet_leaf_133_clk _00518_ net1105 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_149_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14688_ clknet_leaf_135_clk _01393_ net1104 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13639_ clknet_leaf_145_clk _00449_ net1086 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07160_ datapath.rf.registers\[3\]\[28\] net773 net712 datapath.rf.registers\[11\]\[28\]
+ _01995_ vssd1 vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__a221o_1
XFILLER_145_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07091_ datapath.rf.registers\[24\]\[29\] net857 net793 datapath.rf.registers\[31\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_117_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11500__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08212__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout206 _05641_ vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__buf_1
Xfanout217 _05628_ vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__dlymetal6s2s_1
X_09801_ _03893_ _04636_ _03676_ vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__mux2_1
Xfanout228 _04712_ vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__clkbuf_2
XFILLER_87_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06712__A_N mmio.memload_or_instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload10_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout239 net240 vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__clkbuf_2
X_07993_ datapath.rf.registers\[3\]\[10\] net984 net928 vssd1 vssd1 vccd1 vccd1 _02829_
+ sky130_fd_sc_hd__and3_1
XFILLER_86_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09732_ net357 _04071_ vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__nand2_1
XFILLER_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06944_ _01591_ net891 vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__nand2_1
XANTENNA__07318__A2 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12311__A2 _04207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09663_ net357 _04163_ vssd1 vssd1 vccd1 vccd1 _04499_ sky130_fd_sc_hd__nand2_1
XANTENNA__10322__A1 _04207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06875_ _01630_ _01639_ _01657_ net961 vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__nor4_1
XANTENNA_fanout273_A _05564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08614_ _02636_ _03446_ _02637_ _02544_ _02590_ vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__a2111o_1
XPHY_EDGE_ROW_19_Left_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09594_ _03425_ _03558_ vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__xor2_1
XANTENNA__08279__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08545_ _03364_ _03378_ _03379_ _03380_ vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__nor4_1
XFILLER_36_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_128_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_128_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1182_A net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08818__A2 _03417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout159_X net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout538_A net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13162__S net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08764__B _01604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06829__A1 _01505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06829__B2 datapath.ru.latched_instruction\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11822__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08476_ datapath.rf.registers\[6\]\[1\] _01753_ net814 datapath.rf.registers\[23\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03312_ sky130_fd_sc_hd__a22o_1
XFILLER_51_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07427_ _02257_ _02259_ _02261_ _02262_ vssd1 vssd1 vccd1 vccd1 _02263_ sky130_fd_sc_hd__or4_1
XANTENNA__14648__RESET_B net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07358_ datapath.rf.registers\[2\]\[23\] net887 net845 datapath.rf.registers\[1\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__a22o_1
XFILLER_148_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08780__A net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09243__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10389__A1 _05223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_28_Left_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12506__S net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07289_ datapath.rf.registers\[0\]\[25\] net868 _02124_ vssd1 vssd1 vccd1 vccd1 _02125_
+ sky130_fd_sc_hd__o21a_4
XANTENNA__11410__S net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09028_ _03831_ _03832_ _03863_ vssd1 vssd1 vccd1 vccd1 _03864_ sky130_fd_sc_hd__a21o_1
XFILLER_156_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout695_X net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14290__Q datapath.rf.registers\[0\]\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold260 datapath.rf.registers\[8\]\[30\] vssd1 vssd1 vccd1 vccd1 net1608 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold271 datapath.rf.registers\[27\]\[17\] vssd1 vssd1 vccd1 vccd1 net1619 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09400__C1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold282 datapath.rf.registers\[1\]\[4\] vssd1 vssd1 vccd1 vccd1 net1630 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold293 datapath.rf.registers\[12\]\[14\] vssd1 vssd1 vccd1 vccd1 net1641 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout862_X net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout740 net741 vssd1 vssd1 vccd1 vccd1 net740 sky130_fd_sc_hd__buf_4
Xfanout751 _01804_ vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__buf_2
Xfanout762 net765 vssd1 vssd1 vccd1 vccd1 net762 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_148_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13990_ clknet_leaf_112_clk _00767_ net1219 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout773 _01798_ vssd1 vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_148_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout784 net785 vssd1 vssd1 vccd1 vccd1 net784 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07309__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout795 _01775_ vssd1 vssd1 vccd1 vccd1 net795 sky130_fd_sc_hd__clkbuf_8
X_12941_ net264 net2114 net395 vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_37_Left_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07562__C net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12872_ net275 net2512 net400 vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__mux2_1
XANTENNA__09403__X _04239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14611_ clknet_leaf_34_clk _01316_ net1128 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11823_ _01497_ net1017 net315 net335 datapath.ru.latched_instruction\[29\] vssd1
+ vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_119_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_119_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_45_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13072__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14542_ clknet_leaf_6_clk _01247_ net1067 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11813__A1 datapath.ru.latched_instruction\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11754_ net1494 net145 net140 _02680_ vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__a22o_1
XANTENNA__08019__X _02855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09482__A2 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10705_ net1473 _02876_ net571 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i_n\[10\]
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14473_ clknet_leaf_92_clk _01178_ net1234 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11685_ _05177_ net152 net151 net1432 vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_81_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13424_ clknet_leaf_25_clk _00234_ net1159 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12369__A2 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10636_ _05430_ _05454_ _05455_ vssd1 vssd1 vccd1 vccd1 _05456_ sky130_fd_sc_hd__a21bo_1
XANTENNA__08690__A _02705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload108 clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 clkload108/Y sky130_fd_sc_hd__inv_8
Xclkload119 clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 clkload119/Y sky130_fd_sc_hd__bufinv_16
Xmax_cap1046 _01532_ vssd1 vssd1 vccd1 vccd1 net1046 sky130_fd_sc_hd__buf_2
X_13355_ clknet_leaf_46_clk _00165_ net1171 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10567_ screen.register.currentXbus\[9\] screen.register.currentXbus\[8\] screen.register.currentXbus\[11\]
+ screen.register.currentXbus\[10\] vssd1 vssd1 vccd1 vccd1 _05391_ sky130_fd_sc_hd__or4_1
XANTENNA__06922__B net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11320__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12306_ _05585_ _06253_ vssd1 vssd1 vccd1 vccd1 _06285_ sky130_fd_sc_hd__nand2_1
XFILLER_143_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13286_ clknet_leaf_11_clk _00096_ net1083 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10498_ screen.controlBus\[5\] _05315_ _05327_ screen.controlBus\[4\] vssd1 vssd1
+ vccd1 vccd1 _05328_ sky130_fd_sc_hd__or4bb_1
XFILLER_142_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12450__A1_N net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12237_ _06233_ _06234_ vssd1 vssd1 vccd1 vccd1 _00774_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_112_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12168_ _01424_ _06163_ _06170_ _06191_ vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__a31o_1
XANTENNA__13953__RESET_B net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11119_ net264 net2032 net427 vssd1 vssd1 vccd1 vccd1 _00174_ sky130_fd_sc_hd__mux2_1
XFILLER_111_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12099_ screen.register.currentXbus\[7\] net1000 _05757_ screen.register.currentYbus\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06137_ sky130_fd_sc_hd__a22o_1
XANTENNA__09026__A _03850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput6 DAT_I[13] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
XFILLER_49_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10304__A1 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06660_ _01494_ _01495_ _01498_ datapath.ru.latched_instruction\[29\] _01496_ vssd1
+ vssd1 vccd1 vccd1 _01499_ sky130_fd_sc_hd__o221a_1
XANTENNA__07181__B1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07720__A2 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11562__Y _05786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06591_ columns.count\[10\] _01431_ vssd1 vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__nand2_1
XANTENNA__12387__A _05944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08584__B _03419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08330_ datapath.rf.registers\[25\]\[4\] net726 net687 datapath.rf.registers\[31\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03166_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_119_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08261_ datapath.rf.registers\[4\]\[5\] net864 _03095_ _03096_ vssd1 vssd1 vccd1
+ vccd1 _03097_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_15_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07212_ _02026_ _02047_ vssd1 vssd1 vccd1 vccd1 _02048_ sky130_fd_sc_hd__nor2_1
XANTENNA__09696__A net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08192_ _03015_ _03024_ _03027_ net782 datapath.rf.registers\[0\]\[7\] vssd1 vssd1
+ vccd1 vccd1 _03028_ sky130_fd_sc_hd__o32a_4
XFILLER_119_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07143_ _01964_ _01972_ _01976_ _01978_ vssd1 vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_99_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09630__C1 _03613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11230__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07787__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08984__B2 _03818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07074_ _01889_ _01909_ vssd1 vssd1 vccd1 vccd1 _01910_ sky130_fd_sc_hd__nand2_1
XFILLER_134_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10354__B net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1028_A net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07539__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout390_A net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13157__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout488_A _06552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07663__B net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07976_ datapath.rf.registers\[12\]\[11\] net756 net704 datapath.rf.registers\[9\]\[11\]
+ _02811_ vssd1 vssd1 vccd1 vccd1 _02812_ sky130_fd_sc_hd__a221o_1
XFILLER_142_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09715_ _03535_ net623 _03536_ net906 vssd1 vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__a2bb2o_1
X_06927_ datapath.rf.registers\[7\]\[31\] net817 _01761_ _01762_ net872 vssd1 vssd1
+ vccd1 vccd1 _01763_ sky130_fd_sc_hd__a2111o_1
XFILLER_74_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12996__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09646_ net370 _04290_ vssd1 vssd1 vccd1 vccd1 _04482_ sky130_fd_sc_hd__nand2_1
XFILLER_83_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06858_ datapath.ru.latched_instruction\[29\] _01594_ _01614_ datapath.ru.latched_instruction\[12\]
+ vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__a22o_1
XANTENNA__07172__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08775__A _01610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09577_ net460 _04351_ _04412_ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__a21oi_1
X_06789_ _01576_ _01584_ _01624_ vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__nor3_1
XANTENNA_fanout822_A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout443_X net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1185_X net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08494__B net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11405__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08528_ datapath.rf.registers\[24\]\[0\] net858 net834 datapath.rf.registers\[30\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__a22o_1
XANTENNA__07475__B2 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08459_ _03293_ _03294_ vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout610_X net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout708_X net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11470_ net2070 net193 net406 vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__mux2_1
XFILLER_51_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10421_ _03262_ _03321_ net441 vssd1 vssd1 vccd1 vccd1 _05257_ sky130_fd_sc_hd__mux2_1
XFILLER_109_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07778__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13140_ net1684 net263 net383 vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__mux2_1
X_10352_ datapath.PC\[10\] net1249 _05184_ _05187_ vssd1 vssd1 vccd1 vccd1 _05188_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07557__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13071_ net2545 net276 net388 vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__mux2_1
XFILLER_151_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10832__X _05588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10283_ datapath.PC\[6\] _03734_ datapath.PC\[7\] vssd1 vssd1 vccd1 vccd1 _05119_
+ sky130_fd_sc_hd__o21ai_1
X_12022_ screen.register.currentYbus\[2\] _06018_ _06019_ screen.register.currentYbus\[10\]
+ _06064_ vssd1 vssd1 vccd1 vccd1 _06065_ sky130_fd_sc_hd__a221o_1
XFILLER_151_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13067__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_45_Left_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08021__Y _02857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout570 net571 vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13973_ clknet_leaf_105_clk _00751_ net1224 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[16\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_74_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12924_ net1582 net178 net485 vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__mux2_1
XFILLER_46_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08685__A _02612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07702__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12855_ net196 net1946 net488 vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__mux2_1
XANTENNA__11315__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06917__B net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11806_ _01480_ net1017 net315 net335 datapath.ru.latched_instruction\[12\] vssd1
+ vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12786_ net212 net1845 net494 vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__mux2_1
XANTENNA__11798__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14525_ clknet_leaf_144_clk _01230_ net1085 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11737_ net25 net1036 _05889_ net2230 vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_54_Left_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14456_ clknet_leaf_4_clk _01161_ net1070 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11668_ _01405_ _05291_ _05883_ vssd1 vssd1 vccd1 vccd1 _05884_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_12_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06933__A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13407_ clknet_leaf_12_clk _00217_ net1082 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10619_ net38 _05380_ _05434_ net37 vssd1 vssd1 vccd1 vccd1 _05439_ sky130_fd_sc_hd__and4b_1
X_14387_ clknet_leaf_36_clk _01092_ net1135 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11599_ _05297_ _05298_ _05821_ _05822_ vssd1 vssd1 vccd1 vccd1 _05823_ sky130_fd_sc_hd__or4bb_1
XANTENNA__11050__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07769__A2 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13338_ clknet_leaf_3_clk _00148_ net1076 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13269_ clknet_leaf_129_clk _00079_ net1117 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_63_Left_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07830_ datapath.rf.registers\[16\]\[14\] net739 net723 datapath.rf.registers\[18\]\[14\]
+ _02664_ vssd1 vssd1 vccd1 vccd1 _02666_ sky130_fd_sc_hd__a221o_1
XANTENNA__06744__A3 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07761_ datapath.rf.registers\[17\]\[15\] net850 net805 datapath.rf.registers\[28\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02597_ sky130_fd_sc_hd__a22o_1
XFILLER_49_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09500_ _03552_ _03554_ vssd1 vssd1 vccd1 vccd1 _04336_ sky130_fd_sc_hd__xnor2_1
X_06712_ mmio.memload_or_instruction\[24\] mmio.memload_or_instruction\[26\] mmio.memload_or_instruction\[25\]
+ mmio.memload_or_instruction\[23\] vssd1 vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__and4bb_1
X_07692_ datapath.rf.registers\[13\]\[17\] net693 net681 datapath.rf.registers\[6\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__a22o_1
XANTENNA__07154__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09694__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09431_ net339 _04048_ _04266_ vssd1 vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__a21oi_1
X_06643_ net1288 net1283 datapath.ru.latched_instruction\[12\] mmio.memload_or_instruction\[12\]
+ vssd1 vssd1 vccd1 vccd1 _01482_ sky130_fd_sc_hd__or4b_1
XFILLER_37_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11225__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09362_ _04092_ _04197_ net374 vssd1 vssd1 vccd1 vccd1 _04198_ sky130_fd_sc_hd__mux2_1
X_06574_ datapath.rf.registers\[0\]\[28\] vssd1 vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__inv_2
XANTENNA__08882__X _03718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08313_ datapath.rf.registers\[0\]\[4\] net866 _03134_ _03148_ vssd1 vssd1 vccd1
+ vccd1 _03149_ sky130_fd_sc_hd__o22ai_4
XFILLER_32_170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09293_ net455 _04100_ _04101_ vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__and3_1
XANTENNA_11 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout236_A _05616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08244_ net560 _03078_ vssd1 vssd1 vccd1 vccd1 _03080_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_31_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14013__CLK clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07658__B net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08175_ datapath.rf.registers\[14\]\[7\] net776 net712 datapath.rf.registers\[11\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout403_A _06549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07126_ datapath.rf.registers\[19\]\[28\] net855 net844 datapath.rf.registers\[25\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__a22o_1
XFILLER_118_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07057_ datapath.rf.registers\[8\]\[30\] net696 net677 datapath.rf.registers\[29\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__a22o_1
XANTENNA__13804__RESET_B net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout772_A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout393_X net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08185__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07393__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07932__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06735__A3 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12269__A1 _05002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout560_X net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07959_ net874 _02792_ _02793_ _02794_ vssd1 vssd1 vccd1 vccd1 _02795_ sky130_fd_sc_hd__or4_1
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout658_X net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09134__A1 _03667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11924__A _02283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08001__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10970_ _05705_ _05704_ net655 _01443_ vssd1 vssd1 vccd1 vccd1 _05706_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_44_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09629_ net376 _03988_ _03984_ net332 vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__a211o_1
XFILLER_71_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout825_X net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11135__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12640_ net498 _06479_ _06480_ net502 datapath.mulitply_result\[21\] vssd1 vssd1
+ vccd1 vccd1 _00931_ sky130_fd_sc_hd__a32o_1
XANTENNA__10974__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12571_ _06415_ _06416_ _06417_ vssd1 vssd1 vccd1 vccd1 _06423_ sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_50_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_61_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14310_ clknet_leaf_93_clk _01015_ net1212 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[30\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_156_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11522_ _01420_ screen.register.xFill3 _01421_ screen.register.cFill3 net659 vssd1
+ vssd1 vccd1 vccd1 _05747_ sky130_fd_sc_hd__o221a_4
XANTENNA__10546__Y datapath.ack_mul vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14241_ clknet_leaf_124_clk datapath.multiplication_module.multiplier_i_n\[9\] net1214
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i\[9\] sky130_fd_sc_hd__dfrtp_1
X_11453_ net2619 net275 net408 vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__mux2_1
XANTENNA__08948__A1 _02126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10404_ datapath.PC\[0\] _05238_ net1240 vssd1 vssd1 vccd1 vccd1 _05240_ sky130_fd_sc_hd__mux2_2
X_14172_ clknet_leaf_55_clk _00927_ net1174 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_11384_ net2376 net284 net412 vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__mux2_1
X_13123_ net178 net2180 net472 vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__mux2_1
XFILLER_124_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10335_ net1040 _05168_ _05170_ net635 vssd1 vssd1 vccd1 vccd1 _05171_ sky130_fd_sc_hd__a211o_1
XANTENNA__13545__RESET_B net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ net196 net1849 net476 vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__mux2_1
X_10266_ net1043 _05101_ vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__nor2_1
XFILLER_105_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08399__B net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12005_ screen.register.currentYbus\[9\] _05776_ net996 screen.register.currentXbus\[25\]
+ _06048_ vssd1 vssd1 vccd1 vccd1 _06049_ sky130_fd_sc_hd__a221o_1
XANTENNA__08176__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10197_ _04881_ _05032_ net230 vssd1 vssd1 vccd1 vccd1 _05033_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07384__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07923__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13956_ clknet_leaf_103_clk _00734_ net1225 vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07136__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06928__A _01630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07687__A1 datapath.rf.registers\[0\]\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12907_ net2059 net268 net484 vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__mux2_1
X_13887_ clknet_leaf_73_clk _00691_ net1250 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[31\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_17_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11045__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12838_ net280 net2508 net488 vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__mux2_1
XFILLER_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10884__S net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12769_ net295 net1827 net494 vssd1 vssd1 vccd1 vccd1 _01022_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_41_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__10443__B1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14508_ clknet_leaf_14_clk _01213_ net1103 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09310__Y _04146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput20 DAT_I[26] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
XFILLER_147_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput31 DAT_I[7] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
X_14439_ clknet_leaf_137_clk _01144_ net1089 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_96_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold804 datapath.rf.registers\[3\]\[6\] vssd1 vssd1 vccd1 vccd1 net2152 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06950__X _01786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold815 datapath.rf.registers\[14\]\[10\] vssd1 vssd1 vccd1 vccd1 net2163 sky130_fd_sc_hd__dlygate4sd3_1
Xhold826 datapath.rf.registers\[17\]\[3\] vssd1 vssd1 vccd1 vccd1 net2174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold837 datapath.rf.registers\[31\]\[4\] vssd1 vssd1 vccd1 vccd1 net2185 sky130_fd_sc_hd__dlygate4sd3_1
Xhold848 datapath.rf.registers\[8\]\[19\] vssd1 vssd1 vccd1 vccd1 net2196 sky130_fd_sc_hd__dlygate4sd3_1
X_09980_ _04815_ _04814_ vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__and2b_1
Xhold859 datapath.rf.registers\[23\]\[16\] vssd1 vssd1 vccd1 vccd1 net2207 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08931_ net372 _03766_ _03627_ vssd1 vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08167__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08862_ net320 _03693_ _03697_ net322 vssd1 vssd1 vccd1 vccd1 _03698_ sky130_fd_sc_hd__a211o_1
XANTENNA__08102__B _01707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07813_ datapath.rf.registers\[16\]\[14\] net861 net805 datapath.rf.registers\[28\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_127_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08793_ _01666_ _03358_ _03615_ vssd1 vssd1 vccd1 vccd1 _03629_ sky130_fd_sc_hd__mux2_1
XFILLER_84_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07744_ datapath.rf.registers\[24\]\[16\] net766 net726 datapath.rf.registers\[25\]\[16\]
+ _02579_ vssd1 vssd1 vccd1 vccd1 _02580_ sky130_fd_sc_hd__a221o_1
XANTENNA__07941__B net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07127__B1 _01721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08875__A0 _03205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07660__C net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07675_ datapath.rf.registers\[18\]\[17\] net791 _02493_ _02495_ _02507_ vssd1 vssd1
+ vccd1 vccd1 _02511_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_36_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09414_ net454 _04187_ _04248_ net349 vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__a211o_1
X_06626_ net1287 net1282 datapath.ru.latched_instruction\[24\] mmio.memload_or_instruction\[24\]
+ vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__or4b_1
XFILLER_41_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09345_ _03575_ _04179_ vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout520_A net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1262_A _00004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout618_A net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08772__B net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_32_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_21_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09276_ net339 _03851_ _04111_ net322 vssd1 vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__a211o_1
X_08227_ datapath.rf.registers\[10\]\[6\] net706 net660 datapath.rf.registers\[5\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03063_ sky130_fd_sc_hd__a22o_1
XANTENNA__10095__A net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout406_X net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08158_ datapath.rf.registers\[25\]\[7\] net843 net814 datapath.rf.registers\[23\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02994_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout987_A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07109_ datapath.rf.registers\[22\]\[29\] net734 net707 datapath.rf.registers\[10\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__a22o_1
XANTENNA__07602__B2 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08089_ datapath.rf.registers\[3\]\[9\] net772 net670 datapath.rf.registers\[21\]\[9\]
+ _02924_ vssd1 vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__a221o_1
X_10120_ net1043 _03746_ _04955_ net902 vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__a31o_1
XANTENNA__10542__B datapath.multiplication_module.multiplier_i\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout775_X net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_99_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_99_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08158__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10051_ _04823_ _04886_ vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__and2_1
XFILLER_76_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07905__A2 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout942_X net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13810_ clknet_leaf_73_clk _00619_ net1242 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07851__B net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13741_ clknet_leaf_50_clk _00551_ net1176 vssd1 vssd1 vccd1 vccd1 mmio.key_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_3_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08866__A0 _02705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10953_ _05689_ _05690_ vssd1 vssd1 vccd1 vccd1 _05691_ sky130_fd_sc_hd__or2_1
XFILLER_44_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08330__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13672_ clknet_leaf_63_clk _00482_ net1233 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10884_ _04023_ _05631_ net903 vssd1 vssd1 vccd1 vccd1 _05632_ sky130_fd_sc_hd__mux2_2
X_12623_ datapath.mulitply_result\[19\] datapath.multiplication_module.multiplicand_i\[19\]
+ vssd1 vssd1 vccd1 vccd1 _06466_ sky130_fd_sc_hd__and2_1
XANTENNA__13080__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_23_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_8_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12554_ _06407_ _06408_ vssd1 vssd1 vccd1 vccd1 _06409_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11505_ net188 net1950 net511 vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__mux2_1
XFILLER_12_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12485_ net283 net1958 net508 vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__mux2_1
XFILLER_156_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14224_ clknet_leaf_42_clk _00945_ net1144 vssd1 vssd1 vccd1 vccd1 columns.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_138_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11436_ net192 net2158 net514 vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__mux2_1
XANTENNA__06770__X _01607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10728__A1 _02660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14155_ clknet_leaf_90_clk _00910_ net1239 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11367_ net199 net1566 net518 vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__mux2_1
XANTENNA__06930__B net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13106_ net268 net1766 net471 vssd1 vssd1 vccd1 vccd1 _01348_ sky130_fd_sc_hd__mux2_1
XFILLER_3_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10318_ _04836_ _04843_ vssd1 vssd1 vccd1 vccd1 _05154_ sky130_fd_sc_hd__and2b_1
X_14086_ clknet_leaf_109_clk _00852_ net1220 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11298_ net199 net2126 net523 vssd1 vssd1 vccd1 vccd1 _00346_ sky130_fd_sc_hd__mux2_1
X_13037_ net278 net2188 net477 vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__mux2_1
X_10249_ _01417_ _05084_ net1252 vssd1 vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__mux2_2
Xfanout1140 net1143 vssd1 vssd1 vccd1 vccd1 net1140 sky130_fd_sc_hd__clkbuf_4
Xfanout1151 net1152 vssd1 vssd1 vccd1 vccd1 net1151 sky130_fd_sc_hd__clkbuf_2
XFILLER_79_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1162 net1186 vssd1 vssd1 vccd1 vccd1 net1162 sky130_fd_sc_hd__buf_2
Xfanout1173 net1178 vssd1 vssd1 vccd1 vccd1 net1173 sky130_fd_sc_hd__clkbuf_4
XFILLER_67_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_109_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1184 net1185 vssd1 vssd1 vccd1 vccd1 net1184 sky130_fd_sc_hd__clkbuf_2
Xfanout1195 net1196 vssd1 vssd1 vccd1 vccd1 net1195 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07109__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12379__B net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13939_ clknet_leaf_110_clk _00717_ net1222 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13426__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_62_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08321__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07460_ datapath.rf.registers\[16\]\[21\] net860 net793 datapath.rf.registers\[31\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__a22o_1
XFILLER_34_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07391_ datapath.rf.registers\[26\]\[23\] net778 net668 datapath.rf.registers\[21\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_14_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__11503__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09130_ net353 _03842_ _03845_ vssd1 vssd1 vccd1 vccd1 _03966_ sky130_fd_sc_hd__or3_1
XANTENNA_clkbuf_leaf_77_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09061_ net449 _03702_ vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_100_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_120_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07776__X _02612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08012_ datapath.rf.registers\[4\]\[10\] net865 _02834_ _02835_ _02838_ vssd1 vssd1
+ vccd1 vccd1 _02848_ sky130_fd_sc_hd__a2111o_1
XFILLER_129_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09034__B1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold601 datapath.rf.registers\[6\]\[26\] vssd1 vssd1 vccd1 vccd1 net1949 sky130_fd_sc_hd__dlygate4sd3_1
Xhold612 datapath.rf.registers\[8\]\[10\] vssd1 vssd1 vccd1 vccd1 net1960 sky130_fd_sc_hd__dlygate4sd3_1
Xhold623 datapath.rf.registers\[17\]\[17\] vssd1 vssd1 vccd1 vccd1 net1971 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08388__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold634 datapath.rf.registers\[18\]\[1\] vssd1 vssd1 vccd1 vccd1 net1982 sky130_fd_sc_hd__dlygate4sd3_1
Xhold645 datapath.rf.registers\[25\]\[28\] vssd1 vssd1 vccd1 vccd1 net1993 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11392__A1 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold656 datapath.rf.registers\[21\]\[9\] vssd1 vssd1 vccd1 vccd1 net2004 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07596__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold667 datapath.rf.registers\[17\]\[16\] vssd1 vssd1 vccd1 vccd1 net2015 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold678 datapath.rf.registers\[9\]\[5\] vssd1 vssd1 vccd1 vccd1 net2026 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07060__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09963_ _04763_ _04798_ vssd1 vssd1 vccd1 vccd1 _04799_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_135_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold689 datapath.rf.registers\[24\]\[4\] vssd1 vssd1 vccd1 vccd1 net2037 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08914_ datapath.PC\[28\] _03749_ vssd1 vssd1 vccd1 vccd1 _03750_ sky130_fd_sc_hd__or2_1
XFILLER_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09894_ datapath.PC\[19\] net604 _04728_ vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__or3_1
XFILLER_131_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1010_A net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07348__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_15_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1301 mmio.memload_or_instruction\[12\] vssd1 vssd1 vccd1 vccd1 net2649 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08845_ _02126_ _02170_ net444 vssd1 vssd1 vccd1 vccd1 _03681_ sky130_fd_sc_hd__mux2_1
XANTENNA__11695__A2 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout470_A net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08560__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07671__B net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08776_ _03611_ vssd1 vssd1 vccd1 vccd1 _03612_ sky130_fd_sc_hd__inv_2
XFILLER_150_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07727_ datapath.rf.registers\[20\]\[16\] net839 _02546_ _02551_ _02562_ vssd1 vssd1
+ vccd1 vccd1 _02563_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10104__C1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout735_A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07658_ datapath.rf.registers\[8\]\[17\] net955 _01712_ vssd1 vssd1 vccd1 vccd1 _02494_
+ sky130_fd_sc_hd__and3_1
X_06609_ net1286 net1281 mmio.memload_or_instruction\[4\] vssd1 vssd1 vccd1 vccd1
+ _01448_ sky130_fd_sc_hd__or3_1
Xclkbuf_4_8_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_8_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_13_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12509__S net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout523_X net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07589_ datapath.rf.registers\[7\]\[19\] net673 net670 datapath.rf.registers\[21\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout902_A net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11413__S net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09328_ _03931_ _04163_ net361 vssd1 vssd1 vccd1 vccd1 _04164_ sky130_fd_sc_hd__mux2_1
XFILLER_40_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09273__B1 _03770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09259_ net370 _03956_ _04093_ net327 vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__a211oi_1
XFILLER_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07686__X _02522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09025__B1 _03859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12270_ datapath.PC\[4\] net308 _06256_ _06258_ vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__a22o_1
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11221_ net255 net2067 net529 vssd1 vssd1 vccd1 vccd1 _00271_ sky130_fd_sc_hd__mux2_1
XANTENNA__08379__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07587__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11152_ net268 net1991 net532 vssd1 vssd1 vccd1 vccd1 _00205_ sky130_fd_sc_hd__mux2_1
XFILLER_1_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07565__C net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10103_ _03915_ _04606_ _04624_ _03864_ _03830_ vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_8_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11083_ net270 net1798 net536 vssd1 vssd1 vccd1 vccd1 _00140_ sky130_fd_sc_hd__mux2_1
XFILLER_110_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07339__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input31_A DAT_I[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10034_ _04729_ _04730_ vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__and2b_1
XFILLER_76_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13075__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08396__C _01744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06909__C _01630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11985_ screen.register.currentXbus\[24\] net996 net995 screen.register.currentXbus\[0\]
+ _06029_ vssd1 vssd1 vccd1 vccd1 _06030_ sky130_fd_sc_hd__a221o_1
XFILLER_84_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08303__A2 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13724_ clknet_leaf_8_clk _00534_ net1071 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10936_ _01497_ net620 _05675_ _05676_ vssd1 vssd1 vccd1 vccd1 _05677_ sky130_fd_sc_hd__a22o_2
XFILLER_16_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10867_ datapath.PC\[20\] _05611_ vssd1 vssd1 vccd1 vccd1 _05617_ sky130_fd_sc_hd__and2_1
X_13655_ clknet_leaf_126_clk _00465_ net1206 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11323__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12606_ datapath.mulitply_result\[16\] datapath.multiplication_module.multiplicand_i\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06452_ sky130_fd_sc_hd__or2_1
X_13586_ clknet_leaf_32_clk _00396_ net1123 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10798_ net277 net1903 net543 vssd1 vssd1 vccd1 vccd1 _00011_ sky130_fd_sc_hd__mux2_1
XANTENNA__10949__B2 _01477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10447__B _05270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12537_ net500 _06393_ _06394_ net504 datapath.mulitply_result\[4\] vssd1 vssd1 vccd1
+ vccd1 _00914_ sky130_fd_sc_hd__a32o_1
XFILLER_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12468_ net166 _05984_ net128 screen.register.currentXbus\[24\] vssd1 vssd1 vccd1
+ vccd1 _00870_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09567__A1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14207_ clknet_leaf_47_clk datapath.multiplication_module.multiplicand_i_n\[18\]
+ net1173 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_11419_ net275 net2553 net516 vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__mux2_1
X_12399_ _05956_ net158 vssd1 vssd1 vccd1 vccd1 _06347_ sky130_fd_sc_hd__nor2_1
XFILLER_153_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14138_ clknet_leaf_9_clk _00895_ net1080 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07042__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08790__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14069_ clknet_leaf_111_clk _00836_ net1196 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_06960_ net968 net909 _01795_ vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__and3_2
XFILLER_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_3_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_8
X_06891_ net961 _01657_ net980 vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__and3b_1
XFILLER_121_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08630_ _03463_ _03465_ vssd1 vssd1 vccd1 vccd1 _03466_ sky130_fd_sc_hd__nand2_1
XANTENNA__08542__A2 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08561_ datapath.rf.registers\[31\]\[0\] net966 _01825_ vssd1 vssd1 vccd1 vccd1 _03397_
+ sky130_fd_sc_hd__and3_1
X_07512_ datapath.rf.registers\[29\]\[20\] net973 net917 vssd1 vssd1 vccd1 vccd1 _02348_
+ sky130_fd_sc_hd__and3_1
X_08492_ datapath.rf.registers\[12\]\[1\] net757 _03325_ _03326_ _03327_ vssd1 vssd1
+ vccd1 vccd1 _03328_ sky130_fd_sc_hd__a2111o_1
X_07443_ datapath.rf.registers\[15\]\[22\] net664 net660 datapath.rf.registers\[5\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__a22o_1
XFILLER_11_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11233__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout149_A net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07374_ datapath.rf.registers\[20\]\[23\] net839 _02193_ _02195_ _02199_ vssd1 vssd1
+ vccd1 vccd1 _02210_ sky130_fd_sc_hd__a2111o_1
XFILLER_148_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09113_ _03824_ _03948_ net616 vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__o21a_1
XFILLER_129_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1058_A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09044_ net331 _03879_ net312 vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_135_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07281__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09558__A1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold420 datapath.rf.registers\[24\]\[6\] vssd1 vssd1 vccd1 vccd1 net1768 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07666__B net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09558__B2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold431 datapath.rf.registers\[9\]\[4\] vssd1 vssd1 vccd1 vccd1 net1779 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07569__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1225_A net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold442 datapath.rf.registers\[16\]\[16\] vssd1 vssd1 vccd1 vccd1 net1790 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold453 datapath.rf.registers\[1\]\[14\] vssd1 vssd1 vccd1 vccd1 net1801 sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 datapath.rf.registers\[7\]\[18\] vssd1 vssd1 vccd1 vccd1 net1812 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12999__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold475 datapath.rf.registers\[20\]\[0\] vssd1 vssd1 vccd1 vccd1 net1823 sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 datapath.rf.registers\[2\]\[30\] vssd1 vssd1 vccd1 vccd1 net1834 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout900 net903 vssd1 vssd1 vccd1 vccd1 net900 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout685_A net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold497 datapath.rf.registers\[23\]\[22\] vssd1 vssd1 vccd1 vccd1 net1845 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout911 net913 vssd1 vssd1 vccd1 vccd1 net911 sky130_fd_sc_hd__clkbuf_2
Xfanout922 net923 vssd1 vssd1 vccd1 vccd1 net922 sky130_fd_sc_hd__buf_1
XANTENNA__09881__B net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09946_ datapath.PC\[1\] _03322_ _03323_ vssd1 vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__or3_1
Xfanout933 _01725_ vssd1 vssd1 vccd1 vccd1 net933 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08778__A _03601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout944 _01715_ vssd1 vssd1 vccd1 vccd1 net944 sky130_fd_sc_hd__buf_2
XFILLER_131_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout955 net956 vssd1 vssd1 vccd1 vccd1 net955 sky130_fd_sc_hd__clkbuf_4
Xfanout966 net967 vssd1 vssd1 vccd1 vccd1 net966 sky130_fd_sc_hd__buf_2
Xfanout977 net979 vssd1 vssd1 vccd1 vccd1 net977 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10325__C1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09877_ net633 _04710_ _03670_ vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__a21o_1
Xhold1120 datapath.rf.registers\[10\]\[23\] vssd1 vssd1 vccd1 vccd1 net2468 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout852_A _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout473_X net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08497__B net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout988 net989 vssd1 vssd1 vccd1 vccd1 net988 sky130_fd_sc_hd__clkbuf_4
Xfanout999 _05788_ vssd1 vssd1 vccd1 vccd1 net999 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11408__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1131 datapath.rf.registers\[3\]\[16\] vssd1 vssd1 vccd1 vccd1 net2479 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08533__A2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1142 screen.register.currentYbus\[31\] vssd1 vssd1 vccd1 vccd1 net2490 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1153 datapath.rf.registers\[3\]\[15\] vssd1 vssd1 vccd1 vccd1 net2501 sky130_fd_sc_hd__dlygate4sd3_1
X_08828_ _03642_ _03661_ net347 net650 vssd1 vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__o31a_1
Xhold1164 datapath.rf.registers\[2\]\[9\] vssd1 vssd1 vccd1 vccd1 net2512 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07741__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1175 screen.register.currentYbus\[15\] vssd1 vssd1 vccd1 vccd1 net2523 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1186 datapath.rf.registers\[29\]\[21\] vssd1 vssd1 vccd1 vccd1 net2534 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1197 datapath.rf.registers\[5\]\[9\] vssd1 vssd1 vccd1 vccd1 net2545 sky130_fd_sc_hd__dlygate4sd3_1
X_08759_ _03487_ _03489_ _03594_ vssd1 vssd1 vccd1 vccd1 _03595_ sky130_fd_sc_hd__and3_1
XFILLER_72_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout738_X net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11770_ net1502 net145 net140 _01908_ vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__a22o_1
XFILLER_14_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10721_ net1915 _03008_ net572 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[7\]
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_24_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout905_X net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11143__S net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13440_ clknet_leaf_136_clk _00250_ net1090 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10652_ button\[1\] _01435_ vssd1 vssd1 vccd1 vccd1 _05471_ sky130_fd_sc_hd__nand2_1
XANTENNA__10982__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13371_ clknet_leaf_37_clk _00181_ net1138 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10835__X _05590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10583_ _02634_ _02680_ _02725_ _02771_ vssd1 vssd1 vccd1 vccd1 _05406_ sky130_fd_sc_hd__or4_1
X_12322_ _06294_ _06296_ datapath.PC\[18\] net310 vssd1 vssd1 vccd1 vccd1 _00797_
+ sky130_fd_sc_hd__a2bb2o_1
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12253_ _01590_ _01670_ _05901_ vssd1 vssd1 vccd1 vccd1 _06244_ sky130_fd_sc_hd__a21oi_1
XFILLER_123_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11204_ net175 net2047 net424 vssd1 vssd1 vccd1 vccd1 _00256_ sky130_fd_sc_hd__mux2_1
X_12184_ _06166_ _06172_ _06178_ vssd1 vssd1 vccd1 vccd1 _06201_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_71_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11135_ net176 net2533 net428 vssd1 vssd1 vccd1 vccd1 _00190_ sky130_fd_sc_hd__mux2_1
XFILLER_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14177__RESET_B net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12305__B1 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07980__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11066_ net179 net1873 net433 vssd1 vssd1 vccd1 vccd1 _00126_ sky130_fd_sc_hd__mux2_1
XANTENNA__08040__X _02876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10316__C1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11318__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10017_ _04756_ _04757_ vssd1 vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08200__B net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_86_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14756_ net1291 vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_102_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11968_ _06002_ _06005_ _06013_ _05848_ vssd1 vssd1 vccd1 vccd1 _06014_ sky130_fd_sc_hd__o211a_1
XANTENNA__09312__A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13707_ clknet_leaf_57_clk _00517_ net1167 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10919_ _03865_ _05661_ net902 vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__mux2_1
X_11899_ screen.register.currentYbus\[14\] net161 vssd1 vssd1 vccd1 vccd1 _05963_
+ sky130_fd_sc_hd__nand2_1
X_14687_ clknet_leaf_3_clk _01392_ net1077 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11053__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13638_ clknet_leaf_29_clk _00448_ net1133 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_146_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07248__C1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13569_ clknet_leaf_46_clk _00379_ net1147 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07799__B1 _01787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07090_ datapath.rf.registers\[21\]\[29\] net815 _01923_ _01924_ _01925_ vssd1 vssd1
+ vccd1 vccd1 _01926_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_117_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07015__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09800_ _03685_ _03680_ net449 vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__mux2_1
Xfanout207 net208 vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__clkbuf_2
Xfanout218 net221 vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout229 net230 vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__clkbuf_4
X_07992_ datapath.rf.registers\[20\]\[10\] net959 net925 vssd1 vssd1 vccd1 vccd1 _02828_
+ sky130_fd_sc_hd__and3_1
XFILLER_87_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07971__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06943_ datapath.rf.registers\[0\]\[31\] net866 _01752_ _01778_ vssd1 vssd1 vccd1
+ vccd1 _01779_ sky130_fd_sc_hd__o22ai_4
X_09731_ _03571_ _04566_ net580 vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__o21ai_1
XFILLER_140_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11228__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08515__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09662_ _04414_ _04419_ net354 vssd1 vssd1 vccd1 vccd1 _04498_ sky130_fd_sc_hd__mux2_1
X_06874_ _01657_ net961 vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__nor2_1
XFILLER_95_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08885__X _03721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07723__B1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08613_ _02544_ _02589_ vssd1 vssd1 vccd1 vccd1 _03449_ sky130_fd_sc_hd__nand2b_1
X_09593_ _04396_ _04428_ vssd1 vssd1 vccd1 vccd1 _04429_ sky130_fd_sc_hd__nor2_1
XFILLER_131_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08544_ datapath.rf.registers\[6\]\[0\] _01753_ net816 datapath.rf.registers\[21\]\[0\]
+ _03362_ vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__a221o_1
XFILLER_82_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08475_ datapath.rf.registers\[8\]\[1\] net878 net835 datapath.rf.registers\[30\]\[1\]
+ _03310_ vssd1 vssd1 vccd1 vccd1 _03311_ sky130_fd_sc_hd__a221o_1
XANTENNA__10368__A _05085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1175_A net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07426_ datapath.rf.registers\[17\]\[22\] net849 net801 datapath.rf.registers\[3\]\[22\]
+ _02249_ vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__a221o_1
XFILLER_51_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09779__A1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07357_ datapath.rf.registers\[4\]\[23\] net957 net932 vssd1 vssd1 vccd1 vccd1 _02193_
+ sky130_fd_sc_hd__and3_1
XFILLER_149_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08780__B net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07677__A net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07254__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07288_ _02114_ _02119_ _02123_ vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__or3_4
XFILLER_152_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09027_ net608 _03829_ _03862_ net556 vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__o211ai_1
XFILLER_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09892__A _01585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07006__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold250 datapath.rf.registers\[23\]\[19\] vssd1 vssd1 vccd1 vccd1 net1598 sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 datapath.rf.registers\[6\]\[3\] vssd1 vssd1 vccd1 vccd1 net1609 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold272 datapath.rf.registers\[29\]\[27\] vssd1 vssd1 vccd1 vccd1 net1620 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout688_X net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold283 datapath.rf.registers\[6\]\[13\] vssd1 vssd1 vccd1 vccd1 net1631 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11927__A net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold294 datapath.rf.registers\[28\]\[2\] vssd1 vssd1 vccd1 vccd1 net1642 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout730 _01811_ vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__clkbuf_8
Xfanout741 _01808_ vssd1 vssd1 vccd1 vccd1 net741 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06765__B2 _01466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_130_Right_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout752 _01804_ vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__buf_4
X_09929_ datapath.PC\[8\] _02981_ vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_148_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout763 net765 vssd1 vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_148_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout774 _01796_ vssd1 vssd1 vccd1 vccd1 net774 sky130_fd_sc_hd__buf_4
XANTENNA_fanout855_X net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11138__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout785 _01791_ vssd1 vssd1 vccd1 vccd1 net785 sky130_fd_sc_hd__clkbuf_4
Xfanout796 net798 vssd1 vssd1 vccd1 vccd1 net796 sky130_fd_sc_hd__clkbuf_8
X_12940_ net269 net2618 net396 vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__mux2_1
XFILLER_19_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10977__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12871_ net279 net2549 net400 vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__mux2_1
X_14610_ clknet_leaf_32_clk _01315_ net1123 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09467__A0 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11822_ net1045 net1014 net313 net333 datapath.ru.latched_instruction\[28\] vssd1
+ vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__a32o_1
XFILLER_27_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11753_ net1481 net146 net141 _02725_ vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__a22o_1
X_14541_ clknet_leaf_132_clk _01246_ net1113 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10704_ net1446 _02934_ net570 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i_n\[9\]
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11684_ _05106_ net152 net151 net1456 vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__a22o_1
XANTENNA__07493__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14472_ clknet_leaf_64_clk _01177_ net1235 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_81_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10635_ _05428_ _05443_ vssd1 vssd1 vccd1 vccd1 _05455_ sky130_fd_sc_hd__nor2_1
X_13423_ clknet_leaf_25_clk _00233_ net1138 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_128_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload109 clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 clkload109/Y sky130_fd_sc_hd__inv_8
X_13354_ clknet_leaf_61_clk _00164_ net1165 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xmax_cap1047 _01456_ vssd1 vssd1 vccd1 vccd1 net1047 sky130_fd_sc_hd__buf_1
X_10566_ screen.register.currentXbus\[1\] screen.register.currentXbus\[0\] screen.register.currentXbus\[3\]
+ screen.register.currentXbus\[2\] vssd1 vssd1 vccd1 vccd1 _05390_ sky130_fd_sc_hd__or4_1
X_12305_ net890 _04861_ net190 vssd1 vssd1 vccd1 vccd1 _06284_ sky130_fd_sc_hd__a21o_1
X_13285_ clknet_leaf_141_clk _00095_ net1188 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10497_ screen.controlBus\[7\] screen.controlBus\[6\] _05326_ vssd1 vssd1 vccd1 vccd1
+ _05327_ sky130_fd_sc_hd__nor3_1
XFILLER_108_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12236_ net2414 _06232_ net602 vssd1 vssd1 vccd1 vccd1 _06234_ sky130_fd_sc_hd__o21ai_1
XFILLER_108_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12167_ _06162_ net567 _06179_ net1273 vssd1 vssd1 vccd1 vccd1 _06191_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_112_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06756__A1 _01477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11118_ net268 net2197 net428 vssd1 vssd1 vccd1 vccd1 _00173_ sky130_fd_sc_hd__mux2_1
X_12098_ screen.register.currentXbus\[23\] _05769_ _05837_ screen.register.currentYbus\[23\]
+ _06135_ vssd1 vssd1 vccd1 vccd1 _06136_ sky130_fd_sc_hd__a221o_1
XANTENNA__11048__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11049_ net266 net2264 net432 vssd1 vssd1 vccd1 vccd1 _00109_ sky130_fd_sc_hd__mux2_1
Xinput7 DAT_I[14] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10887__S net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06590_ columns.count\[7\] columns.count\[6\] columns.count\[9\] columns.count\[8\]
+ vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__and4_1
XFILLER_64_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12387__B net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08130__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08260_ datapath.rf.registers\[9\]\[5\] net885 net829 datapath.rf.registers\[14\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03096_ sky130_fd_sc_hd__a22o_1
XANTENNA__07484__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08881__A _01610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07211_ net610 _02045_ _01787_ vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__o21ai_2
XFILLER_20_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08191_ _03017_ _03019_ _03020_ _03026_ vssd1 vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__or4_1
XFILLER_146_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07142_ datapath.rf.registers\[9\]\[28\] _01716_ net835 datapath.rf.registers\[30\]\[28\]
+ _01977_ vssd1 vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__a221o_1
XANTENNA__07497__A _02311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07236__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07073_ net613 _01908_ net565 vssd1 vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__a21o_1
XANTENNA__08105__B net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14028__RESET_B net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11740__B2 _03417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07663__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07975_ datapath.rf.registers\[30\]\[11\] net760 net752 datapath.rf.registers\[28\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__a22o_1
XANTENNA__10370__B net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout383_A net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06926_ datapath.rf.registers\[2\]\[31\] net887 net879 datapath.rf.registers\[10\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__a22o_1
X_09714_ _03663_ _04541_ _04543_ net574 vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__o211a_1
X_06857_ datapath.ru.latched_instruction\[20\] net992 _01692_ vssd1 vssd1 vccd1 vccd1
+ _01693_ sky130_fd_sc_hd__a21oi_1
X_09645_ net647 _04480_ _03770_ vssd1 vssd1 vccd1 vccd1 _04481_ sky130_fd_sc_hd__o21a_1
XFILLER_16_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1292_A _01436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout269_X net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout648_A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08775__B _01614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09576_ net457 _04214_ _04215_ vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__and3_1
X_06788_ _01579_ _01587_ vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__nand2_1
XFILLER_24_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08527_ datapath.rf.registers\[7\]\[0\] net942 net936 vssd1 vssd1 vccd1 vccd1 _03363_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout815_A net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout436_X net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1178_X net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08458_ net614 _03265_ vssd1 vssd1 vccd1 vccd1 _03294_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_46_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07409_ datapath.rf.registers\[22\]\[22\] net954 net921 vssd1 vssd1 vccd1 vccd1 _02245_
+ sky130_fd_sc_hd__and3_1
X_08389_ _03218_ _03220_ _03222_ _03224_ vssd1 vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__or4_2
XFILLER_7_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11421__S net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10420_ net362 _04325_ _04441_ net371 vssd1 vssd1 vccd1 vccd1 _05256_ sky130_fd_sc_hd__o211a_1
XANTENNA__07227__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10351_ net222 _05186_ net1292 vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__a21o_1
X_13070_ net1907 net278 net389 vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__mux2_1
X_10282_ datapath.PC\[7\] _04495_ net468 vssd1 vssd1 vccd1 vccd1 _05118_ sky130_fd_sc_hd__mux2_1
XFILLER_133_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08188__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12021_ screen.register.currentYbus\[26\] _05757_ _05769_ screen.register.currentXbus\[18\]
+ vssd1 vssd1 vccd1 vccd1 _06064_ sky130_fd_sc_hd__a22o_1
XFILLER_151_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout560 _03057_ vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09137__C1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout571 _05367_ vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13972_ clknet_leaf_105_clk _00750_ net1224 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_76_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12923_ net2574 net187 net483 vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__mux2_1
XANTENNA__07699__C1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13083__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12854_ net202 net2112 net486 vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11805_ _01474_ net1017 net315 net335 datapath.ru.latched_instruction\[11\] vssd1
+ vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__a32o_1
X_12785_ net216 net2101 net494 vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__mux2_1
XANTENNA__08112__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_1_Left_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07869__X _02705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14524_ clknet_leaf_10_clk _01229_ net1073 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11736_ net23 net1034 net1024 net2282 vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__o22a_1
XANTENNA__06773__X _01610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07466__A2 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14455_ clknet_leaf_124_clk _01160_ net1208 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11667_ mmio.wishbone.curr_state\[0\] _05289_ vssd1 vssd1 vccd1 vccd1 _05883_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_12_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11331__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06933__B net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13406_ clknet_leaf_148_clk _00216_ net1060 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10618_ _05431_ net1013 _05437_ vssd1 vssd1 vccd1 vccd1 _05438_ sky130_fd_sc_hd__or3_1
X_11598_ screen.counter.ct\[7\] net1279 screen.counter.ct\[15\] screen.counter.ct\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05822_ sky130_fd_sc_hd__and4b_1
X_14386_ clknet_leaf_32_clk _01091_ net1126 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09612__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10549_ keypad.debounce.debounce\[2\] _05374_ _05375_ vssd1 vssd1 vccd1 vccd1 _05376_
+ sky130_fd_sc_hd__and3_1
XFILLER_128_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13337_ clknet_leaf_31_clk _00147_ net1122 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13268_ clknet_leaf_93_clk _00078_ net1212 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09915__A1 _01613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12219_ screen.counter.currentCt\[9\] screen.counter.currentCt\[10\] _06219_ vssd1
+ vssd1 vccd1 vccd1 _06223_ sky130_fd_sc_hd__and3_1
XFILLER_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13199_ clknet_leaf_26_clk _00009_ net1135 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_151_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07926__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07760_ datapath.rf.registers\[14\]\[15\] net831 net808 datapath.rf.registers\[27\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02596_ sky130_fd_sc_hd__a22o_1
XFILLER_65_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12278__A2 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06711_ _01541_ _01542_ _01549_ vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__nor3_1
X_07691_ datapath.rf.registers\[24\]\[17\] net768 net752 datapath.rf.registers\[28\]\[17\]
+ _02524_ vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__a221o_1
XFILLER_65_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11506__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09430_ net339 _04052_ vssd1 vssd1 vccd1 vccd1 _04266_ sky130_fd_sc_hd__nor2_1
X_06642_ mmio.memload_or_instruction\[12\] net1050 vssd1 vssd1 vccd1 vccd1 _01481_
+ sky130_fd_sc_hd__nand2_1
XFILLER_53_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09361_ net364 _04124_ _04196_ vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__a21oi_1
X_06573_ datapath.ru.latched_instruction\[23\] vssd1 vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__inv_2
XANTENNA__11789__A1 _05747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08103__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08312_ _03136_ _03137_ _03142_ _03147_ vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__or4_1
XANTENNA__07457__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09292_ net330 _04127_ net311 vssd1 vssd1 vccd1 vccd1 _04128_ sky130_fd_sc_hd__a21o_1
XFILLER_21_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_12 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08243_ _03078_ vssd1 vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout131_A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07939__B net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06843__B _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout229_A net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11241__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08174_ datapath.rf.registers\[13\]\[7\] net693 net685 datapath.rf.registers\[27\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03010_ sky130_fd_sc_hd__a22o_1
XANTENNA__07658__C _01712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10213__A1 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07125_ datapath.rf.registers\[21\]\[28\] net945 net926 vssd1 vssd1 vccd1 vccd1 _01961_
+ sky130_fd_sc_hd__and3_1
XFILLER_137_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1040_A net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1138_A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07056_ datapath.rf.registers\[18\]\[30\] net724 net673 datapath.rf.registers\[7\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__a22o_1
XANTENNA__09367__C1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout598_A net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07917__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08489__C _01823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout386_X net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12800__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07958_ datapath.rf.registers\[17\]\[11\] net851 _02777_ _02778_ _02788_ vssd1 vssd1
+ vccd1 vccd1 _02794_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12269__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06909_ net962 _01639_ _01630_ _01656_ vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__and4b_1
XANTENNA_fanout932_A net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07889_ datapath.rf.registers\[0\]\[13\] net784 _02724_ vssd1 vssd1 vccd1 vccd1 _02725_
+ sky130_fd_sc_hd__o21a_2
XANTENNA__11416__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07145__B2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09628_ net329 _04230_ _04462_ _04463_ vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_48_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07696__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout720_X net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09559_ _04393_ _04394_ vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout818_X net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12977__A0 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12570_ _06420_ _06421_ vssd1 vssd1 vccd1 vccd1 _06422_ sky130_fd_sc_hd__nand2_1
XANTENNA__07448__A2 _02283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11521_ _05360_ _05743_ _05745_ net1010 _05304_ vssd1 vssd1 vccd1 vccd1 _05746_ sky130_fd_sc_hd__a32oi_1
XANTENNA__14632__RESET_B net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09767__D _04600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11151__S net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06753__B _01579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14240_ clknet_leaf_124_clk datapath.multiplication_module.multiplier_i_n\[8\] net1214
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i\[8\] sky130_fd_sc_hd__dfrtp_1
X_11452_ net1661 net279 net409 vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__mux2_1
XFILLER_149_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07568__C net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10204__A1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10403_ datapath.PC\[0\] _03384_ vssd1 vssd1 vccd1 vccd1 _05239_ sky130_fd_sc_hd__or2_1
X_14171_ clknet_leaf_55_clk _00926_ net1179 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10843__X _05597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10990__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11383_ net1678 net290 net410 vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__mux2_1
XANTENNA__10755__A2 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10334_ _03740_ _05169_ net1040 vssd1 vssd1 vccd1 vccd1 _05170_ sky130_fd_sc_hd__a21oi_1
X_13122_ net185 net1830 net473 vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__mux2_1
XANTENNA__07081__B1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07620__A2 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13078__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13053_ net199 net1664 net474 vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__mux2_1
X_10265_ datapath.PC\[13\] _04272_ net467 vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_76_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07908__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12004_ screen.register.currentYbus\[25\] _05786_ net999 screen.register.currentXbus\[9\]
+ _05781_ vssd1 vssd1 vccd1 vccd1 _06048_ sky130_fd_sc_hd__a221o_1
XANTENNA__08399__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10196_ _04878_ _04880_ vssd1 vssd1 vccd1 vccd1 _05032_ sky130_fd_sc_hd__or2_1
XFILLER_79_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08696__A _02805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout390 net391 vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__buf_4
X_13955_ clknet_leaf_104_clk _00733_ net1225 vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__dfrtp_1
XFILLER_47_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06928__B _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11326__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload7_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12906_ net1579 net273 net484 vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__mux2_1
XFILLER_46_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13886_ clknet_leaf_74_clk _00690_ net1242 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[30\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_17_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13915__SET_B net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06895__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12837_ net282 net1717 net488 vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__mux2_1
XFILLER_62_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07439__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12768_ net300 net2060 net495 vssd1 vssd1 vccd1 vccd1 _01021_ sky130_fd_sc_hd__mux2_1
XFILLER_30_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14507_ clknet_leaf_59_clk _01212_ net1168 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11719_ net5 net1034 net1024 net2649 vssd1 vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__o22a_1
XFILLER_147_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12699_ net2578 net503 net499 _06529_ vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__a22o_1
XANTENNA__11061__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput10 DAT_I[17] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
X_14438_ clknet_leaf_11_clk _01143_ net1083 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput21 DAT_I[27] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
Xinput32 DAT_I[8] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_1
XFILLER_128_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold805 datapath.rf.registers\[8\]\[29\] vssd1 vssd1 vccd1 vccd1 net2153 sky130_fd_sc_hd__dlygate4sd3_1
X_14369_ clknet_leaf_25_clk _01074_ net1159 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold816 datapath.rf.registers\[25\]\[21\] vssd1 vssd1 vccd1 vccd1 net2164 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07072__B1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold827 datapath.rf.registers\[10\]\[9\] vssd1 vssd1 vccd1 vccd1 net2175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold838 datapath.rf.registers\[26\]\[8\] vssd1 vssd1 vccd1 vccd1 net2186 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07611__A2 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold849 datapath.rf.registers\[9\]\[11\] vssd1 vssd1 vccd1 vccd1 net2197 sky130_fd_sc_hd__dlygate4sd3_1
X_08930_ net368 _03765_ _03764_ vssd1 vssd1 vccd1 vccd1 _03766_ sky130_fd_sc_hd__a21boi_2
XFILLER_115_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08861_ net344 _03682_ net338 _03696_ vssd1 vssd1 vccd1 vccd1 _03697_ sky130_fd_sc_hd__o211a_1
XANTENNA__08102__C net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07812_ datapath.rf.registers\[1\]\[14\] net846 net795 datapath.rf.registers\[31\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02648_ sky130_fd_sc_hd__a22o_1
X_08792_ net972 _03359_ _03615_ vssd1 vssd1 vccd1 vccd1 _03628_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_127_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07743_ datapath.rf.registers\[2\]\[16\] net742 net664 datapath.rf.registers\[15\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02579_ sky130_fd_sc_hd__a22o_1
XFILLER_38_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07941__C net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08324__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11236__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout179_A _05670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07674_ datapath.rf.registers\[29\]\[17\] net797 net794 datapath.rf.registers\[31\]\[17\]
+ _02497_ vssd1 vssd1 vccd1 vccd1 _02510_ sky130_fd_sc_hd__a221o_1
XANTENNA__08893__X _03729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07678__A2 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08875__A1 _03263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06625_ net1288 net1284 mmio.memload_or_instruction\[24\] vssd1 vssd1 vccd1 vccd1
+ _01464_ sky130_fd_sc_hd__or3b_1
X_09413_ net454 _04187_ _04248_ vssd1 vssd1 vccd1 vccd1 _04249_ sky130_fd_sc_hd__a21o_1
XANTENNA__10928__X _05670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09344_ _03446_ _04179_ vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__xor2_1
XFILLER_32_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09275_ net339 _03856_ vssd1 vssd1 vccd1 vccd1 _04111_ sky130_fd_sc_hd__nor2_1
XANTENNA__07669__B net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout513_A _05735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08226_ _03060_ _03061_ vssd1 vssd1 vccd1 vccd1 _03062_ sky130_fd_sc_hd__or2_1
XFILLER_20_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08157_ datapath.rf.registers\[14\]\[7\] net830 net791 datapath.rf.registers\[18\]\[7\]
+ _02988_ vssd1 vssd1 vccd1 vccd1 _02993_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1043_X net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07108_ datapath.rf.registers\[18\]\[29\] net723 net688 datapath.rf.registers\[31\]\[29\]
+ _01943_ vssd1 vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__a221o_1
XANTENNA__07063__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08088_ datapath.rf.registers\[2\]\[9\] net744 net685 datapath.rf.registers\[27\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02924_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout882_A net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07039_ _01864_ _01868_ _01870_ _01874_ vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__or4_1
XFILLER_115_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10050_ net1264 datapath.PC\[25\] net594 vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11698__B1 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout670_X net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout768_X net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09760__C1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_82_Left_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout935_X net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11146__S net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08315__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13740_ clknet_leaf_51_clk _00550_ net1181 vssd1 vssd1 vccd1 vccd1 mmio.key_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_723 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08866__A1 _02751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10952_ _01649_ _03264_ vssd1 vssd1 vccd1 vccd1 _05690_ sky130_fd_sc_hd__or2_1
XFILLER_73_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13671_ clknet_leaf_145_clk _00481_ net1087 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10985__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10883_ _05629_ _05630_ vssd1 vssd1 vccd1 vccd1 _05631_ sky130_fd_sc_hd__nor2_1
X_12622_ net498 _06464_ _06465_ net502 net2531 vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__a32o_1
XANTENNA__09815__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06764__A _01593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12553_ _06402_ _06403_ _06400_ vssd1 vssd1 vccd1 vccd1 _06408_ sky130_fd_sc_hd__o21a_1
XFILLER_8_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11504_ net195 net1929 net510 vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__mux2_1
XANTENNA__07841__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12484_ net290 net2073 net506 vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_91_Left_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11669__X _05885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14223_ clknet_leaf_42_clk _00944_ net1144 vssd1 vssd1 vccd1 vccd1 columns.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_22_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11435_ _05653_ net2605 net516 vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__mux2_1
XANTENNA__10189__B1 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07054__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14154_ clknet_leaf_77_clk net1374 net1246 vssd1 vssd1 vccd1 vccd1 datapath.pc_module.i_ack2
+ sky130_fd_sc_hd__dfrtp_1
X_11366_ net203 net2208 net519 vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__mux2_1
XFILLER_99_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13105_ net271 net2590 net471 vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__mux2_1
X_10317_ net892 _05148_ _05152_ net229 vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__o211a_1
X_14085_ clknet_leaf_109_clk _00851_ net1220 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11297_ net204 net2305 net522 vssd1 vssd1 vccd1 vccd1 _00345_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08203__B net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13036_ net284 net2191 net476 vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__mux2_1
X_10248_ _05076_ _05083_ net227 vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__mux2_1
Xfanout1130 net1153 vssd1 vssd1 vccd1 vccd1 net1130 sky130_fd_sc_hd__clkbuf_2
Xfanout1141 net1143 vssd1 vssd1 vccd1 vccd1 net1141 sky130_fd_sc_hd__clkbuf_4
Xfanout1152 net1153 vssd1 vssd1 vccd1 vccd1 net1152 sky130_fd_sc_hd__clkbuf_2
X_10179_ net641 _04607_ _05014_ _05013_ net225 vssd1 vssd1 vccd1 vccd1 _05015_ sky130_fd_sc_hd__a311oi_1
Xfanout1163 net1166 vssd1 vssd1 vccd1 vccd1 net1163 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06939__A net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1174 net1178 vssd1 vssd1 vccd1 vccd1 net1174 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_109_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1185 net1186 vssd1 vssd1 vccd1 vccd1 net1185 sky130_fd_sc_hd__clkbuf_2
Xfanout1196 net1204 vssd1 vssd1 vccd1 vccd1 net1196 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11056__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13938_ clknet_leaf_109_clk _00716_ net1218 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10895__S net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13869_ clknet_leaf_74_clk _00673_ net1242 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_23_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07390_ datapath.rf.registers\[30\]\[23\] net758 net750 datapath.rf.registers\[28\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__a22o_1
XFILLER_31_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10416__A1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09282__A1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08085__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09282__B2 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09060_ _03895_ vssd1 vssd1 vccd1 vccd1 _03896_ sky130_fd_sc_hd__inv_2
XANTENNA__07293__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07832__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06961__X _01797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08011_ datapath.rf.registers\[11\]\[10\] net884 net834 datapath.rf.registers\[30\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02847_ sky130_fd_sc_hd__a22o_1
XFILLER_129_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold602 datapath.rf.registers\[19\]\[27\] vssd1 vssd1 vccd1 vccd1 net1950 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold613 datapath.rf.registers\[29\]\[16\] vssd1 vssd1 vccd1 vccd1 net1961 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold624 datapath.rf.registers\[3\]\[3\] vssd1 vssd1 vccd1 vccd1 net1972 sky130_fd_sc_hd__dlygate4sd3_1
Xhold635 datapath.rf.registers\[29\]\[11\] vssd1 vssd1 vccd1 vccd1 net1983 sky130_fd_sc_hd__dlygate4sd3_1
Xhold646 datapath.rf.registers\[12\]\[17\] vssd1 vssd1 vccd1 vccd1 net1994 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08793__A0 _01666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold657 datapath.rf.registers\[3\]\[5\] vssd1 vssd1 vccd1 vccd1 net2005 sky130_fd_sc_hd__dlygate4sd3_1
Xhold668 datapath.rf.registers\[17\]\[20\] vssd1 vssd1 vccd1 vccd1 net2016 sky130_fd_sc_hd__dlygate4sd3_1
Xhold679 datapath.rf.registers\[24\]\[22\] vssd1 vssd1 vccd1 vccd1 net2027 sky130_fd_sc_hd__dlygate4sd3_1
X_09962_ net1267 _02935_ _04794_ _04795_ _04765_ vssd1 vssd1 vccd1 vccd1 _04798_ sky130_fd_sc_hd__a221o_1
X_08913_ net1263 datapath.PC\[27\] _03748_ vssd1 vssd1 vccd1 vccd1 _03749_ sky130_fd_sc_hd__or3_1
XANTENNA__09337__A2 _03718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_139_Left_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09893_ net604 _04728_ datapath.PC\[19\] vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__o21a_1
XANTENNA__12341__A1 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout296_A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1302 screen.register.currentXbus\[2\] vssd1 vssd1 vccd1 vccd1 net2650 sky130_fd_sc_hd__dlygate4sd3_1
X_08844_ _02026_ _02070_ net447 vssd1 vssd1 vccd1 vccd1 _03680_ sky130_fd_sc_hd__mux2_1
XANTENNA__07671__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08775_ _01610_ _01614_ _01618_ vssd1 vssd1 vccd1 vccd1 _03611_ sky130_fd_sc_hd__or3b_2
XANTENNA_fanout463_A _03149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07726_ datapath.rf.registers\[21\]\[16\] net815 _02548_ _02549_ _02550_ vssd1 vssd1
+ vccd1 vccd1 _02562_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_0_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08848__A1 _01647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07657_ datapath.rf.registers\[10\]\[17\] net984 net937 vssd1 vssd1 vccd1 vccd1 _02493_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout630_A _01706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout728_A _01812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06608_ datapath.ru.latched_instruction\[13\] _01446_ vssd1 vssd1 vccd1 vccd1 _01447_
+ sky130_fd_sc_hd__xor2_1
X_07588_ datapath.rf.registers\[16\]\[19\] net740 net732 datapath.rf.registers\[19\]\[19\]
+ _02423_ vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__a221o_1
XFILLER_40_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09327_ _04070_ _04162_ net355 vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__mux2_1
XANTENNA__09273__A1 _01609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout516_X net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07967__X _02803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07284__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09258_ net370 _03956_ _04093_ vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_153_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08209_ datapath.rf.registers\[12\]\[6\] net826 _03034_ _03044_ vssd1 vssd1 vccd1
+ vccd1 _03045_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_153_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09189_ _03458_ _04024_ vssd1 vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__xnor2_2
XANTENNA__09025__A1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11220_ net264 net2020 net529 vssd1 vssd1 vccd1 vccd1 _00270_ sky130_fd_sc_hd__mux2_1
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout885_X net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08784__B1 _03613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11151_ net270 net2391 net532 vssd1 vssd1 vccd1 vccd1 _00204_ sky130_fd_sc_hd__mux2_1
XFILLER_134_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10102_ net893 _04935_ _04937_ vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_73_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11082_ net276 net2342 net536 vssd1 vssd1 vccd1 vccd1 _00139_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08536__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10033_ _04733_ _04811_ vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input24_A DAT_I[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12096__B1 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06909__D _01656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11984_ screen.register.currentYbus\[0\] _05778_ net999 screen.register.currentXbus\[8\]
+ _06028_ vssd1 vssd1 vccd1 vccd1 _06029_ sky130_fd_sc_hd__a221o_1
X_13723_ clknet_leaf_36_clk _00533_ net1136 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10935_ datapath.mulitply_result\[29\] net615 net652 vssd1 vssd1 vccd1 vccd1 _05676_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_104_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13091__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13654_ clknet_leaf_140_clk _00464_ net1095 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10866_ net235 net2110 net543 vssd1 vssd1 vccd1 vccd1 _00021_ sky130_fd_sc_hd__mux2_1
XFILLER_90_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12605_ datapath.mulitply_result\[16\] datapath.multiplication_module.multiplicand_i\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06451_ sky130_fd_sc_hd__nand2_1
XANTENNA__08067__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13585_ clknet_leaf_40_clk _00395_ net1140 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10797_ _05557_ _05556_ net655 _01536_ vssd1 vssd1 vccd1 vccd1 _05558_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__07275__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12536_ _06390_ _06391_ _06392_ vssd1 vssd1 vccd1 vccd1 _06394_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07814__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13947__RESET_B net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12467_ net164 _05982_ net126 screen.register.currentXbus\[23\] vssd1 vssd1 vccd1
+ vccd1 _00869_ sky130_fd_sc_hd__a2bb2o_1
XPHY_EDGE_ROW_144_Right_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14206_ clknet_leaf_55_clk datapath.multiplication_module.multiplicand_i_n\[17\]
+ net1179 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_144_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11418_ net281 net1921 net516 vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__mux2_1
X_12398_ net1383 net132 _06346_ vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__a21o_1
XFILLER_152_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14137_ clknet_leaf_4_clk _00894_ net1069 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11349_ net290 net2209 net519 vssd1 vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__mux2_1
XFILLER_125_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14068_ clknet_leaf_111_clk _00835_ net1196 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_140_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09724__C1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13019_ net1539 net199 net390 vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__mux2_1
X_06890_ net957 net931 vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__and2_2
XFILLER_67_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10334__B1 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12087__B1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08560_ datapath.rf.registers\[30\]\[0\] net761 _03393_ _03394_ _03395_ vssd1 vssd1
+ vccd1 vccd1 _03396_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08884__A _01613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07511_ datapath.rf.registers\[20\]\[20\] net957 net922 vssd1 vssd1 vccd1 vccd1 _02347_
+ sky130_fd_sc_hd__and3_1
X_08491_ datapath.rf.registers\[30\]\[1\] net966 net909 _01795_ vssd1 vssd1 vccd1
+ vccd1 _03327_ sky130_fd_sc_hd__and4_1
X_07442_ datapath.rf.registers\[8\]\[22\] net694 net675 datapath.rf.registers\[29\]\[22\]
+ _02277_ vssd1 vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__a221o_1
XFILLER_63_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07373_ datapath.rf.registers\[22\]\[23\] net821 _02196_ _02197_ _02198_ vssd1 vssd1
+ vccd1 vccd1 _02209_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09255__A1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09112_ _03461_ _03497_ vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__xor2_1
XFILLER_148_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09043_ net327 _03877_ _03623_ vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_135_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07947__B net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout309_A _06246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12011__B1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold410 datapath.rf.registers\[25\]\[3\] vssd1 vssd1 vccd1 vccd1 net1758 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_111_Right_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold421 datapath.rf.registers\[16\]\[17\] vssd1 vssd1 vccd1 vccd1 net1769 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07666__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_6_0_clk_X clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold432 datapath.rf.registers\[15\]\[7\] vssd1 vssd1 vccd1 vccd1 net1780 sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 datapath.rf.registers\[5\]\[10\] vssd1 vssd1 vccd1 vccd1 net1791 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold454 datapath.mulitply_result\[11\] vssd1 vssd1 vccd1 vccd1 net1802 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_147_Left_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold465 datapath.rf.registers\[1\]\[24\] vssd1 vssd1 vccd1 vccd1 net1813 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08230__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1120_A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10092__C _03914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold476 datapath.rf.registers\[18\]\[28\] vssd1 vssd1 vccd1 vccd1 net1824 sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 datapath.rf.registers\[26\]\[22\] vssd1 vssd1 vccd1 vccd1 net1835 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout901 net902 vssd1 vssd1 vccd1 vccd1 net901 sky130_fd_sc_hd__buf_4
Xhold498 datapath.rf.registers\[24\]\[3\] vssd1 vssd1 vccd1 vccd1 net1846 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout912 net913 vssd1 vssd1 vccd1 vccd1 net912 sky130_fd_sc_hd__buf_1
X_09945_ datapath.PC\[0\] _03384_ vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__nand2_1
Xfanout923 _01739_ vssd1 vssd1 vccd1 vccd1 net923 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout934 net935 vssd1 vssd1 vccd1 vccd1 net934 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout945 net948 vssd1 vssd1 vccd1 vccd1 net945 sky130_fd_sc_hd__buf_4
Xfanout956 _01709_ vssd1 vssd1 vccd1 vccd1 net956 sky130_fd_sc_hd__clkbuf_2
X_09876_ net633 _04710_ _03670_ vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__a21oi_2
XFILLER_86_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout967 _01676_ vssd1 vssd1 vccd1 vccd1 net967 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11522__C1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1110 datapath.rf.registers\[9\]\[13\] vssd1 vssd1 vccd1 vccd1 net2458 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout978 net979 vssd1 vssd1 vccd1 vccd1 net978 sky130_fd_sc_hd__buf_1
Xhold1121 datapath.rf.registers\[18\]\[10\] vssd1 vssd1 vccd1 vccd1 net2469 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09191__B1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout989 _01650_ vssd1 vssd1 vccd1 vccd1 net989 sky130_fd_sc_hd__clkbuf_2
Xhold1132 datapath.rf.registers\[8\]\[20\] vssd1 vssd1 vccd1 vccd1 net2480 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08497__C _01823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08827_ net971 _03172_ _03643_ vssd1 vssd1 vccd1 vccd1 _03663_ sky130_fd_sc_hd__mux2_1
Xhold1143 datapath.rf.registers\[12\]\[2\] vssd1 vssd1 vccd1 vccd1 net2491 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout466_X net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout845_A _01737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1154 datapath.rf.registers\[9\]\[0\] vssd1 vssd1 vccd1 vccd1 net2502 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1165 datapath.mulitply_result\[14\] vssd1 vssd1 vccd1 vccd1 net2513 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1176 datapath.rf.registers\[13\]\[16\] vssd1 vssd1 vccd1 vccd1 net2524 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1187 datapath.rf.registers\[21\]\[15\] vssd1 vssd1 vccd1 vccd1 net2535 sky130_fd_sc_hd__dlygate4sd3_1
X_08758_ _03492_ _03494_ _03591_ _03490_ _03488_ vssd1 vssd1 vccd1 vccd1 _03594_ sky130_fd_sc_hd__a311o_1
Xhold1198 datapath.rf.registers\[8\]\[31\] vssd1 vssd1 vccd1 vccd1 net2546 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_156_Left_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07709_ _02522_ _02543_ vssd1 vssd1 vccd1 vccd1 _02545_ sky130_fd_sc_hd__or2_1
XFILLER_54_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08297__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout633_X net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08689_ _02705_ _02726_ vssd1 vssd1 vccd1 vccd1 _03525_ sky130_fd_sc_hd__nand2_1
XANTENNA__11424__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10720_ _03057_ net572 _05512_ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[6\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10651_ keypad.alpha _05470_ _05463_ vssd1 vssd1 vccd1 vccd1 keypad.decode.button_n\[0\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_9_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout800_X net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13370_ clknet_leaf_14_clk _00180_ net1079 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09797__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10582_ _05396_ _05399_ _05402_ _05404_ vssd1 vssd1 vccd1 vccd1 _05405_ sky130_fd_sc_hd__or4_1
X_12321_ _05606_ _06254_ _06295_ net191 vssd1 vssd1 vccd1 vccd1 _06296_ sky130_fd_sc_hd__o22a_1
XFILLER_126_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07009__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12252_ net1379 _06242_ _06243_ vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12002__B1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11203_ net181 net1947 net423 vssd1 vssd1 vccd1 vccd1 _00255_ sky130_fd_sc_hd__mux2_1
X_12183_ _06200_ _06198_ screen.counter.ct\[19\] vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__mux2_1
XFILLER_150_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_61_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11134_ net187 net2351 net427 vssd1 vssd1 vccd1 vccd1 _00189_ sky130_fd_sc_hd__mux2_1
XANTENNA__13086__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11065_ net186 datapath.rf.registers\[8\]\[27\] net431 vssd1 vssd1 vccd1 vccd1 _00125_
+ sky130_fd_sc_hd__mux2_1
XFILLER_48_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10016_ _04835_ _04851_ vssd1 vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_76_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08200__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12069__B1 _05786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06776__X _01613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14755_ net1291 vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_86_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11967_ _05999_ _06012_ _05819_ vssd1 vssd1 vccd1 vccd1 _06013_ sky130_fd_sc_hd__o21ai_1
XFILLER_44_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11334__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06936__B net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13706_ clknet_leaf_58_clk _00516_ net1168 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10918_ _05660_ vssd1 vssd1 vccd1 vccd1 _05661_ sky130_fd_sc_hd__inv_2
XANTENNA__07496__B1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14686_ clknet_leaf_1_clk _01391_ net1062 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11898_ net134 _05962_ _05961_ vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_leaf_134_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13637_ clknet_leaf_118_clk _00447_ net1192 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10849_ _05600_ _05601_ vssd1 vssd1 vccd1 vccd1 _05602_ sky130_fd_sc_hd__or2_1
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_14_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13568_ clknet_leaf_135_clk _00378_ net1090 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06952__A _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07799__A1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12519_ net500 _06378_ _06379_ net504 datapath.mulitply_result\[1\] vssd1 vssd1 vccd1
+ vccd1 _00911_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_117_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13499_ clknet_leaf_38_clk _00309_ net1145 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_149_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_29_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08212__A2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10761__X _05527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07420__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout208 _05700_ vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__buf_2
XFILLER_114_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout219 net221 vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__clkbuf_2
XFILLER_99_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07991_ _02804_ _02825_ vssd1 vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__and2_1
XANTENNA__11509__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_7_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_7_0_clk sky130_fd_sc_hd__clkbuf_8
X_09730_ _03531_ _03570_ _03530_ vssd1 vssd1 vccd1 vccd1 _04566_ sky130_fd_sc_hd__a21oi_1
X_06942_ _01757_ _01763_ _01770_ _01777_ vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__or4_1
X_09661_ _03564_ _03565_ vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__xor2_1
X_06873_ net980 _01656_ net961 vssd1 vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__nor3_1
XFILLER_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08612_ _02589_ _03447_ _02590_ vssd1 vssd1 vccd1 vccd1 _03448_ sky130_fd_sc_hd__o21bai_2
X_09592_ net630 _04397_ _04425_ _04427_ vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__o22ai_4
XFILLER_82_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08543_ datapath.rf.registers\[20\]\[0\] _01740_ net814 datapath.rf.registers\[23\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__a22o_1
XANTENNA__08279__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout161_A _05933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11244__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout259_A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07487__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08474_ datapath.rf.registers\[16\]\[1\] net862 net830 datapath.rf.registers\[14\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__a22o_1
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11822__A3 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07425_ datapath.rf.registers\[5\]\[22\] net819 _02246_ _02248_ _02260_ vssd1 vssd1
+ vccd1 vccd1 _02261_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_137_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1070_A net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10936__X _05677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout426_A _05716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07239__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07356_ datapath.rf.registers\[10\]\[23\] net879 net804 datapath.rf.registers\[28\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__a22o_1
XFILLER_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08780__C _03614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07287_ _02120_ _02121_ _02122_ vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_150_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08125__Y _02961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09026_ _03850_ _03854_ _03860_ _03861_ vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__or4b_1
XFILLER_156_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold240 datapath.rf.registers\[28\]\[1\] vssd1 vssd1 vccd1 vccd1 net1588 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12803__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold251 datapath.rf.registers\[19\]\[6\] vssd1 vssd1 vccd1 vccd1 net1599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 datapath.rf.registers\[7\]\[23\] vssd1 vssd1 vccd1 vccd1 net1610 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold273 datapath.rf.registers\[11\]\[0\] vssd1 vssd1 vccd1 vccd1 net1621 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11927__B screen.counter.ack vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold284 datapath.rf.registers\[7\]\[25\] vssd1 vssd1 vccd1 vccd1 net1632 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 datapath.rf.registers\[4\]\[18\] vssd1 vssd1 vccd1 vccd1 net1643 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout962_A _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout720 net721 vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__buf_4
XANTENNA__11419__S net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout731 _01811_ vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__buf_2
Xfanout742 net745 vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__buf_4
X_09928_ net1267 _02935_ vssd1 vssd1 vccd1 vccd1 _04764_ sky130_fd_sc_hd__nand2_1
Xfanout753 _01804_ vssd1 vssd1 vccd1 vccd1 net753 sky130_fd_sc_hd__buf_2
Xfanout764 net765 vssd1 vssd1 vccd1 vccd1 net764 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_148_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout775 _01796_ vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout786 net789 vssd1 vssd1 vccd1 vccd1 net786 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout750_X net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09859_ _03361_ _04678_ _03297_ _03360_ vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__o211a_1
Xfanout797 net798 vssd1 vssd1 vccd1 vccd1 net797 sky130_fd_sc_hd__buf_4
XFILLER_46_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout848_X net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12870_ net282 net2565 net400 vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__mux2_1
X_11821_ datapath.ru.latched_instruction\[27\] net335 net315 _01597_ vssd1 vssd1 vccd1
+ vccd1 _00687_ sky130_fd_sc_hd__a22o_1
XANTENNA__09467__A1 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11154__S net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07478__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14540_ clknet_leaf_134_clk _01245_ net1104 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_81_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11752_ net1466 net146 net141 _02771_ vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__a22o_1
XFILLER_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10703_ net1505 _02980_ net571 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i_n\[8\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA__10993__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14471_ clknet_leaf_145_clk _01176_ net1086 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11683_ _05146_ net152 net151 net1420 vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__a22o_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13422_ clknet_leaf_4_clk _00232_ net1069 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10634_ _05432_ _05433_ _05437_ vssd1 vssd1 vccd1 vccd1 _05454_ sky130_fd_sc_hd__or3_1
XANTENNA__06772__A _01575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13353_ clknet_leaf_92_clk _00163_ net1232 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xmax_cap1037 _05442_ vssd1 vssd1 vccd1 vccd1 net1037 sky130_fd_sc_hd__buf_1
X_10565_ screen.register.currentXbus\[5\] screen.register.currentXbus\[4\] screen.register.currentXbus\[7\]
+ screen.register.currentXbus\[6\] vssd1 vssd1 vccd1 vccd1 _05389_ sky130_fd_sc_hd__or4_1
XANTENNA__08442__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12304_ datapath.PC\[13\] net307 _06283_ _05099_ vssd1 vssd1 vccd1 vccd1 _00792_
+ sky130_fd_sc_hd__o22a_1
XFILLER_127_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13284_ clknet_leaf_18_clk _00094_ net1116 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10496_ screen.controlBus\[0\] screen.controlBus\[1\] screen.controlBus\[2\] screen.controlBus\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05326_ sky130_fd_sc_hd__or4_2
X_12235_ screen.counter.currentCt\[16\] _06232_ vssd1 vssd1 vccd1 vccd1 _06233_ sky130_fd_sc_hd__and2_1
XANTENNA__08699__A _02857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12166_ _06162_ net567 _06179_ _06190_ vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_112_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11329__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11117_ net272 net1644 net428 vssd1 vssd1 vccd1 vccd1 _00172_ sky130_fd_sc_hd__mux2_1
X_12097_ screen.register.currentYbus\[7\] _06018_ _06019_ screen.register.currentYbus\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06135_ sky130_fd_sc_hd__a22o_1
X_11048_ net270 net1960 net432 vssd1 vssd1 vccd1 vccd1 _00108_ sky130_fd_sc_hd__mux2_1
Xinput8 DAT_I[15] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11853__A _05281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07181__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12999_ net1880 net298 net390 vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__mux2_1
XANTENNA__11064__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10068__A2 _01593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07469__B1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10188__B _04146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14669_ clknet_leaf_126_clk _01374_ net1205 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_119_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07210_ _02045_ vssd1 vssd1 vccd1 vccd1 _02046_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_15_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08190_ datapath.rf.registers\[17\]\[7\] net748 net724 datapath.rf.registers\[18\]\[7\]
+ _03025_ vssd1 vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__a221o_1
X_07141_ datapath.rf.registers\[17\]\[28\] net851 net830 datapath.rf.registers\[14\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__a22o_1
XFILLER_146_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10776__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07641__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07072_ _01899_ _01905_ _01907_ net785 datapath.rf.registers\[0\]\[30\] vssd1 vssd1
+ vccd1 vccd1 _01908_ sky130_fd_sc_hd__o32a_4
XFILLER_146_778 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06718__C_N _01500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08105__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07944__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11239__S net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07974_ datapath.rf.registers\[16\]\[11\] net740 net724 datapath.rf.registers\[18\]\[11\]
+ _02807_ vssd1 vssd1 vccd1 vccd1 _02810_ sky130_fd_sc_hd__a221o_1
X_09713_ net438 _04544_ _04548_ _03614_ vssd1 vssd1 vccd1 vccd1 _04549_ sky130_fd_sc_hd__o22a_1
X_06925_ datapath.rf.registers\[21\]\[31\] net815 net813 datapath.rf.registers\[23\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__a22o_1
XFILLER_56_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09644_ net346 _03967_ _04476_ _04479_ vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__a22o_1
X_06856_ net993 _01631_ datapath.ru.latched_instruction\[20\] vssd1 vssd1 vccd1 vccd1
+ _01692_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07172__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09575_ net381 _04061_ _04067_ _04410_ _03614_ vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__a311o_1
XFILLER_83_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_143_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06787_ net616 vssd1 vssd1 vccd1 vccd1 datapath.MUL_EN sky130_fd_sc_hd__inv_2
XANTENNA_fanout543_A net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08526_ datapath.rf.registers\[4\]\[0\] net960 net936 vssd1 vssd1 vccd1 vccd1 _03362_
+ sky130_fd_sc_hd__and3_1
XFILLER_24_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout710_A net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08457_ net610 _03266_ net581 vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout808_A net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout429_X net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07408_ datapath.rf.registers\[9\]\[22\] net981 net943 vssd1 vssd1 vccd1 vccd1 _02244_
+ sky130_fd_sc_hd__and3_1
XANTENNA__06683__B2 datapath.ru.latched_instruction\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__07880__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08388_ datapath.rf.registers\[26\]\[3\] net781 net693 datapath.rf.registers\[13\]\[3\]
+ _03223_ vssd1 vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__a221o_1
XFILLER_149_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07339_ datapath.rf.registers\[12\]\[24\] net755 net695 datapath.rf.registers\[8\]\[24\]
+ _02174_ vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__a221o_1
XFILLER_137_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10350_ _04852_ _05185_ vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__nand2b_1
XANTENNA__07632__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout798_X net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09009_ net459 _03843_ _03844_ vssd1 vssd1 vccd1 vccd1 _03845_ sky130_fd_sc_hd__and3_1
XFILLER_151_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10281_ _04475_ _04495_ vssd1 vssd1 vccd1 vccd1 _05117_ sky130_fd_sc_hd__and2_1
XANTENNA__10842__A net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12020_ _06059_ _06060_ _06061_ _06062_ vssd1 vssd1 vccd1 vccd1 _06063_ sky130_fd_sc_hd__or4_1
XFILLER_105_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11657__B _05874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout965_X net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11149__S net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout550 _03655_ vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09137__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout572 net573 vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10988__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13971_ clknet_leaf_105_clk _00749_ net1224 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_101_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout594 net595 vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__buf_2
X_12922_ net2117 net193 net482 vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__mux2_1
XFILLER_132_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12853_ net206 net1973 net486 vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__mux2_1
XFILLER_62_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ net2373 net1050 net315 net335 datapath.ru.latched_instruction\[10\] vssd1
+ vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__a32o_1
X_12784_ net231 net2172 net494 vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__mux2_1
XANTENNA__11798__A2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14523_ clknet_leaf_36_clk _01228_ net1135 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_11735_ net22 net1033 net1024 net1388 vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__o22a_1
X_14454_ clknet_leaf_141_clk _01159_ net1095 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_11666_ net2319 _05875_ _05882_ vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__a21o_1
XANTENNA__07871__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_14_0_clk_X clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13405_ clknet_leaf_147_clk _00215_ net1088 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10617_ net35 net36 _05382_ _05434_ vssd1 vssd1 vccd1 vccd1 _05437_ sky130_fd_sc_hd__and4b_2
XANTENNA__09612__A1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14385_ clknet_leaf_40_clk _01090_ net1140 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11597_ net1280 _01423_ screen.counter.ct\[9\] net1277 vssd1 vssd1 vccd1 vccd1 _05821_
+ sky130_fd_sc_hd__and4_1
Xwire951 _01711_ vssd1 vssd1 vccd1 vccd1 net951 sky130_fd_sc_hd__clkbuf_2
XFILLER_128_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07623__B1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13336_ clknet_leaf_6_clk _00146_ net1067 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_114_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10548_ keypad.debounce.debounce\[1\] keypad.debounce.debounce\[0\] keypad.debounce.debounce\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05375_ sky130_fd_sc_hd__and3_1
XFILLER_143_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13267_ clknet_leaf_41_clk _00077_ net1141 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10479_ screen.controlBus\[25\] screen.controlBus\[24\] screen.controlBus\[27\] screen.controlBus\[26\]
+ vssd1 vssd1 vccd1 vccd1 _05309_ sky130_fd_sc_hd__or4_1
X_12218_ _06221_ _06222_ vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_94_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13198_ clknet_leaf_3_clk _00008_ net1076 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11722__A2 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11059__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_102_Left_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12149_ _06154_ _06172_ vssd1 vssd1 vccd1 vccd1 _06180_ sky130_fd_sc_hd__and2_1
XFILLER_69_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09679__A1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06948__Y _01784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06710_ _01543_ _01544_ _01547_ _01548_ vssd1 vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__or4_1
XFILLER_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07690_ datapath.rf.registers\[3\]\[17\] net772 net716 datapath.rf.registers\[4\]\[17\]
+ _02525_ vssd1 vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__a221o_1
XANTENNA__08887__C1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07154__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06641_ mmio.memload_or_instruction\[12\] net1050 vssd1 vssd1 vccd1 vccd1 _01480_
+ sky130_fd_sc_hd__and2_1
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09360_ net561 net442 _04195_ net367 vssd1 vssd1 vccd1 vccd1 _04196_ sky130_fd_sc_hd__o211a_1
XFILLER_80_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06572_ datapath.ru.latched_instruction\[15\] vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__inv_2
XANTENNA__06964__X _01800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08311_ datapath.rf.registers\[23\]\[4\] net814 _03143_ _03146_ vssd1 vssd1 vccd1
+ vccd1 _03147_ sky130_fd_sc_hd__a211o_1
XANTENNA__09300__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_111_Left_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09291_ _03878_ _04126_ net376 vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__mux2_1
XANTENNA_13 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08242_ _03076_ _03077_ net611 vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__mux2_1
XANTENNA__07862__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07939__C net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08173_ datapath.rf.registers\[0\]\[7\] net867 net583 _03007_ vssd1 vssd1 vccd1 vccd1
+ _03009_ sky130_fd_sc_hd__a2bb2o_4
XANTENNA__09603__A1 _02857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07614__B1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07124_ datapath.rf.registers\[22\]\[28\] net954 net926 vssd1 vssd1 vccd1 vccd1 _01960_
+ sky130_fd_sc_hd__and3_1
XFILLER_146_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07055_ datapath.rf.registers\[26\]\[30\] net780 net760 datapath.rf.registers\[30\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__a22o_1
XFILLER_134_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput120 net120 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
XANTENNA__09367__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_120_Left_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout493_A _06551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11713__A2 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10921__B1 _05662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09119__A0 _02169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07393__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_145_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07957_ datapath.rf.registers\[2\]\[11\] net889 _02774_ _02780_ _02787_ vssd1 vssd1
+ vccd1 vccd1 _02793_ sky130_fd_sc_hd__a2111o_1
XFILLER_56_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout660_A net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout758_A _01802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06908_ _01629_ _01638_ vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__nor2_2
X_07888_ _02714_ _02723_ vssd1 vssd1 vccd1 vccd1 _02724_ sky130_fd_sc_hd__or2_1
XFILLER_16_607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13884__RESET_B net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09627_ net373 _04373_ net377 vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__o21ai_1
X_06839_ _01463_ net1002 net1018 net1026 datapath.ru.latched_instruction\[24\] vssd1
+ vssd1 vccd1 vccd1 _01675_ sky130_fd_sc_hd__a32oi_2
XFILLER_56_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout546_X net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout925_A net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09898__A _01585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09558_ net555 _04390_ _04392_ _04339_ net631 vssd1 vssd1 vccd1 vccd1 _04394_ sky130_fd_sc_hd__a32o_1
X_08509_ datapath.rf.registers\[6\]\[1\] net682 _03342_ _03343_ _03344_ vssd1 vssd1
+ vccd1 vccd1 _03345_ sky130_fd_sc_hd__a2111o_1
XFILLER_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09489_ net560 net464 net441 vssd1 vssd1 vccd1 vccd1 _04325_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout713_X net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07302__C1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11432__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11520_ _05333_ _05356_ _05737_ _05744_ vssd1 vssd1 vccd1 vccd1 _05745_ sky130_fd_sc_hd__and4_1
XFILLER_12_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07853__B1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11451_ net1868 net285 net408 vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__mux2_1
XFILLER_109_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10402_ datapath.PC\[0\] _05237_ _05212_ vssd1 vssd1 vccd1 vccd1 _05238_ sky130_fd_sc_hd__mux2_1
X_14170_ clknet_leaf_55_clk _00925_ net1179 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11382_ net1889 net294 net411 vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__mux2_1
X_13121_ net192 net2621 net470 vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__mux2_1
X_10333_ datapath.PC\[14\] _03739_ vssd1 vssd1 vccd1 vccd1 _05169_ sky130_fd_sc_hd__nand2_1
XFILLER_3_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10572__A _02612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08313__Y _03149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13052_ net203 net1727 net475 vssd1 vssd1 vccd1 vccd1 _01296_ sky130_fd_sc_hd__mux2_1
X_10264_ _04582_ _05099_ _05098_ vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_76_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08042__A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12003_ screen.register.currentYbus\[17\] _05773_ net997 screen.register.currentXbus\[17\]
+ _06046_ vssd1 vssd1 vccd1 vccd1 _06047_ sky130_fd_sc_hd__a221o_1
XANTENNA__08030__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10195_ datapath.PC\[17\] net1256 _05027_ _05030_ vssd1 vssd1 vccd1 vccd1 _05031_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08977__A net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07384__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout380 net381 vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__clkbuf_2
XFILLER_93_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout391 net393 vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__clkbuf_8
X_13954_ clknet_leaf_99_clk _00732_ net1229 vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10125__D1 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07136__A2 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12905_ net1792 net277 net484 vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__mux2_1
XANTENNA__10140__A1 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13885_ clknet_leaf_74_clk _00689_ net1247 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[29\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_19_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12836_ net291 net2008 net486 vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__mux2_1
XFILLER_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12767_ net302 net1902 net497 vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__mux2_1
XANTENNA__10747__A _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06944__B net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14506_ clknet_leaf_59_clk _01211_ net1169 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11718_ net4 net1034 net1024 net2116 vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__o22a_1
X_12698_ _06527_ _06528_ vssd1 vssd1 vccd1 vccd1 _06529_ sky130_fd_sc_hd__xnor2_1
XFILLER_147_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07121__A _01935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14437_ clknet_leaf_116_clk _01142_ net1188 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput11 DAT_I[18] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
X_11649_ screen.screenLogic.currentWrx _05872_ _05870_ vssd1 vssd1 vccd1 vccd1 _00548_
+ sky130_fd_sc_hd__mux2_1
Xinput22 DAT_I[28] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
XFILLER_128_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput33 DAT_I[9] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_96_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14368_ clknet_leaf_137_clk _01073_ net1097 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold806 datapath.rf.registers\[11\]\[21\] vssd1 vssd1 vccd1 vccd1 net2154 sky130_fd_sc_hd__dlygate4sd3_1
Xhold817 datapath.rf.registers\[29\]\[23\] vssd1 vssd1 vccd1 vccd1 net2165 sky130_fd_sc_hd__dlygate4sd3_1
X_13319_ clknet_leaf_142_clk _00129_ net1087 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold828 datapath.rf.registers\[26\]\[7\] vssd1 vssd1 vccd1 vccd1 net2176 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07072__B2 datapath.rf.registers\[0\]\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold839 datapath.rf.registers\[1\]\[10\] vssd1 vssd1 vccd1 vccd1 net2187 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14299_ clknet_leaf_91_clk _01004_ net1241 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[19\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_143_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09048__A _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12353__C1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08860_ net342 _03695_ vssd1 vssd1 vccd1 vccd1 _03696_ sky130_fd_sc_hd__or2_1
XANTENNA__08021__B1 _02855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12901__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07811_ datapath.rf.registers\[22\]\[14\] net822 net817 datapath.rf.registers\[7\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02647_ sky130_fd_sc_hd__a22o_1
X_08791_ _03617_ net375 vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_127_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07742_ datapath.rf.registers\[14\]\[16\] net774 net718 datapath.rf.registers\[20\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__a22o_1
XANTENNA__07127__A2 _01713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07673_ datapath.rf.registers\[1\]\[17\] net847 net838 datapath.rf.registers\[26\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02509_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_140_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09412_ _04245_ _04246_ net455 vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__a21oi_1
X_06624_ mmio.memload_or_instruction\[24\] net1049 vssd1 vssd1 vccd1 vccd1 _01463_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_140_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10419__C1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09343_ _03519_ _03521_ vssd1 vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__nand2_2
XANTENNA__08088__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11252__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07835__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09274_ _03667_ _04108_ _04109_ _04098_ vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07669__C net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08225_ datapath.rf.registers\[22\]\[6\] net734 net668 datapath.rf.registers\[21\]\[6\]
+ _03059_ vssd1 vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__a221o_1
XFILLER_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout127_X net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout506_A net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1248_A net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08156_ datapath.rf.registers\[17\]\[7\] net851 net847 datapath.rf.registers\[1\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__a22o_1
XANTENNA__10198__A1 _03978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06870__A _01579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07107_ datapath.rf.registers\[29\]\[29\] net676 net661 datapath.rf.registers\[5\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__a22o_1
XANTENNA__08260__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08087_ datapath.rf.registers\[16\]\[9\] net740 _02920_ _02922_ net788 vssd1 vssd1
+ vccd1 vccd1 _02923_ sky130_fd_sc_hd__a2111oi_1
X_07038_ datapath.rf.registers\[1\]\[30\] net847 _01871_ _01872_ _01873_ vssd1 vssd1
+ vccd1 vccd1 _01874_ sky130_fd_sc_hd__a2111o_1
XFILLER_122_718 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14012__RESET_B net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout496_X net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout875_A _01723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12811__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09392__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09760__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout663_X net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08989_ _03470_ _03487_ _03824_ vssd1 vssd1 vccd1 vccd1 _03825_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11427__S net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07118__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout830_X net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10951_ _01644_ _01663_ vssd1 vssd1 vccd1 vccd1 _05689_ sky130_fd_sc_hd__nand2_1
XANTENNA__10122__A1 _04057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout928_X net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11951__A _01854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13670_ clknet_leaf_23_clk _00480_ net1154 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10882_ datapath.PC\[21\] _05617_ net1265 vssd1 vssd1 vccd1 vccd1 _05630_ sky130_fd_sc_hd__a21oi_1
X_12621_ _06457_ _06463_ _06462_ _06461_ vssd1 vssd1 vccd1 vccd1 _06465_ sky130_fd_sc_hd__o211ai_2
XANTENNA__08079__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11162__S net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_125_Right_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07826__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12552_ _06405_ _06406_ vssd1 vssd1 vccd1 vccd1 _06407_ sky130_fd_sc_hd__nor2_1
XFILLER_8_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11503_ net196 net1765 net512 vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__mux2_1
XFILLER_7_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12483_ net294 datapath.rf.registers\[31\]\[5\] net506 vssd1 vssd1 vccd1 vccd1 _00883_
+ sky130_fd_sc_hd__mux2_1
X_14222_ clknet_leaf_41_clk _00943_ net1153 vssd1 vssd1 vccd1 vccd1 columns.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_22_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11434_ net201 net2466 net515 vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13089__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14153_ clknet_leaf_78_clk MemWrite net1248 vssd1 vssd1 vccd1 vccd1 datapath.ru.n_memwrite
+ sky130_fd_sc_hd__dfrtp_4
X_11365_ net212 net1651 net519 vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__mux2_1
XANTENNA__08251__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_100_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_100_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_98_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13104_ net274 net2557 net471 vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__mux2_1
X_10316_ net1044 _05151_ _05150_ net639 vssd1 vssd1 vccd1 vccd1 _05152_ sky130_fd_sc_hd__a211o_1
X_14084_ clknet_leaf_108_clk _00850_ net1218 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11296_ net213 net1754 net522 vssd1 vssd1 vccd1 vccd1 _00344_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08203__C net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13035_ net290 net2575 net475 vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__mux2_1
XFILLER_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10247_ net892 _05078_ _05080_ _05082_ vssd1 vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__o22a_1
XFILLER_67_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1120 net1121 vssd1 vssd1 vccd1 vccd1 net1120 sky130_fd_sc_hd__buf_2
XANTENNA__12350__A2 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1131 net1139 vssd1 vssd1 vccd1 vccd1 net1131 sky130_fd_sc_hd__clkbuf_4
Xfanout1142 net1143 vssd1 vssd1 vccd1 vccd1 net1142 sky130_fd_sc_hd__clkbuf_2
Xfanout1153 net1186 vssd1 vssd1 vccd1 vccd1 net1153 sky130_fd_sc_hd__clkbuf_4
X_10178_ _03950_ _04605_ vssd1 vssd1 vccd1 vccd1 _05014_ sky130_fd_sc_hd__or2_1
XANTENNA__11337__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1164 net1166 vssd1 vssd1 vccd1 vccd1 net1164 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06939__B net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1175 net1178 vssd1 vssd1 vccd1 vccd1 net1175 sky130_fd_sc_hd__clkbuf_4
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1186 _00004_ vssd1 vssd1 vccd1 vccd1 net1186 sky130_fd_sc_hd__clkbuf_4
Xfanout1197 net1204 vssd1 vssd1 vccd1 vccd1 net1197 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07109__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13937_ clknet_leaf_108_clk _00715_ net1218 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11861__A _03357_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13868_ clknet_leaf_75_clk _00672_ net1246 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[12\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_35_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06955__A net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12819_ net1772 net212 net490 vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__mux2_1
X_13799_ clknet_leaf_52_clk _00608_ net1183 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07817__B1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08010_ net874 _02843_ _02844_ _02845_ vssd1 vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_100_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold603 datapath.rf.registers\[26\]\[4\] vssd1 vssd1 vccd1 vccd1 net1951 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08242__A0 _03076_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold614 datapath.rf.registers\[8\]\[4\] vssd1 vssd1 vccd1 vccd1 net1962 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold625 datapath.rf.registers\[30\]\[23\] vssd1 vssd1 vccd1 vccd1 net1973 sky130_fd_sc_hd__dlygate4sd3_1
Xhold636 datapath.rf.registers\[27\]\[5\] vssd1 vssd1 vccd1 vccd1 net1984 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08793__A1 _03358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold647 datapath.rf.registers\[3\]\[7\] vssd1 vssd1 vccd1 vccd1 net1995 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07596__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold658 datapath.rf.registers\[19\]\[20\] vssd1 vssd1 vccd1 vccd1 net2006 sky130_fd_sc_hd__dlygate4sd3_1
X_09961_ _04794_ _04795_ _04765_ vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__a21o_1
Xhold669 datapath.rf.registers\[30\]\[20\] vssd1 vssd1 vccd1 vccd1 net2017 sky130_fd_sc_hd__dlygate4sd3_1
X_08912_ net1264 datapath.PC\[25\] _03747_ vssd1 vssd1 vccd1 vccd1 _03748_ sky130_fd_sc_hd__or3b_2
X_09892_ _01585_ net900 net979 vssd1 vssd1 vccd1 vccd1 _04728_ sky130_fd_sc_hd__and3_1
XFILLER_134_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07348__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09742__B1 _04575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08843_ _03419_ net992 _03671_ vssd1 vssd1 vccd1 vccd1 _03679_ sky130_fd_sc_hd__mux2_1
XANTENNA__07952__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1303 datapath.PC\[5\] vssd1 vssd1 vccd1 vccd1 net2651 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11247__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08774_ _01605_ net651 net646 net631 vssd1 vssd1 vccd1 vccd1 _03610_ sky130_fd_sc_hd__a31o_1
X_07725_ datapath.rf.registers\[16\]\[16\] net860 net810 datapath.rf.registers\[13\]\[16\]
+ _02560_ vssd1 vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__a221o_1
XFILLER_72_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_2_0_clk_X clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1198_A net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07656_ datapath.rf.registers\[20\]\[17\] net959 net925 vssd1 vssd1 vccd1 vccd1 _02492_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07520__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06607_ net1288 net1283 mmio.memload_or_instruction\[13\] vssd1 vssd1 vccd1 vccd1
+ _01446_ sky130_fd_sc_hd__nor3b_2
XFILLER_43_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07587_ datapath.rf.registers\[8\]\[19\] net696 net677 datapath.rf.registers\[29\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__a22o_1
XFILLER_43_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09326_ _04158_ _04160_ net461 vssd1 vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__mux2_1
XANTENNA__07808__B1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09257_ net364 _04090_ _04091_ net374 vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout411_X net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08481__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12806__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1153_X net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06871__Y _01707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout509_X net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08208_ net872 _03041_ _03042_ _03043_ vssd1 vssd1 vccd1 vccd1 _03044_ sky130_fd_sc_hd__or4_1
XFILLER_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09188_ _02333_ _03455_ vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__and2b_1
XANTENNA__08144__X _02980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08233__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08139_ datapath.rf.registers\[12\]\[8\] net756 net673 datapath.rf.registers\[7\]\[8\]
+ _02974_ vssd1 vssd1 vccd1 vccd1 _02975_ sky130_fd_sc_hd__a221o_1
XFILLER_134_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07587__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11150_ net276 net2250 net532 vssd1 vssd1 vccd1 vccd1 _00203_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout780_X net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout878_X net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10101_ _03749_ _04936_ net1042 vssd1 vssd1 vccd1 vccd1 _04937_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_73_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12868__A0 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11081_ net278 net2122 net537 vssd1 vssd1 vccd1 vccd1 _00138_ sky130_fd_sc_hd__mux2_1
XFILLER_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07339__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10032_ _04864_ _04865_ _04867_ vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__or3b_2
XANTENNA__11665__B _05874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11157__S net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10894__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input17_A DAT_I[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10996__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_149_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_149_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11983_ screen.register.currentYbus\[8\] _05776_ net997 screen.register.currentXbus\[16\]
+ _06027_ vssd1 vssd1 vccd1 vccd1 _06028_ sky130_fd_sc_hd__a221o_1
XFILLER_84_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13722_ clknet_leaf_2_clk _00532_ net1065 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_90_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10934_ net898 _04645_ _05674_ net600 vssd1 vssd1 vccd1 vccd1 _05675_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_104_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13653_ clknet_leaf_129_clk _00463_ net1117 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_896 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10865_ _01469_ net652 _05614_ _05615_ vssd1 vssd1 vccd1 vccd1 _05616_ sky130_fd_sc_hd__o22a_2
XTAP_TAPCELL_ROW_27_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12604_ net499 _06449_ _06450_ net503 net2161 vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__a32o_1
X_13584_ clknet_leaf_24_clk _00394_ net1158 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10796_ datapath.mulitply_result\[9\] net598 net620 vssd1 vssd1 vccd1 vccd1 _05557_
+ sky130_fd_sc_hd__a21oi_1
X_12535_ _06390_ _06391_ _06392_ vssd1 vssd1 vccd1 vccd1 _06393_ sky130_fd_sc_hd__or3_1
XANTENNA__08472__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06781__Y _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12466_ net164 _05980_ net126 screen.register.currentXbus\[22\] vssd1 vssd1 vccd1
+ vccd1 _00868_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14205_ clknet_leaf_55_clk datapath.multiplication_module.multiplicand_i_n\[16\]
+ net1180 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11417_ net284 net2582 net516 vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__mux2_1
XANTENNA__08224__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12397_ _05954_ net159 vssd1 vssd1 vccd1 vccd1 _06346_ sky130_fd_sc_hd__nor2_1
XFILLER_126_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14136_ clknet_leaf_126_clk _00893_ net1206 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11348_ net295 net1979 net518 vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__mux2_1
XANTENNA__07983__C1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14067_ clknet_leaf_111_clk _00834_ net1198 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_3_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11279_ net296 net2492 net522 vssd1 vssd1 vccd1 vccd1 _00327_ sky130_fd_sc_hd__mux2_1
X_13018_ net1540 net203 net391 vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__mux2_1
XANTENNA__11067__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08884__B _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07510_ datapath.rf.registers\[4\]\[20\] net957 net932 vssd1 vssd1 vccd1 vccd1 _02346_
+ sky130_fd_sc_hd__and3_1
XFILLER_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08490_ datapath.rf.registers\[1\]\[1\] net914 _01800_ vssd1 vssd1 vccd1 vccd1 _03326_
+ sky130_fd_sc_hd__and3_1
X_07441_ datapath.rf.registers\[23\]\[22\] net698 net671 datapath.rf.registers\[7\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__a22o_1
X_07372_ datapath.rf.registers\[9\]\[23\] net885 net799 datapath.rf.registers\[15\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_40_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09111_ _03918_ _03946_ net632 vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__a21o_2
XFILLER_148_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire581_X net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09042_ _03877_ vssd1 vssd1 vccd1 vccd1 _03878_ sky130_fd_sc_hd__inv_2
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07947__C net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold400 datapath.rf.registers\[4\]\[17\] vssd1 vssd1 vccd1 vccd1 net1748 sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 datapath.rf.registers\[22\]\[24\] vssd1 vssd1 vccd1 vccd1 net1759 sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 datapath.rf.registers\[4\]\[6\] vssd1 vssd1 vccd1 vccd1 net1770 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout204_A _05641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07569__A2 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold433 datapath.rf.registers\[8\]\[8\] vssd1 vssd1 vccd1 vccd1 net1781 sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 datapath.rf.registers\[16\]\[9\] vssd1 vssd1 vccd1 vccd1 net1792 sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 datapath.rf.registers\[12\]\[23\] vssd1 vssd1 vccd1 vccd1 net1803 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold466 datapath.rf.registers\[7\]\[7\] vssd1 vssd1 vccd1 vccd1 net1814 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold477 datapath.rf.registers\[31\]\[27\] vssd1 vssd1 vccd1 vccd1 net1825 sky130_fd_sc_hd__dlygate4sd3_1
Xhold488 datapath.rf.registers\[11\]\[1\] vssd1 vssd1 vccd1 vccd1 net1836 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09944_ _03322_ _03323_ datapath.PC\[1\] vssd1 vssd1 vccd1 vccd1 _04780_ sky130_fd_sc_hd__o21a_1
Xfanout902 net903 vssd1 vssd1 vccd1 vccd1 net902 sky130_fd_sc_hd__clkbuf_4
Xfanout913 _01789_ vssd1 vssd1 vccd1 vccd1 net913 sky130_fd_sc_hd__clkbuf_2
Xhold499 datapath.rf.registers\[25\]\[2\] vssd1 vssd1 vccd1 vccd1 net1847 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout924 net926 vssd1 vssd1 vccd1 vccd1 net924 sky130_fd_sc_hd__buf_2
XANTENNA__12314__A2 _06253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07308__X _02144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout935 net936 vssd1 vssd1 vccd1 vccd1 net935 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout946 net948 vssd1 vssd1 vccd1 vccd1 net946 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input9_A DAT_I[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09875_ net633 _04710_ vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__and2_2
Xfanout957 net960 vssd1 vssd1 vccd1 vccd1 net957 sky130_fd_sc_hd__buf_2
XANTENNA__10325__A1 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1100 datapath.rf.registers\[31\]\[21\] vssd1 vssd1 vccd1 vccd1 net2448 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout968 net969 vssd1 vssd1 vccd1 vccd1 net968 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout573_A _05367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1111 datapath.rf.registers\[16\]\[22\] vssd1 vssd1 vccd1 vccd1 net2459 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout979 net980 vssd1 vssd1 vccd1 vccd1 net979 sky130_fd_sc_hd__buf_4
Xhold1122 datapath.rf.registers\[31\]\[22\] vssd1 vssd1 vccd1 vccd1 net2470 sky130_fd_sc_hd__dlygate4sd3_1
X_08826_ net967 _03171_ _03643_ vssd1 vssd1 vccd1 vccd1 _03662_ sky130_fd_sc_hd__mux2_1
Xhold1133 screen.register.currentYbus\[13\] vssd1 vssd1 vccd1 vccd1 net2481 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1144 datapath.rf.registers\[25\]\[5\] vssd1 vssd1 vccd1 vccd1 net2492 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1155 datapath.rf.registers\[26\]\[15\] vssd1 vssd1 vccd1 vccd1 net2503 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07741__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1166 screen.register.currentYbus\[2\] vssd1 vssd1 vccd1 vccd1 net2514 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1177 datapath.rf.registers\[30\]\[12\] vssd1 vssd1 vccd1 vccd1 net2525 sky130_fd_sc_hd__dlygate4sd3_1
X_08757_ _03492_ _03494_ _03591_ _03490_ vssd1 vssd1 vccd1 vccd1 _03593_ sky130_fd_sc_hd__a31o_1
Xhold1188 datapath.rf.registers\[29\]\[29\] vssd1 vssd1 vccd1 vccd1 net2536 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout740_A net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1199 mmio.wishbone.curr_state\[1\] vssd1 vssd1 vccd1 vccd1 net2547 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06866__Y _01702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10089__B1 _01702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout838_A _01743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07708_ _02522_ _02543_ vssd1 vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__and2_1
XANTENNA__11825__A1 _01477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08688_ _03522_ _03523_ vssd1 vssd1 vccd1 vccd1 _03524_ sky130_fd_sc_hd__nor2_2
XFILLER_81_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07639_ datapath.rf.registers\[30\]\[18\] net758 net734 datapath.rf.registers\[22\]\[18\]
+ _02474_ vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__a221o_1
XFILLER_41_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout626_X net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10650_ _05435_ _05445_ _05468_ _05469_ _05467_ vssd1 vssd1 vccd1 vccd1 _05470_ sky130_fd_sc_hd__o311a_1
XFILLER_10_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09309_ net607 _04120_ _04144_ net556 vssd1 vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__o211a_1
XANTENNA__09797__A3 _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10581_ _01934_ _05400_ _05401_ _05403_ vssd1 vssd1 vccd1 vccd1 _05404_ sky130_fd_sc_hd__or4_1
XANTENNA__11440__S net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12320_ net640 _04869_ vssd1 vssd1 vccd1 vccd1 _06295_ sky130_fd_sc_hd__nor2_1
XFILLER_6_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout995_X net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08206__B1 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12251_ net1379 _06242_ net602 vssd1 vssd1 vccd1 vccd1 _06243_ sky130_fd_sc_hd__o21ai_1
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11202_ net177 net1906 net424 vssd1 vssd1 vccd1 vccd1 _00254_ sky130_fd_sc_hd__mux2_1
XFILLER_135_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12182_ _06159_ net601 vssd1 vssd1 vccd1 vccd1 _06200_ sky130_fd_sc_hd__and2_1
XFILLER_108_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11133_ net193 net2336 net426 vssd1 vssd1 vccd1 vccd1 _00188_ sky130_fd_sc_hd__mux2_1
XANTENNA__10580__A _02418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07980__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11064_ net192 net2295 net430 vssd1 vssd1 vccd1 vccd1 _00124_ sky130_fd_sc_hd__mux2_1
XFILLER_135_83 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10316__A1 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10015_ _04846_ _04847_ _04850_ vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__or3_2
XANTENNA__07193__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07732__A2 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14754_ net1291 vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__clkbuf_1
X_11966_ net1010 _05794_ _05798_ _06006_ _06011_ vssd1 vssd1 vccd1 vccd1 _06012_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_86_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10917_ datapath.PC\[27\] _05654_ vssd1 vssd1 vccd1 vccd1 _05660_ sky130_fd_sc_hd__xnor2_1
X_13705_ clknet_leaf_20_clk _00515_ net1165 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07496__A1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14685_ clknet_leaf_146_clk _01390_ net1088 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11897_ _02725_ net657 vssd1 vssd1 vccd1 vccd1 _05962_ sky130_fd_sc_hd__nand2_1
XFILLER_32_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13636_ clknet_leaf_21_clk _00446_ net1163 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10848_ datapath.PC\[17\] _05593_ vssd1 vssd1 vccd1 vccd1 _05601_ sky130_fd_sc_hd__nor2_1
XFILLER_13_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13567_ clknet_leaf_14_clk _00377_ net1078 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08445__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10779_ net1268 datapath.PC\[7\] _05530_ vssd1 vssd1 vccd1 vccd1 _05542_ sky130_fd_sc_hd__and3_1
XANTENNA__06952__B net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11350__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07799__A2 _02633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12518_ datapath.mulitply_result\[0\] datapath.multiplication_module.multiplicand_i\[0\]
+ _06376_ vssd1 vssd1 vccd1 vccd1 _06379_ sky130_fd_sc_hd__a21o_1
X_13498_ clknet_leaf_3_clk _00308_ net1076 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_117_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12449_ net165 _05946_ net127 screen.register.currentXbus\[5\] vssd1 vssd1 vccd1
+ vccd1 _00851_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14119_ clknet_leaf_75_clk net1510 net1246 vssd1 vssd1 vccd1 vccd1 datapath.ru.n_memwrite2
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13750__RESET_B net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07990_ _02804_ _02825_ vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__or2_1
Xfanout209 _05700_ vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__clkbuf_2
XFILLER_87_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07971__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06941_ datapath.rf.registers\[31\]\[31\] net793 net790 datapath.rf.registers\[18\]\[31\]
+ _01774_ vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__a221o_1
XFILLER_113_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09660_ _04475_ _04495_ vssd1 vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__nor2_1
X_06872_ _01656_ net962 vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__nor2_1
XANTENNA__07184__B1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07723__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08611_ _02636_ _03446_ _02637_ vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__a21oi_1
XFILLER_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09591_ _03637_ _04403_ _04426_ _04400_ vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__a31o_1
XANTENNA__06931__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08542_ datapath.rf.registers\[2\]\[0\] net889 net795 datapath.rf.registers\[31\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__a22o_1
X_08473_ net875 _03304_ _03306_ _03308_ vssd1 vssd1 vccd1 vccd1 _03309_ sky130_fd_sc_hd__or4_1
XFILLER_62_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout154_A net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07424_ datapath.rf.registers\[6\]\[22\] net824 _02243_ _02245_ _02247_ vssd1 vssd1
+ vccd1 vccd1 _02260_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_137_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07355_ _02170_ _02190_ vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__nor2_1
XANTENNA__11260__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout419_A _05722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07286_ datapath.rf.registers\[29\]\[25\] net797 _02097_ _02107_ _02108_ vssd1 vssd1
+ vccd1 vccd1 _02122_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_150_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09025_ net904 _03828_ _03859_ net318 vssd1 vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__o22a_1
XFILLER_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1230_A net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold230 datapath.rf.registers\[4\]\[0\] vssd1 vssd1 vccd1 vccd1 net1578 sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 datapath.rf.registers\[17\]\[13\] vssd1 vssd1 vccd1 vccd1 net1589 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09892__C net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09400__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold252 datapath.multiplication_module.multiplicand_i\[8\] vssd1 vssd1 vccd1 vccd1
+ net1600 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout788_A net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold263 datapath.rf.registers\[10\]\[7\] vssd1 vssd1 vccd1 vccd1 net1611 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold274 datapath.rf.registers\[4\]\[15\] vssd1 vssd1 vccd1 vccd1 net1622 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold285 datapath.rf.registers\[12\]\[20\] vssd1 vssd1 vccd1 vccd1 net1633 sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 datapath.rf.registers\[9\]\[10\] vssd1 vssd1 vccd1 vccd1 net1644 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout710 net713 vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__buf_4
Xfanout721 _01814_ vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__clkbuf_4
XFILLER_49_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout732 _01811_ vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__buf_4
XANTENNA__07962__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09927_ net1267 _02935_ vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__or2_1
Xfanout743 net745 vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__clkbuf_4
Xfanout754 net757 vssd1 vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__buf_4
XANTENNA_fanout576_X net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout955_A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout765 _01801_ vssd1 vssd1 vccd1 vccd1 net765 sky130_fd_sc_hd__clkbuf_4
Xfanout776 _01796_ vssd1 vssd1 vccd1 vccd1 net776 sky130_fd_sc_hd__buf_4
Xfanout787 net789 vssd1 vssd1 vccd1 vccd1 net787 sky130_fd_sc_hd__buf_4
X_09858_ _03466_ _04669_ _04693_ vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06877__X _01713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07175__B1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout798 _01773_ vssd1 vssd1 vccd1 vccd1 net798 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_29_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08809_ _01647_ _03644_ vssd1 vssd1 vccd1 vccd1 _03645_ sky130_fd_sc_hd__nand2_1
X_09789_ _03916_ _04607_ _04624_ vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__or3b_2
XANTENNA_fanout743_X net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06596__Y _01436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11435__S net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11820_ datapath.ru.latched_instruction\[26\] net336 net316 _01503_ vssd1 vssd1 vccd1
+ vccd1 _00686_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_68_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ net1495 net144 net139 _02824_ vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__a22o_1
XFILLER_42_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_80_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_42_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10702_ net1468 _03028_ net570 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i_n\[7\]
+ sky130_fd_sc_hd__mux2_1
X_14470_ clknet_leaf_17_clk _01175_ net1107 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11682_ _05095_ net152 net151 net1455 vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__a22o_1
X_13421_ clknet_leaf_133_clk _00231_ net1112 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_81_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10633_ _05432_ _05433_ vssd1 vssd1 vccd1 vccd1 _05453_ sky130_fd_sc_hd__nor2_1
XANTENNA__08427__B1 _03261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10575__A _03205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11170__S net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06772__B _01607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13352_ clknet_leaf_65_clk _00162_ net1238 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10564_ _05385_ _05387_ vssd1 vssd1 vccd1 vccd1 _05388_ sky130_fd_sc_hd__or2_1
XFILLER_128_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08045__A _02856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12303_ _05579_ _06254_ _06282_ net190 vssd1 vssd1 vccd1 vccd1 _06283_ sky130_fd_sc_hd__o22a_1
XANTENNA__11982__B1 _05786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13283_ clknet_leaf_120_clk _00093_ net1192 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10495_ _05324_ vssd1 vssd1 vccd1 vccd1 _05325_ sky130_fd_sc_hd__inv_2
XFILLER_6_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12234_ _06168_ _06231_ _06232_ vssd1 vssd1 vccd1 vccd1 _00773_ sky130_fd_sc_hd__nor3_1
XANTENNA__09428__X _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Left_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13097__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12165_ screen.counter.ct\[11\] _06186_ net1274 vssd1 vssd1 vccd1 vccd1 _06190_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_112_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11116_ net275 net1806 net428 vssd1 vssd1 vccd1 vccd1 _00171_ sky130_fd_sc_hd__mux2_1
X_12096_ screen.register.currentYbus\[15\] _05776_ net997 screen.register.currentXbus\[23\]
+ _06133_ vssd1 vssd1 vccd1 vccd1 _06134_ sky130_fd_sc_hd__a221o_1
XFILLER_150_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_10_0_clk_X clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11047_ net275 net2054 net432 vssd1 vssd1 vccd1 vccd1 _00107_ sky130_fd_sc_hd__mux2_1
Xinput9 DAT_I[16] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11345__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06947__B net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_24_Left_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12998_ net1567 net303 net393 vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__mux2_1
XFILLER_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10068__A3 _01784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11949_ net134 _05996_ _05995_ vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_71_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08130__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09610__Y _04446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14668_ clknet_leaf_14_clk _01373_ net1102 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06963__A net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13619_ clknet_leaf_34_clk _00429_ net1128 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_14599_ clknet_leaf_137_clk _01304_ net1089 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11080__S net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07140_ _01973_ _01974_ _01975_ vssd1 vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__or3_1
XFILLER_9_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09091__B1 _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13931__RESET_B net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07071_ _01890_ _01891_ _01892_ _01906_ vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_33_Left_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12904__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08402__B net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07973_ datapath.rf.registers\[2\]\[11\] net744 net681 datapath.rf.registers\[6\]\[11\]
+ _02808_ vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__a221o_1
XFILLER_141_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09712_ net379 _04545_ _04546_ _04547_ vssd1 vssd1 vccd1 vccd1 _04548_ sky130_fd_sc_hd__a22o_1
X_06924_ net940 net921 vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__and2_2
XFILLER_142_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07157__B1 _01832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09643_ net359 _04477_ _04478_ net345 vssd1 vssd1 vccd1 vccd1 _04479_ sky130_fd_sc_hd__a31oi_1
X_06855_ datapath.ru.latched_instruction\[6\] _01580_ _01586_ datapath.ru.latched_instruction\[3\]
+ _01690_ vssd1 vssd1 vccd1 vccd1 _01691_ sky130_fd_sc_hd__a221o_1
XFILLER_27_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10700__A1 _03123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout271_A _05564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11255__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09574_ net377 _04407_ _04409_ net330 vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__o211a_1
X_06786_ _01605_ net651 net643 vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_143_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14037__RESET_B net1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08525_ net559 _03358_ vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__nor2_1
XFILLER_70_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10947__X _05686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1180_A net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout536_A net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout157_X net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_62_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_60_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08121__A2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08456_ _03266_ net581 vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__nor2_4
XANTENNA__06873__A net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07407_ datapath.rf.registers\[20\]\[22\] net957 net921 vssd1 vssd1 vccd1 vccd1 _02243_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_34_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08387_ datapath.rf.registers\[12\]\[3\] net756 net704 datapath.rf.registers\[9\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__a22o_1
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout703_A net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout324_X net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07338_ datapath.rf.registers\[23\]\[24\] net699 net672 datapath.rf.registers\[7\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__a22o_1
XANTENNA__09082__B1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_75_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12814__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07269_ datapath.rf.registers\[23\]\[25\] net941 net926 vssd1 vssd1 vccd1 vccd1 _02105_
+ sky130_fd_sc_hd__and3_1
X_09008_ net551 net547 _02025_ vssd1 vssd1 vccd1 vccd1 _03844_ sky130_fd_sc_hd__a21o_1
XANTENNA__09248__X _04084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10280_ net1267 net1254 _05112_ _05115_ vssd1 vssd1 vccd1 vccd1 _05116_ sky130_fd_sc_hd__o22a_1
XFILLER_3_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout693_X net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08188__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07396__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07935__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_133_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout860_X net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout958_X net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout540 net541 vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__clkbuf_8
XFILLER_116_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout551 _03654_ vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__buf_2
X_13970_ clknet_leaf_105_clk _00748_ net1224 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout573 _05367_ vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_13_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07148__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout595 net596 vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__buf_2
XFILLER_101_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12921_ net1854 net196 net484 vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__mux2_1
XFILLER_100_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11165__S net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08360__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_148_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12852_ net210 net2485 net486 vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _01536_ net1016 net316 net336 datapath.ru.latched_instruction\[9\] vssd1
+ vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__a32o_1
X_12783_ net236 net1598 net496 vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_28_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_53_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_15_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08112__A2 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11734_ net21 net1034 net1024 net1786 vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__o22a_1
XFILLER_14_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14522_ clknet_leaf_14_clk _01227_ net1102 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_25_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07320__B1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06783__A _01614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11665_ keypad.apps.app_c\[1\] _05874_ vssd1 vssd1 vccd1 vccd1 _05882_ sky130_fd_sc_hd__and2_1
X_14453_ clknet_leaf_130_clk _01158_ net1116 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_4_6_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_6_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_30_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10616_ net35 net36 _05379_ _05382_ vssd1 vssd1 vccd1 vccd1 _05436_ sky130_fd_sc_hd__and4b_1
X_13404_ clknet_leaf_10_clk _00214_ net1081 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_14384_ clknet_leaf_25_clk _01089_ net1158 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11596_ _05758_ _05775_ vssd1 vssd1 vccd1 vccd1 _05820_ sky130_fd_sc_hd__and2_1
X_13335_ clknet_leaf_130_clk _00145_ net1111 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_127_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10547_ keypad.debounce.debounce\[5\] keypad.debounce.debounce\[4\] keypad.debounce.debounce\[7\]
+ keypad.debounce.debounce\[6\] vssd1 vssd1 vccd1 vccd1 _05374_ sky130_fd_sc_hd__and4_1
XANTENNA__08281__D1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13266_ clknet_leaf_33_clk _00076_ net1125 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10478_ screen.controlBus\[29\] screen.controlBus\[28\] screen.controlBus\[31\] screen.controlBus\[30\]
+ vssd1 vssd1 vccd1 vccd1 _05308_ sky130_fd_sc_hd__or4_1
X_12217_ net2593 _06219_ net602 vssd1 vssd1 vccd1 vccd1 _06222_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_94_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13197_ clknet_leaf_125_clk _00007_ net1207 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07926__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12148_ _06152_ net603 vssd1 vssd1 vccd1 vccd1 _06179_ sky130_fd_sc_hd__or2_1
XFILLER_150_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11864__A _03292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12079_ _06043_ _06116_ _06118_ _06105_ vssd1 vssd1 vccd1 vccd1 _06119_ sky130_fd_sc_hd__or4b_1
XFILLER_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07139__B1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_139_Right_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11075__S net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06640_ net1288 net1284 mmio.memload_or_instruction\[27\] vssd1 vssd1 vccd1 vccd1
+ _01479_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_125_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11870__Y _05944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06571_ datapath.ru.latched_instruction\[7\] vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_44_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_clk sky130_fd_sc_hd__clkbuf_8
X_08310_ datapath.rf.registers\[26\]\[4\] net836 _03144_ _03145_ vssd1 vssd1 vccd1
+ vccd1 _03146_ sky130_fd_sc_hd__a211o_1
XFILLER_61_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08103__A2 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09290_ _04032_ _04125_ net374 vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__mux2_1
XFILLER_33_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08241_ _01595_ _01784_ vssd1 vssd1 vccd1 vccd1 _03077_ sky130_fd_sc_hd__nor2_1
XANTENNA_14 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08172_ net582 _03007_ datapath.rf.registers\[0\]\[7\] net867 vssd1 vssd1 vccd1 vccd1
+ _03008_ sky130_fd_sc_hd__o2bb2a_4
XANTENNA__06980__X _01816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09603__A2 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07123_ datapath.rf.registers\[16\]\[28\] _01707_ net930 vssd1 vssd1 vccd1 vccd1
+ _01959_ sky130_fd_sc_hd__and3_1
XFILLER_146_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07054_ datapath.rf.registers\[16\]\[30\] net740 net720 datapath.rf.registers\[20\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__a22o_1
XANTENNA__07090__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 WE_O sky130_fd_sc_hd__buf_2
Xoutput121 net121 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
XANTENNA__07378__B1 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07917__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09119__A1 _02217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout486_A _06552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07956_ datapath.rf.registers\[9\]\[11\] net886 net881 datapath.rf.registers\[10\]\[11\]
+ _02779_ vssd1 vssd1 vccd1 vccd1 _02792_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_145_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06907_ net977 _01720_ vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__and2_4
XFILLER_46_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07887_ _02716_ _02718_ _02720_ _02722_ vssd1 vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout653_A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_106_Right_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09626_ net371 _04379_ vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__nor2_1
XANTENNA__14354__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06838_ datapath.ru.latched_instruction\[29\] _01497_ net1016 net994 vssd1 vssd1
+ vccd1 vccd1 _01674_ sky130_fd_sc_hd__and4b_1
XFILLER_16_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07550__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09557_ net607 _04339_ vssd1 vssd1 vccd1 vccd1 _04393_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout820_A _01756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06769_ _01571_ _01589_ vssd1 vssd1 vccd1 vccd1 _01606_ sky130_fd_sc_hd__nor2_1
XANTENNA__12809__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09827__C1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout539_X net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_35_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout918_A _01764_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08508_ datapath.rf.registers\[19\]\[1\] _01797_ net907 vssd1 vssd1 vccd1 vccd1 _03344_
+ sky130_fd_sc_hd__and3_1
X_09488_ net463 net441 _04322_ net366 vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__o211a_1
XANTENNA__13853__RESET_B net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08439_ datapath.rf.registers\[25\]\[2\] net729 net720 datapath.rf.registers\[20\]\[2\]
+ _03273_ vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__a221o_1
XFILLER_12_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout706_X net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11450_ net1746 net292 net406 vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__mux2_1
XANTENNA__06890__X _01726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09055__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10401_ _05225_ _05233_ _05236_ vssd1 vssd1 vccd1 vccd1 _05237_ sky130_fd_sc_hd__or3_1
XFILLER_137_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11381_ net1809 net301 net410 vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__mux2_1
X_13120_ net196 net1894 net471 vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__mux2_1
XFILLER_125_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10332_ datapath.PC\[14\] _04239_ net467 vssd1 vssd1 vccd1 vccd1 _05168_ sky130_fd_sc_hd__mux2_1
XANTENNA__07081__A2 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10572__B _02660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13051_ net212 net1976 net475 vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__mux2_1
X_10263_ net635 _04272_ vssd1 vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__and2_1
XFILLER_127_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12002_ screen.register.currentYbus\[1\] _05778_ net995 screen.register.currentXbus\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06046_ sky130_fd_sc_hd__a22o_1
XANTENNA__07908__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10194_ net223 _05029_ net1294 vssd1 vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__a21o_1
XANTENNA__10999__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08581__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout370 net371 vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__buf_2
Xfanout381 _03618_ vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__buf_2
XFILLER_143_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08869__A0 _02913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout392 net393 vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__clkbuf_8
X_13953_ clknet_leaf_104_clk _00731_ net1225 vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__dfrtp_1
X_12904_ net1580 net280 net485 vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__mux2_1
X_13884_ clknet_leaf_54_clk _00688_ net1180 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[28\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07541__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06895__A2 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12835_ net297 net2251 net486 vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__mux2_1
XFILLER_15_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_26_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_8
X_12766_ net286 net1575 net497 vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__mux2_1
XFILLER_15_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10747__B _01663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14505_ clknet_leaf_21_clk _01210_ net1163 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11717_ net3 net1036 net1025 net2373 vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__a22o_1
X_12697_ datapath.mulitply_result\[31\] datapath.multiplication_module.multiplicand_i\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06528_ sky130_fd_sc_hd__xnor2_1
X_11648_ net1001 _05830_ _05867_ _05350_ _05871_ vssd1 vssd1 vccd1 vccd1 _05872_ sky130_fd_sc_hd__a221o_1
X_14436_ clknet_leaf_20_clk _01141_ net1119 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput12 DAT_I[19] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
Xinput23 DAT_I[29] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
Xinput34 en vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_96_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11579_ net1270 _01425_ _05801_ _05802_ vssd1 vssd1 vccd1 vccd1 _05803_ sky130_fd_sc_hd__or4b_1
X_14367_ clknet_leaf_13_clk _01072_ net1080 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold807 datapath.rf.registers\[13\]\[9\] vssd1 vssd1 vccd1 vccd1 net2155 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13318_ clknet_leaf_28_clk _00128_ net1133 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold818 datapath.rf.registers\[6\]\[0\] vssd1 vssd1 vccd1 vccd1 net2166 sky130_fd_sc_hd__dlygate4sd3_1
Xhold829 datapath.rf.registers\[11\]\[22\] vssd1 vssd1 vccd1 vccd1 net2177 sky130_fd_sc_hd__dlygate4sd3_1
X_14298_ clknet_leaf_135_clk _01003_ net1102 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13249_ clknet_leaf_46_clk _00059_ net1147 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08021__A1 datapath.rf.registers\[0\]\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07810_ _02644_ _02645_ vssd1 vssd1 vccd1 vccd1 _02646_ sky130_fd_sc_hd__or2_1
X_08790_ _03296_ net576 _03624_ vssd1 vssd1 vccd1 vccd1 _03626_ sky130_fd_sc_hd__o21ai_1
XFILLER_69_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12105__B1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07780__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07741_ datapath.rf.registers\[11\]\[16\] net710 net702 datapath.rf.registers\[9\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__a22o_1
XFILLER_38_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08324__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07672_ datapath.rf.registers\[16\]\[17\] net862 net828 datapath.rf.registers\[12\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__a22o_1
XFILLER_38_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06975__X _01811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07532__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09411_ _04245_ _04246_ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__nand2_1
XFILLER_93_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06623_ _01459_ _01460_ vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_140_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_17_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_34_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09342_ _04150_ _04176_ _04148_ vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__a21o_1
XFILLER_40_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09285__B1 _03604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09824__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09273_ _01609_ _04108_ _03770_ vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__o21ai_1
XFILLER_138_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout234_A _05623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08224_ datapath.rf.registers\[3\]\[6\] net770 net762 datapath.rf.registers\[1\]\[6\]
+ _03058_ vssd1 vssd1 vccd1 vccd1 _03060_ sky130_fd_sc_hd__a221o_1
XFILLER_138_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07031__B net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10944__Y _05684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08155_ datapath.rf.registers\[8\]\[7\] net878 net800 datapath.rf.registers\[15\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02991_ sky130_fd_sc_hd__a22o_1
XFILLER_146_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1143_A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07599__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07106_ datapath.rf.registers\[1\]\[29\] net762 net719 datapath.rf.registers\[20\]\[29\]
+ _01941_ vssd1 vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__a221o_1
XFILLER_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07063__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08086_ datapath.rf.registers\[17\]\[9\] net748 net732 datapath.rf.registers\[19\]\[9\]
+ _02921_ vssd1 vssd1 vccd1 vccd1 _02922_ sky130_fd_sc_hd__a221o_1
X_07037_ datapath.rf.registers\[30\]\[30\] net973 net919 vssd1 vssd1 vccd1 vccd1 _01873_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_58_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout770_A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout391_X net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout489_X net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08289__S net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08988_ net632 net609 vssd1 vssd1 vccd1 vccd1 _03824_ sky130_fd_sc_hd__nor2_2
XANTENNA__07771__B1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07939_ datapath.rf.registers\[11\]\[11\] net987 net938 vssd1 vssd1 vccd1 vccd1 _02775_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08315__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10950_ net169 net2591 net545 vssd1 vssd1 vccd1 vccd1 _00033_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06885__X _01721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07523__B1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11951__B screen.counter.ack vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09609_ net331 _04034_ _04444_ _03613_ vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__o211a_1
X_10881_ datapath.PC\[21\] net1265 _05617_ vssd1 vssd1 vccd1 vccd1 _05629_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout823_X net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12620_ _06461_ _06462_ _06463_ _06457_ vssd1 vssd1 vccd1 vccd1 _06464_ sky130_fd_sc_hd__a211o_1
XANTENNA__09815__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12551_ datapath.mulitply_result\[7\] datapath.multiplication_module.multiplicand_i\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06406_ sky130_fd_sc_hd__nor2_1
XANTENNA__10830__A0 _04239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11502_ net199 net1964 net511 vssd1 vssd1 vccd1 vccd1 _00538_ sky130_fd_sc_hd__mux2_1
X_12482_ net300 net2185 net507 vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__mux2_1
XFILLER_138_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14221_ clknet_leaf_41_clk _00942_ net1144 vssd1 vssd1 vccd1 vccd1 columns.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_22_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11433_ net206 net1879 net514 vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10583__A _02634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14152_ clknet_leaf_143_clk _00909_ net1093 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11364_ net216 net1869 net519 vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__mux2_1
XFILLER_4_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07054__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13103_ net280 net2331 net472 vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__mux2_1
X_10315_ net1268 _03734_ vssd1 vssd1 vccd1 vccd1 _05151_ sky130_fd_sc_hd__xnor2_1
X_14083_ clknet_leaf_96_clk _00849_ net1226 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11295_ net215 net2164 net522 vssd1 vssd1 vccd1 vccd1 _00343_ sky130_fd_sc_hd__mux2_1
XFILLER_152_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08988__A net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13034_ net295 net2347 net474 vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09436__X _04272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10246_ net1044 _03733_ _05081_ net634 vssd1 vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__a31o_1
Xfanout1110 net1120 vssd1 vssd1 vccd1 vccd1 net1110 sky130_fd_sc_hd__buf_2
XFILLER_67_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1121 _00004_ vssd1 vssd1 vccd1 vccd1 net1121 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10897__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1132 net1139 vssd1 vssd1 vccd1 vccd1 net1132 sky130_fd_sc_hd__buf_2
X_10177_ _05010_ _05011_ _05012_ net1041 net895 vssd1 vssd1 vccd1 vccd1 _05013_ sky130_fd_sc_hd__o221a_1
Xfanout1143 net1153 vssd1 vssd1 vccd1 vccd1 net1143 sky130_fd_sc_hd__clkbuf_2
XFILLER_67_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07762__B1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1154 net1162 vssd1 vssd1 vccd1 vccd1 net1154 sky130_fd_sc_hd__clkbuf_4
Xfanout1165 net1166 vssd1 vssd1 vccd1 vccd1 net1165 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1176 net1177 vssd1 vssd1 vccd1 vccd1 net1176 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_109_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1187 net1188 vssd1 vssd1 vccd1 vccd1 net1187 sky130_fd_sc_hd__clkbuf_4
Xfanout1198 net1204 vssd1 vssd1 vccd1 vccd1 net1198 sky130_fd_sc_hd__buf_2
X_13936_ clknet_leaf_111_clk _00714_ net1198 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07514__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11861__B net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13867_ clknet_leaf_75_clk _00671_ net1242 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_122_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11353__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12818_ net1822 net215 net490 vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__mux2_1
XFILLER_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13798_ clknet_leaf_73_clk _00607_ net1243 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_12749_ net1750 net219 net402 vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__mux2_1
XFILLER_8_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07293__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06971__A net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14419_ clknet_leaf_39_clk _01124_ net1141 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_7_Left_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold604 datapath.rf.registers\[27\]\[28\] vssd1 vssd1 vccd1 vccd1 net1952 sky130_fd_sc_hd__dlygate4sd3_1
Xwire590 _02428_ vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__clkbuf_2
Xhold615 datapath.multiplication_module.multiplicand_i\[9\] vssd1 vssd1 vccd1 vccd1
+ net1963 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold626 datapath.rf.registers\[19\]\[3\] vssd1 vssd1 vccd1 vccd1 net1974 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold637 datapath.rf.registers\[30\]\[30\] vssd1 vssd1 vccd1 vccd1 net1985 sky130_fd_sc_hd__dlygate4sd3_1
Xhold648 datapath.rf.registers\[1\]\[29\] vssd1 vssd1 vccd1 vccd1 net1996 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12912__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold659 datapath.rf.registers\[17\]\[23\] vssd1 vssd1 vccd1 vccd1 net2007 sky130_fd_sc_hd__dlygate4sd3_1
X_09960_ _04765_ _04795_ vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__nand2b_1
Xclkbuf_leaf_6_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_8
X_08911_ net1265 datapath.PC\[23\] _03746_ vssd1 vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__nor3_1
X_09891_ _01703_ _01780_ _01593_ vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__o21ba_1
XANTENNA__09742__A1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08842_ _03358_ _01666_ _03671_ vssd1 vssd1 vccd1 vccd1 _03678_ sky130_fd_sc_hd__mux2_1
Xhold1304 datapath.rf.registers\[28\]\[31\] vssd1 vssd1 vccd1 vccd1 net2652 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_774 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10352__A2 net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08410__B _01712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08773_ net600 net633 vssd1 vssd1 vccd1 vccd1 _03609_ sky130_fd_sc_hd__nor2_1
XFILLER_84_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout184_A _05677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07724_ datapath.rf.registers\[14\]\[16\] net829 net796 datapath.rf.registers\[29\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__a22o_1
XFILLER_38_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07026__B net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_894 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06859__A2 _01571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07655_ _02490_ vssd1 vssd1 vccd1 vccd1 _02491_ sky130_fd_sc_hd__inv_2
XFILLER_81_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11263__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06606_ _01411_ _01441_ _01444_ datapath.ru.latched_instruction\[2\] _01439_ vssd1
+ vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__a221o_1
X_07586_ datapath.rf.registers\[2\]\[19\] net744 net685 datapath.rf.registers\[27\]\[19\]
+ _02421_ vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__a221o_1
XFILLER_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09325_ _02522_ net453 _04159_ vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout1260_A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10812__A0 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09256_ net364 _04090_ _04091_ vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__o21a_1
XANTENNA__07284__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08425__X _03261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06881__A _01656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08207_ datapath.rf.registers\[2\]\[6\] net887 net832 datapath.rf.registers\[30\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03043_ sky130_fd_sc_hd__a22o_1
XFILLER_154_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09187_ net630 _03979_ _03981_ _04022_ vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__a2bb2o_2
XTAP_TAPCELL_ROW_153_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout404_X net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08138_ datapath.rf.registers\[23\]\[8\] net701 net693 datapath.rf.registers\[13\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02974_ sky130_fd_sc_hd__a22o_1
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout985_A net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08069_ datapath.rf.registers\[20\]\[9\] net840 _02889_ _02891_ _02896_ vssd1 vssd1
+ vccd1 vccd1 _02905_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12822__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10100_ net1263 _03748_ datapath.PC\[27\] vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_73_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11080_ net282 net1627 net536 vssd1 vssd1 vccd1 vccd1 _00137_ sky130_fd_sc_hd__mux2_1
XFILLER_150_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06599__Y _01438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout773_X net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10031_ _04809_ _04866_ vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11438__S net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08536__A2 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10879__B1 _05626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07744__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout940_X net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11982_ screen.register.currentYbus\[16\] _05773_ _05786_ screen.register.currentYbus\[24\]
+ _05781_ vssd1 vssd1 vccd1 vccd1 _06027_ sky130_fd_sc_hd__a221o_1
XFILLER_90_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13721_ clknet_leaf_31_clk _00531_ net1124 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10933_ net898 _05673_ vssd1 vssd1 vccd1 vccd1 _05674_ sky130_fd_sc_hd__nor2_1
XANTENNA__10578__A net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10864_ datapath.mulitply_result\[19\] net597 net617 vssd1 vssd1 vccd1 vccd1 _05615_
+ sky130_fd_sc_hd__a21o_1
X_13652_ clknet_leaf_93_clk _00462_ net1211 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_27_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12603_ _06440_ _06444_ _06448_ vssd1 vssd1 vccd1 vccd1 _06450_ sky130_fd_sc_hd__nand3_1
XANTENNA__10865__X _05616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13583_ clknet_leaf_26_clk _00393_ net1135 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10795_ _04537_ _05555_ net901 vssd1 vssd1 vccd1 vccd1 _05556_ sky130_fd_sc_hd__mux2_1
X_12534_ _06386_ _06388_ _06385_ vssd1 vssd1 vccd1 vccd1 _06392_ sky130_fd_sc_hd__o21ba_1
XANTENNA__07275__A2 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06791__A _01585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12465_ net164 _05978_ net126 screen.register.currentXbus\[21\] vssd1 vssd1 vccd1
+ vccd1 _00867_ sky130_fd_sc_hd__a2bb2o_1
X_14204_ clknet_leaf_54_clk datapath.multiplication_module.multiplicand_i_n\[15\]
+ net1179 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11416_ net292 net1768 net514 vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__mux2_1
XANTENNA__09421__A0 _02661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12396_ net1381 net131 _06345_ vssd1 vssd1 vccd1 vccd1 _00822_ sky130_fd_sc_hd__a21o_1
X_14135_ clknet_leaf_142_clk _00892_ net1093 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_11347_ net299 net2418 net518 vssd1 vssd1 vccd1 vccd1 _00390_ sky130_fd_sc_hd__mux2_1
XANTENNA__12732__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14066_ clknet_leaf_122_clk _00833_ net1200 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_11278_ net300 net1767 net522 vssd1 vssd1 vccd1 vccd1 _00326_ sky130_fd_sc_hd__mux2_1
XANTENNA__11348__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13017_ net1568 net212 net391 vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__mux2_1
X_10229_ _03750_ _05064_ net1038 vssd1 vssd1 vccd1 vccd1 _05065_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07735__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13956__RESET_B net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1 screen.register.cFill1 vssd1 vssd1 vccd1 vccd1 net1349 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12087__A2 _05773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13919_ clknet_leaf_96_clk _00697_ net1226 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11083__S net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08160__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07440_ datapath.rf.registers\[16\]\[22\] net738 net691 datapath.rf.registers\[13\]\[22\]
+ _02266_ vssd1 vssd1 vccd1 vccd1 _02276_ sky130_fd_sc_hd__a221o_1
XFILLER_90_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07371_ datapath.rf.registers\[18\]\[23\] net790 _02192_ _02206_ vssd1 vssd1 vccd1
+ vccd1 _02207_ sky130_fd_sc_hd__a211oi_1
XANTENNA_max_cap950_A net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12907__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09110_ _03935_ _03939_ _03944_ _03945_ vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_40_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08392__S net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09041_ _03874_ _03876_ net374 vssd1 vssd1 vccd1 vccd1 _03877_ sky130_fd_sc_hd__mux2_1
XANTENNA__10270__B2 net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08405__B net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07018__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold401 datapath.rf.registers\[5\]\[5\] vssd1 vssd1 vccd1 vccd1 net1749 sky130_fd_sc_hd__dlygate4sd3_1
Xhold412 datapath.rf.registers\[13\]\[22\] vssd1 vssd1 vccd1 vccd1 net1760 sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 datapath.rf.registers\[15\]\[24\] vssd1 vssd1 vccd1 vccd1 net1771 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold434 datapath.rf.registers\[12\]\[4\] vssd1 vssd1 vccd1 vccd1 net1782 sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 datapath.rf.registers\[4\]\[5\] vssd1 vssd1 vccd1 vccd1 net1793 sky130_fd_sc_hd__dlygate4sd3_1
Xhold456 datapath.rf.registers\[22\]\[13\] vssd1 vssd1 vccd1 vccd1 net1804 sky130_fd_sc_hd__dlygate4sd3_1
Xhold467 datapath.rf.registers\[24\]\[18\] vssd1 vssd1 vccd1 vccd1 net1815 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07974__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11770__B2 _01908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold478 datapath.rf.registers\[24\]\[28\] vssd1 vssd1 vccd1 vccd1 net1826 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold489 datapath.rf.registers\[26\]\[24\] vssd1 vssd1 vccd1 vccd1 net1837 sky130_fd_sc_hd__dlygate4sd3_1
X_09943_ _01416_ _03265_ vssd1 vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__or2_1
XFILLER_132_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout903 _01625_ vssd1 vssd1 vccd1 vccd1 net903 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout914 _01788_ vssd1 vssd1 vccd1 vccd1 net914 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11258__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout925 net926 vssd1 vssd1 vccd1 vccd1 net925 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout399_A net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout936 _01725_ vssd1 vssd1 vccd1 vccd1 net936 sky130_fd_sc_hd__buf_2
XANTENNA__09715__B2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09874_ _04667_ _04684_ _04709_ vssd1 vssd1 vccd1 vccd1 _04710_ sky130_fd_sc_hd__o21ai_2
Xfanout947 net948 vssd1 vssd1 vccd1 vccd1 net947 sky130_fd_sc_hd__clkbuf_4
Xfanout958 net960 vssd1 vssd1 vccd1 vccd1 net958 sky130_fd_sc_hd__clkbuf_2
Xhold1101 datapath.rf.registers\[12\]\[22\] vssd1 vssd1 vccd1 vccd1 net2449 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1106_A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout969 net970 vssd1 vssd1 vccd1 vccd1 net969 sky130_fd_sc_hd__clkbuf_2
Xhold1112 datapath.rf.registers\[27\]\[21\] vssd1 vssd1 vccd1 vccd1 net2460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1123 datapath.rf.registers\[16\]\[21\] vssd1 vssd1 vccd1 vccd1 net2471 sky130_fd_sc_hd__dlygate4sd3_1
X_08825_ net357 net350 _03660_ vssd1 vssd1 vccd1 vccd1 _03661_ sky130_fd_sc_hd__or3b_2
XFILLER_85_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1134 datapath.rf.registers\[20\]\[11\] vssd1 vssd1 vccd1 vccd1 net2482 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout566_A _01779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1145 datapath.rf.registers\[16\]\[12\] vssd1 vssd1 vccd1 vccd1 net2493 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1156 datapath.rf.registers\[21\]\[16\] vssd1 vssd1 vccd1 vccd1 net2504 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1167 datapath.rf.registers\[25\]\[31\] vssd1 vssd1 vccd1 vccd1 net2515 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1178 datapath.rf.registers\[24\]\[19\] vssd1 vssd1 vccd1 vccd1 net2526 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08756_ _03492_ _03494_ _03591_ vssd1 vssd1 vccd1 vccd1 _03592_ sky130_fd_sc_hd__and3_1
XANTENNA__06876__A _01630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1189 datapath.mulitply_result\[30\] vssd1 vssd1 vccd1 vccd1 net2537 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09252__A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07707_ net612 _02542_ net564 vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__a21oi_2
XANTENNA__11825__A2 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout733_A _01811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08687_ _02660_ _02681_ vssd1 vssd1 vccd1 vccd1 _03523_ sky130_fd_sc_hd__nor2_1
XANTENNA__10398__A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07638_ datapath.rf.registers\[16\]\[18\] net738 net722 datapath.rf.registers\[18\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02474_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout900_A net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout521_X net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07569_ datapath.rf.registers\[16\]\[19\] net862 net843 datapath.rf.registers\[25\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__a22o_1
XANTENNA__12817__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout619_X net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09308_ _04137_ _04138_ _04140_ _04143_ vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__o211ai_1
X_10580_ _02418_ _02466_ _02522_ _02567_ vssd1 vssd1 vccd1 vccd1 _05403_ sky130_fd_sc_hd__or4_1
XANTENNA__09651__B1 _03721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09239_ _03667_ _04073_ _04074_ _04068_ vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__o22a_1
XFILLER_108_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12250_ _06168_ _06241_ _06242_ vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__nor3_1
XANTENNA__07009__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12002__A2 _05778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11201_ net188 net2227 net423 vssd1 vssd1 vccd1 vccd1 _00253_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout988_X net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12181_ _06198_ _06199_ vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__and2_1
XFILLER_135_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11761__B2 _02331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11132_ net198 net2444 net428 vssd1 vssd1 vccd1 vccd1 _00187_ sky130_fd_sc_hd__mux2_1
XFILLER_123_858 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold990 datapath.rf.registers\[15\]\[25\] vssd1 vssd1 vccd1 vccd1 net2338 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_79_Left_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10580__B _02466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11168__S net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08509__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11063_ net197 net2266 net432 vssd1 vssd1 vccd1 vccd1 _00123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07717__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10014_ _04797_ _04849_ vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12069__A2 _05778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14753_ net1291 vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__clkbuf_1
X_11965_ _05751_ _05852_ _05853_ _05777_ _05358_ vssd1 vssd1 vccd1 vccd1 _06011_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_86_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_864 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08142__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13704_ clknet_leaf_65_clk _00514_ net1235 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10916_ net192 net2528 net542 vssd1 vssd1 vccd1 vccd1 _00028_ sky130_fd_sc_hd__mux2_1
XFILLER_72_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14684_ clknet_leaf_8_clk _01389_ net1071 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07496__A2 _02331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11896_ net2481 net160 vssd1 vssd1 vccd1 vccd1 _05961_ sky130_fd_sc_hd__nand2_1
XFILLER_17_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_88_Left_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13635_ clknet_leaf_120_clk _00445_ net1193 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10847_ datapath.PC\[17\] _05593_ vssd1 vssd1 vccd1 vccd1 _05600_ sky130_fd_sc_hd__and2_1
XANTENNA__07248__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13566_ clknet_leaf_148_clk _00376_ net1059 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10778_ net292 net2215 net542 vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__mux2_1
XANTENNA__06952__C net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12517_ _06377_ vssd1 vssd1 vccd1 vccd1 _06378_ sky130_fd_sc_hd__inv_2
X_13497_ clknet_leaf_31_clk _00307_ net1122 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_117_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12448_ net165 _05944_ net127 net2653 vssd1 vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_117_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11867__A _03226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06759__A1 _01503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12379_ _05936_ net159 vssd1 vssd1 vccd1 vccd1 _06337_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_97_Left_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07956__B1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11752__B2 _02771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14118_ clknet_leaf_75_clk net1375 net1246 vssd1 vssd1 vccd1 vccd1 datapath.ru.n_memread2
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07420__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08241__A _01595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11078__S net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06940_ net973 net949 vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__and2_1
XFILLER_86_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14049_ clknet_leaf_100_clk _00816_ net1228 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_06871_ _01630_ _01639_ vssd1 vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__nor2_4
XANTENNA__08381__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08610_ _02683_ _03440_ _03443_ _02682_ vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__a31o_1
X_09590_ _03639_ _04422_ _04423_ _03640_ _04411_ vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__a32o_1
XFILLER_94_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07144__X _01980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08541_ _03374_ _03375_ _03376_ vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__or3_1
XANTENNA__11807__A2 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08133__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08472_ datapath.rf.registers\[9\]\[1\] _01716_ net792 datapath.rf.registers\[18\]\[1\]
+ _03307_ vssd1 vssd1 vccd1 vccd1 _03308_ sky130_fd_sc_hd__a221o_1
XANTENNA__07487__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07423_ datapath.rf.registers\[11\]\[22\] net882 net853 datapath.rf.registers\[19\]\[22\]
+ _02258_ vssd1 vssd1 vccd1 vccd1 _02259_ sky130_fd_sc_hd__a221o_1
XANTENNA__07798__Y _02634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout147_A _05886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07354_ net612 _02189_ net564 vssd1 vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__a21o_2
XANTENNA__07239__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07644__C1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07285_ datapath.rf.registers\[2\]\[25\] net889 net858 datapath.rf.registers\[24\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_150_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1056_A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11991__A1 _05335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09024_ _03488_ net628 _03721_ _03489_ net645 vssd1 vssd1 vccd1 vccd1 _03860_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_150_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold220 datapath.rf.registers\[4\]\[22\] vssd1 vssd1 vccd1 vccd1 net1568 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09397__C1 _03613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12372__S net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold231 datapath.rf.registers\[16\]\[10\] vssd1 vssd1 vccd1 vccd1 net1579 sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 datapath.rf.registers\[21\]\[21\] vssd1 vssd1 vccd1 vccd1 net1590 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1223_A net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12940__A0 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold253 datapath.rf.registers\[3\]\[1\] vssd1 vssd1 vccd1 vccd1 net1601 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 datapath.multiplication_module.multiplicand_i\[21\] vssd1 vssd1 vccd1 vccd1
+ net1612 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11743__B2 _03227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold275 datapath.rf.registers\[21\]\[13\] vssd1 vssd1 vccd1 vccd1 net1623 sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 datapath.rf.registers\[13\]\[21\] vssd1 vssd1 vccd1 vccd1 net1634 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout683_A net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout700 net701 vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__buf_4
Xhold297 datapath.rf.registers\[23\]\[23\] vssd1 vssd1 vccd1 vccd1 net1645 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout711 net713 vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13807__RESET_B net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout722 net725 vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__buf_4
X_09926_ _04761_ vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1011_X net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout733 _01811_ vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__buf_2
Xfanout744 net745 vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__clkbuf_8
Xfanout755 net757 vssd1 vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07990__A _02804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout766 net769 vssd1 vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__buf_4
XANTENNA_fanout850_A _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout777 _01796_ vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__buf_2
X_09857_ _04670_ _04690_ _04692_ vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__o21ai_1
Xfanout788 net789 vssd1 vssd1 vccd1 vccd1 net788 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout471_X net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout799 net800 vssd1 vssd1 vccd1 vccd1 net799 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08372__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08808_ net647 _03642_ vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__or2_4
XFILLER_86_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09788_ _04611_ _04623_ _04609_ vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__a21oi_2
X_08739_ _03524_ _03525_ _03573_ _03522_ vssd1 vssd1 vccd1 vccd1 _03575_ sky130_fd_sc_hd__a31o_1
XANTENNA__12895__X _06554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout736_X net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07478__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11750_ net1524 net143 net138 _02876_ vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__a22o_1
XANTENNA__09872__A0 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10701_ net1467 _03076_ net570 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i_n\[6\]
+ sky130_fd_sc_hd__mux2_1
X_11681_ _05188_ net152 net151 net1441 vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout903_X net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11451__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13420_ clknet_leaf_133_clk _00230_ net1104 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_81_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10632_ _05432_ _05449_ _05450_ _05445_ vssd1 vssd1 vccd1 vccd1 _05452_ sky130_fd_sc_hd__o211a_1
XANTENNA__10575__B _03263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10563_ _05383_ _05384_ _05386_ vssd1 vssd1 vccd1 vccd1 _05387_ sky130_fd_sc_hd__or3_1
X_13351_ clknet_leaf_145_clk _00161_ net1089 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_12302_ net635 _04859_ vssd1 vssd1 vccd1 vccd1 _06282_ sky130_fd_sc_hd__nor2_1
XFILLER_6_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13282_ clknet_leaf_151_clk _00092_ net1052 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10494_ screen.controlBus\[2\] screen.controlBus\[3\] _05314_ _05322_ vssd1 vssd1
+ vccd1 vccd1 _05324_ sky130_fd_sc_hd__and4b_2
XFILLER_108_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12233_ screen.counter.currentCt\[15\] screen.counter.currentCt\[14\] _06228_ vssd1
+ vssd1 vccd1 vccd1 _06232_ sky130_fd_sc_hd__and3_1
XFILLER_108_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12164_ _06189_ _06187_ screen.counter.ct\[11\] vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__mux2_1
XANTENNA__07402__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11115_ net279 net1942 net428 vssd1 vssd1 vccd1 vccd1 _00170_ sky130_fd_sc_hd__mux2_1
XFILLER_111_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12095_ screen.register.currentYbus\[7\] _05778_ _05786_ screen.register.currentYbus\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06133_ sky130_fd_sc_hd__a22o_1
XFILLER_49_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11046_ net280 net1781 net432 vssd1 vssd1 vccd1 vccd1 _00106_ sky130_fd_sc_hd__mux2_1
XFILLER_65_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12997_ net1655 net286 net393 vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__mux2_1
XANTENNA__08115__B1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07124__B net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07469__A2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11948_ _01908_ net656 vssd1 vssd1 vccd1 vccd1 _05996_ sky130_fd_sc_hd__nand2_1
XFILLER_60_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14667_ clknet_leaf_57_clk _01372_ net1161 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11879_ _03028_ net656 vssd1 vssd1 vccd1 vccd1 _05950_ sky130_fd_sc_hd__nand2_1
XANTENNA__11361__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13618_ clknet_leaf_33_clk _00428_ net1125 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14598_ clknet_leaf_29_clk _01303_ net1133 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_13549_ clknet_leaf_138_clk _00359_ net1100 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10776__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07070_ datapath.rf.registers\[28\]\[30\] net752 net736 datapath.rf.registers\[22\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01906_ sky130_fd_sc_hd__a22o_1
XFILLER_145_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07641__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07929__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08402__C net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12920__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07972_ datapath.rf.registers\[11\]\[11\] net712 net673 datapath.rf.registers\[7\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__a22o_1
XFILLER_101_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09711_ net329 _04374_ net332 vssd1 vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__o21a_1
X_06923_ net945 net921 vssd1 vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__and2_1
X_09642_ net454 _04247_ _04281_ net353 vssd1 vssd1 vccd1 vccd1 _04478_ sky130_fd_sc_hd__a211o_1
X_06854_ datapath.ru.latched_instruction\[7\] _01643_ _01673_ net993 _01681_ vssd1
+ vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__a221o_1
X_09573_ net373 _04405_ _04408_ net329 vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__a211o_1
X_06785_ _01610_ net906 vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__nand2_1
XFILLER_83_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout264_A _05575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08524_ net559 _03358_ vssd1 vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__nand2_1
XFILLER_35_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09530__A net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07602__X _02438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08455_ _03282_ _03287_ _03289_ _03290_ vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__nor4_1
XANTENNA_fanout431_A net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1173_A net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11271__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06873__B _01656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout529_A _05721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07406_ _02218_ _02240_ vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_63_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08386_ datapath.rf.registers\[2\]\[3\] net744 net666 datapath.rf.registers\[15\]\[3\]
+ _03221_ vssd1 vssd1 vccd1 vccd1 _03222_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_34_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07880__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08146__A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10395__B net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07337_ datapath.rf.registers\[25\]\[24\] net727 net719 datapath.rf.registers\[20\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__a22o_1
XANTENNA__11964__A1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07268_ datapath.rf.registers\[21\]\[25\] net947 net924 vssd1 vssd1 vccd1 vccd1 _02104_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07632__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout898_A _01626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09007_ _01980_ net553 net549 vssd1 vssd1 vccd1 vccd1 _03843_ sky130_fd_sc_hd__or3_1
X_07199_ datapath.rf.registers\[19\]\[27\] net731 net665 datapath.rf.registers\[15\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02035_ sky130_fd_sc_hd__a22o_1
XFILLER_145_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout686_X net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12830__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout530 net531 vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09137__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout541 _05709_ vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__buf_4
X_09909_ datapath.PC\[14\] _04744_ vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__and2_1
Xfanout552 _03654_ vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__buf_2
Xfanout563 _02264_ vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout853_X net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout574 net575 vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__buf_2
XFILLER_19_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11446__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12920_ net2210 net201 net483 vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__mux2_1
XFILLER_74_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout596 _01785_ vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__clkbuf_4
XFILLER_47_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07699__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08896__A1 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12851_ net214 net2465 net486 vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__mux2_1
XFILLER_132_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ mmio.memload_or_instruction\[8\] net1050 net315 net335 net2611 vssd1 vssd1
+ vccd1 vccd1 _00668_ sky130_fd_sc_hd__a32o_1
XFILLER_15_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_83_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ net221 net1934 net494 vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__mux2_1
XFILLER_15_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14521_ clknet_leaf_9_clk _01226_ net1073 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_11733_ net20 net1036 _05889_ net2548 vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__a22o_1
XANTENNA__10586__A _03227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06783__B _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11181__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14452_ clknet_leaf_94_clk _01157_ net1212 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11664_ net1472 _05875_ _05881_ vssd1 vssd1 vccd1 vccd1 _00554_ sky130_fd_sc_hd__a21o_1
XANTENNA__07871__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13403_ clknet_leaf_38_clk _00213_ net1146 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10615_ _05431_ net1013 vssd1 vssd1 vccd1 vccd1 _05435_ sky130_fd_sc_hd__nor2_1
XANTENNA__10873__X _05623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14383_ clknet_leaf_28_clk _01088_ net1134 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11595_ net1009 _05785_ vssd1 vssd1 vccd1 vccd1 _05819_ sky130_fd_sc_hd__or2_2
XFILLER_128_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13334_ clknet_leaf_140_clk _00144_ net1097 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07623__A2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10546_ net570 _05373_ vssd1 vssd1 vccd1 vccd1 datapath.ack_mul sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_114_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13265_ clknet_leaf_41_clk _00075_ net1142 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_142_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10477_ _05305_ _05306_ vssd1 vssd1 vccd1 vccd1 _05307_ sky130_fd_sc_hd__nor2_1
XANTENNA__08503__B _01800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13650__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12216_ screen.counter.currentCt\[9\] screen.counter.currentCt\[8\] _06217_ vssd1
+ vssd1 vccd1 vccd1 _06221_ sky130_fd_sc_hd__and3_1
X_13196_ clknet_leaf_18_clk _00006_ net1109 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12740__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12147_ _06152_ net603 vssd1 vssd1 vccd1 vccd1 _06178_ sky130_fd_sc_hd__nor2_2
XFILLER_2_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11864__B net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12078_ _06115_ _06117_ _05324_ vssd1 vssd1 vccd1 vccd1 _06118_ sky130_fd_sc_hd__o21a_1
XANTENNA__11356__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11029_ net197 net2647 net540 vssd1 vssd1 vccd1 vccd1 _00091_ sky130_fd_sc_hd__mux2_1
XANTENNA__10143__B1 net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06898__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06570_ datapath.ru.latched_instruction\[5\] vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__inv_2
XFILLER_33_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09300__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11091__S net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08240_ _03062_ _03066_ _03075_ net782 datapath.rf.registers\[0\]\[6\] vssd1 vssd1
+ vccd1 vccd1 _03076_ sky130_fd_sc_hd__o32a_4
XANTENNA__07862__A2 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_15 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08171_ _03006_ _02987_ net867 _03003_ vssd1 vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__and4b_1
XANTENNA__12915__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07122_ datapath.rf.registers\[20\]\[28\] net960 net926 vssd1 vssd1 vccd1 vccd1 _01958_
+ sky130_fd_sc_hd__and3_1
XFILLER_119_747 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07614__A2 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08811__A1 _03228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07053_ datapath.rf.registers\[0\]\[30\] net870 _01887_ vssd1 vssd1 vccd1 vccd1 _01889_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_134_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput100 net100 vssd1 vssd1 vccd1 vccd1 DAT_O[5] sky130_fd_sc_hd__buf_2
Xoutput111 net111 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
Xoutput122 net122 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
XANTENNA__09367__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12371__A1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07029__B net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07955_ datapath.rf.registers\[16\]\[11\] net862 net794 datapath.rf.registers\[31\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02791_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_145_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11266__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08327__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout479_A _06556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06906_ datapath.rf.registers\[1\]\[31\] net845 net842 datapath.rf.registers\[25\]\[31\]
+ _01741_ vssd1 vssd1 vccd1 vccd1 _01742_ sky130_fd_sc_hd__a221o_1
XFILLER_96_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07886_ datapath.rf.registers\[2\]\[13\] net743 net672 datapath.rf.registers\[7\]\[13\]
+ _02721_ vssd1 vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__a221o_1
X_09625_ net650 _04460_ net439 vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__a21oi_1
X_06837_ _01671_ _01672_ _01473_ vssd1 vssd1 vccd1 vccd1 _01673_ sky130_fd_sc_hd__or3b_1
XANTENNA__12293__A1_N net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07550__A1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09556_ _03551_ _04391_ _03604_ vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__a21o_1
X_06768_ _01601_ _01603_ _01604_ vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__nor3_1
XANTENNA__09898__C _01630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14649__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08507_ datapath.rf.registers\[5\]\[1\] net970 _01831_ vssd1 vssd1 vccd1 vccd1 _03343_
+ sky130_fd_sc_hd__and3_1
X_06699_ _01409_ _01502_ _01533_ _01535_ _01537_ vssd1 vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__o2111a_1
XANTENNA_fanout813_A net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout434_X net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09487_ net463 net441 _04322_ vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__o21a_1
XFILLER_24_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07051__Y _01887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08438_ datapath.rf.registers\[27\]\[2\] net967 _01816_ vssd1 vssd1 vccd1 vccd1 _03274_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07853__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09055__A1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout601_X net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12825__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08369_ datapath.rf.registers\[0\]\[3\] net868 _03203_ vssd1 vssd1 vccd1 vccd1 _03205_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_149_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07066__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10400_ _03420_ _04678_ _05234_ _05235_ vssd1 vssd1 vccd1 vccd1 _05236_ sky130_fd_sc_hd__o22a_1
X_11380_ net2279 net305 net413 vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__mux2_1
XANTENNA__09460__D1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10331_ datapath.PC\[15\] net1255 _05163_ _05166_ vssd1 vssd1 vccd1 vccd1 _05167_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10572__C _02704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10262_ net890 _04272_ _04582_ vssd1 vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__nor3_1
X_13050_ net216 net1590 net475 vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__mux2_1
XFILLER_152_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout970_X net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12001_ _05759_ _05851_ _05855_ _05846_ vssd1 vssd1 vccd1 vccd1 _06045_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_76_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09763__C1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10193_ _04868_ _05028_ vssd1 vssd1 vccd1 vccd1 _05029_ sky130_fd_sc_hd__nand2_1
XANTENNA__08030__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10373__B1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08318__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout360 net361 vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__buf_2
XFILLER_143_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout371 _03626_ vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__buf_2
XANTENNA__11176__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout382 net383 vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__buf_4
X_13952_ clknet_leaf_99_clk _00730_ net1229 vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__dfrtp_1
XFILLER_47_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout393 _06557_ vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__buf_4
XANTENNA__08869__A1 _02961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12903_ net2259 net283 net485 vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__mux2_1
X_13883_ clknet_leaf_75_clk _00687_ net1246 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[27\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_19_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12834_ net300 net2368 net489 vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__mux2_1
XANTENNA__09818__A0 _01889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ net259 net2096 net497 vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__mux2_1
X_14504_ clknet_leaf_65_clk _01209_ net1235 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11716_ net33 net1034 net1023 net1490 vssd1 vssd1 vccd1 vccd1 _00597_ sky130_fd_sc_hd__o22a_1
XFILLER_15_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07844__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12696_ _06522_ _06526_ vssd1 vssd1 vccd1 vccd1 _06527_ sky130_fd_sc_hd__nand2_1
X_14435_ clknet_leaf_120_clk _01140_ net1192 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11647_ _05846_ _05864_ net1010 _05845_ vssd1 vssd1 vccd1 vccd1 _05871_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12735__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput13 DAT_I[1] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11928__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput24 DAT_I[2] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07057__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput35 gpio_in[5] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__buf_1
X_14366_ clknet_leaf_148_clk _01071_ net1061 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11578_ net1271 net1272 vssd1 vssd1 vccd1 vccd1 _05802_ sky130_fd_sc_hd__and2b_1
XFILLER_6_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold808 datapath.rf.registers\[26\]\[14\] vssd1 vssd1 vccd1 vccd1 net2156 sky130_fd_sc_hd__dlygate4sd3_1
X_13317_ clknet_leaf_114_clk _00127_ net1190 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10529_ _05350_ _05358_ screen.counter.ct\[16\] vssd1 vssd1 vccd1 vccd1 _05359_ sky130_fd_sc_hd__o21ai_1
Xhold819 datapath.rf.registers\[25\]\[0\] vssd1 vssd1 vccd1 vccd1 net2167 sky130_fd_sc_hd__dlygate4sd3_1
X_14297_ clknet_leaf_92_clk _01002_ net1232 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[17\]
+ sky130_fd_sc_hd__dfrtp_4
X_13248_ clknet_leaf_136_clk _00058_ net1088 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_124_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13179_ net2634 vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_96_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06969__A _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08309__B1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11086__S net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07740_ datapath.rf.registers\[17\]\[16\] net746 net722 datapath.rf.registers\[18\]\[16\]
+ _02575_ vssd1 vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__a221o_1
XFILLER_77_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_74_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07671_ datapath.rf.registers\[15\]\[17\] net984 net915 vssd1 vssd1 vccd1 vccd1 _02507_
+ sky130_fd_sc_hd__and3_1
XFILLER_93_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09410_ net551 net547 _02704_ vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__a21o_1
X_06622_ _01459_ _01460_ vssd1 vssd1 vccd1 vccd1 _01461_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_36_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12408__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09341_ _04150_ _04176_ _04148_ vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__a21oi_2
XANTENNA__08088__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08408__B net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07296__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09272_ net346 _04107_ vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__nor2_1
XANTENNA__06991__X _01827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07835__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_132_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08223_ datapath.rf.registers\[14\]\[6\] net774 net742 datapath.rf.registers\[2\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__a22o_1
XANTENNA__07031__C net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07048__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12041__B1 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_12_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08154_ datapath.rf.registers\[12\]\[7\] net955 net920 vssd1 vssd1 vccd1 vccd1 _02990_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_155_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07105_ datapath.rf.registers\[30\]\[29\] net759 net750 datapath.rf.registers\[28\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__a22o_1
XFILLER_146_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08085_ datapath.rf.registers\[23\]\[9\] net700 net693 datapath.rf.registers\[13\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02921_ sky130_fd_sc_hd__a22o_1
XANTENNA__08260__A2 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_147_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1136_A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07036_ datapath.rf.registers\[26\]\[30\] net975 net937 vssd1 vssd1 vccd1 vccd1 _01872_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_58_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_27_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1244_A datapath.mulitply_result\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08012__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07220__B1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09760__A2 _03718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout763_A net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08987_ _03470_ _03487_ vssd1 vssd1 vccd1 vccd1 _03823_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout384_X net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_5_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_5_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_29_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07938_ datapath.rf.registers\[26\]\[11\] net976 net937 vssd1 vssd1 vccd1 vccd1 _02774_
+ sky130_fd_sc_hd__and3_1
XANTENNA__11855__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07869_ datapath.rf.registers\[0\]\[13\] net870 net589 net587 vssd1 vssd1 vccd1 vccd1
+ _02705_ sky130_fd_sc_hd__a2bb2o_2
XANTENNA_fanout930_A _01727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout649_X net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09608_ net376 _04260_ _04443_ net331 vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__o211ai_1
X_10880_ net215 net2532 net542 vssd1 vssd1 vccd1 vccd1 _00023_ sky130_fd_sc_hd__mux2_1
XANTENNA__14021__RESET_B net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_51_Left_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09539_ _03205_ _03263_ net441 vssd1 vssd1 vccd1 vccd1 _04375_ sky130_fd_sc_hd__mux2_1
XANTENNA__08079__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout816_X net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12550_ datapath.mulitply_result\[7\] datapath.multiplication_module.multiplicand_i\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06405_ sky130_fd_sc_hd__and2_1
XFILLER_24_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07826__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11501_ net205 net1719 net510 vssd1 vssd1 vccd1 vccd1 _00537_ sky130_fd_sc_hd__mux2_1
X_12481_ net302 net1850 net508 vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__mux2_1
X_14220_ clknet_leaf_47_clk datapath.multiplication_module.multiplicand_i_n\[31\]
+ net1173 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11432_ net212 net2027 net514 vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10583__B _02680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14151_ clknet_leaf_17_clk _00908_ net1107 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11363_ net231 net2048 net519 vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__mux2_1
XANTENNA__08251__A2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10594__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08053__B net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13102_ net282 net2372 net471 vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__mux2_1
XFILLER_153_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10314_ net1268 net468 net1038 _05149_ vssd1 vssd1 vccd1 vccd1 _05150_ sky130_fd_sc_hd__o211a_1
X_14082_ clknet_leaf_101_clk _00848_ net1227 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_60_Left_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11294_ net232 net2623 net524 vssd1 vssd1 vccd1 vccd1 _00342_ sky130_fd_sc_hd__mux2_1
XANTENNA__08539__B1 _01756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08988__B net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13033_ net301 net1970 net474 vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07892__B net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10245_ datapath.PC\[2\] datapath.PC\[3\] datapath.PC\[4\] vssd1 vssd1 vccd1 vccd1
+ _05081_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10346__B1 net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1100 net1101 vssd1 vssd1 vccd1 vccd1 net1100 sky130_fd_sc_hd__clkbuf_4
XFILLER_154_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1111 net1115 vssd1 vssd1 vccd1 vccd1 net1111 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09165__A net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07211__B1 _01787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10176_ net1264 _03747_ vssd1 vssd1 vccd1 vccd1 _05012_ sky130_fd_sc_hd__xnor2_1
Xfanout1122 net1123 vssd1 vssd1 vccd1 vccd1 net1122 sky130_fd_sc_hd__clkbuf_4
Xfanout1133 net1139 vssd1 vssd1 vccd1 vccd1 net1133 sky130_fd_sc_hd__clkbuf_4
Xfanout1144 net1153 vssd1 vssd1 vccd1 vccd1 net1144 sky130_fd_sc_hd__clkbuf_4
XFILLER_79_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1155 net1162 vssd1 vssd1 vccd1 vccd1 net1155 sky130_fd_sc_hd__clkbuf_4
Xfanout1166 net1186 vssd1 vssd1 vccd1 vccd1 net1166 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_109_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1177 net1178 vssd1 vssd1 vccd1 vccd1 net1177 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1188 net1204 vssd1 vssd1 vccd1 vccd1 net1188 sky130_fd_sc_hd__buf_2
Xfanout190 _06252_ vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__clkbuf_4
Xfanout1199 net1203 vssd1 vssd1 vccd1 vccd1 net1199 sky130_fd_sc_hd__clkbuf_4
X_13935_ clknet_leaf_122_clk _00713_ net1201 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_75_862 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload5_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13866_ clknet_leaf_73_clk _00670_ net1244 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_122_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12817_ net2454 net232 net492 vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__mux2_1
X_13797_ clknet_leaf_52_clk _00606_ net1181 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07817__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12748_ net1535 net241 net404 vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__mux2_1
XANTENNA__12271__B1 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07700__X _02536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12679_ datapath.mulitply_result\[28\] datapath.multiplication_module.multiplicand_i\[28\]
+ vssd1 vssd1 vccd1 vccd1 _06513_ sky130_fd_sc_hd__or2_1
XFILLER_8_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14418_ clknet_leaf_30_clk _01123_ net1124 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08244__A net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10493__B _05314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14349_ clknet_leaf_124_clk _01054_ net1207 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire591 _02041_ vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__clkbuf_1
Xhold605 datapath.rf.registers\[6\]\[4\] vssd1 vssd1 vccd1 vccd1 net1953 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold616 datapath.rf.registers\[19\]\[24\] vssd1 vssd1 vccd1 vccd1 net1964 sky130_fd_sc_hd__dlygate4sd3_1
Xhold627 datapath.rf.registers\[15\]\[22\] vssd1 vssd1 vccd1 vccd1 net1975 sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 screen.counter.currentCt\[8\] vssd1 vssd1 vccd1 vccd1 net1986 sky130_fd_sc_hd__dlygate4sd3_1
Xhold649 datapath.rf.registers\[24\]\[21\] vssd1 vssd1 vccd1 vccd1 net1997 sky130_fd_sc_hd__dlygate4sd3_1
X_08910_ datapath.PC\[21\] _03745_ vssd1 vssd1 vccd1 vccd1 _03746_ sky130_fd_sc_hd__or2_2
XFILLER_98_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09890_ datapath.PC\[20\] net596 vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__xor2_1
XANTENNA__10713__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07202__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08841_ _03296_ _03671_ _03675_ vssd1 vssd1 vccd1 vccd1 _03677_ sky130_fd_sc_hd__o21ai_1
XFILLER_97_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1305 screen.register.currentXbus\[4\] vssd1 vssd1 vccd1 vccd1 net2653 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08410__C net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08772_ net647 net642 _03601_ vssd1 vssd1 vccd1 vccd1 _03608_ sky130_fd_sc_hd__or3b_2
XFILLER_100_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07723_ datapath.rf.registers\[2\]\[16\] net887 net885 datapath.rf.registers\[9\]\[16\]
+ _02558_ vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_108_Left_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07026__C net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout177_A _05670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07654_ _02467_ _02488_ vssd1 vssd1 vccd1 vccd1 _02490_ sky130_fd_sc_hd__and2_1
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06605_ mmio.key_data\[2\] net1048 _01442_ vssd1 vssd1 vccd1 vccd1 _01444_ sky130_fd_sc_hd__o21ai_2
XANTENNA__07323__A net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07585_ datapath.rf.registers\[12\]\[19\] net756 net708 datapath.rf.registers\[10\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__a22o_1
XFILLER_41_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1086_A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09324_ _02522_ net452 _04159_ vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07808__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09255_ net563 _03761_ _04029_ net367 vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout511_A _05735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout132_X net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08481__A2 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1253_A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout609_A _03607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08206_ datapath.rf.registers\[9\]\[6\] net885 net836 datapath.rf.registers\[26\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_117_Left_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09186_ net609 _03979_ _04021_ net605 vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__a211oi_1
XFILLER_147_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08137_ datapath.rf.registers\[6\]\[8\] net681 net663 datapath.rf.registers\[5\]\[8\]
+ _02972_ vssd1 vssd1 vccd1 vccd1 _02973_ sky130_fd_sc_hd__a221o_1
XANTENNA__08233__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1139_X net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07441__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08068_ datapath.rf.registers\[5\]\[9\] net820 _02887_ _02888_ _02890_ vssd1 vssd1
+ vccd1 vccd1 _02904_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout880_A net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout599_X net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout978_A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07019_ _01854_ vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__inv_2
XFILLER_68_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10030_ _04736_ _04737_ vssd1 vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_8_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10879__A1 _01505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout766_X net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_126_Left_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06896__X _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11981_ _06021_ _06024_ _06025_ vssd1 vssd1 vccd1 vccd1 _06026_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout933_X net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11454__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13720_ clknet_leaf_5_clk _00530_ net1069 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10932_ _05671_ _05672_ vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__or2_1
XFILLER_140_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10578__B _01889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13651_ clknet_leaf_33_clk _00461_ net1129 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10863_ _04118_ _05613_ net902 vssd1 vssd1 vccd1 vccd1 _05614_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_27_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12602_ _06440_ _06444_ _06448_ vssd1 vssd1 vccd1 vccd1 _06449_ sky130_fd_sc_hd__a21o_1
X_13582_ clknet_leaf_0_clk _00392_ net1055 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10794_ datapath.PC\[9\] _05548_ vssd1 vssd1 vccd1 vccd1 _05555_ sky130_fd_sc_hd__xnor2_1
XFILLER_9_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12533_ datapath.mulitply_result\[4\] datapath.multiplication_module.multiplicand_i\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06391_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_135_Left_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08472__A2 _01716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06791__B net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12005__B1 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12464_ net164 _05976_ net126 screen.register.currentXbus\[20\] vssd1 vssd1 vccd1
+ vccd1 _00866_ sky130_fd_sc_hd__a2bb2o_1
X_14203_ clknet_leaf_70_clk datapath.multiplication_module.multiplicand_i_n\[14\]
+ net1244 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_11415_ net296 datapath.rf.registers\[24\]\[5\] net515 vssd1 vssd1 vccd1 vccd1 _00455_
+ sky130_fd_sc_hd__mux2_1
XFILLER_126_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08224__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12395_ _05952_ net158 vssd1 vssd1 vccd1 vccd1 _06345_ sky130_fd_sc_hd__nor2_1
XANTENNA__09421__A1 _02705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07432__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14134_ clknet_leaf_20_clk _00891_ net1118 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11346_ net304 net2640 net520 vssd1 vssd1 vccd1 vccd1 _00389_ sky130_fd_sc_hd__mux2_1
XFILLER_152_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14065_ clknet_leaf_122_clk _00832_ net1200 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_11277_ net302 net1758 net525 vssd1 vssd1 vccd1 vccd1 _00325_ sky130_fd_sc_hd__mux2_1
X_13016_ net1725 net217 net390 vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__mux2_1
XANTENNA__09724__A2 _04556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10228_ datapath.PC\[28\] _03749_ vssd1 vssd1 vccd1 vccd1 _05064_ sky130_fd_sc_hd__nand2_1
XFILLER_95_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10159_ _04874_ _04994_ vssd1 vssd1 vccd1 vccd1 _04995_ sky130_fd_sc_hd__or2_1
Xhold2 screen.register.xFill1 vssd1 vssd1 vccd1 vccd1 net1350 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11872__B net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09488__A1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11364__S net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13918_ clknet_leaf_101_clk _00696_ net1227 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13849_ clknet_leaf_68_clk mmio.ack_center.key_en net1245 vssd1 vssd1 vccd1 vccd1
+ mmio.key_en1 sky130_fd_sc_hd__dfrtp_1
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07370_ net872 _02203_ _02204_ _02205_ vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__or4_1
XANTENNA__08999__A0 _01980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10775__Y _05539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09040_ _03835_ _03875_ net367 vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__mux2_1
XFILLER_136_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08405__C net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12923__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold402 datapath.rf.registers\[15\]\[18\] vssd1 vssd1 vccd1 vccd1 net1750 sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 datapath.rf.registers\[22\]\[27\] vssd1 vssd1 vccd1 vccd1 net1761 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07423__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold424 datapath.rf.registers\[1\]\[22\] vssd1 vssd1 vccd1 vccd1 net1772 sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 datapath.rf.registers\[10\]\[13\] vssd1 vssd1 vccd1 vccd1 net1783 sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 datapath.rf.registers\[2\]\[1\] vssd1 vssd1 vccd1 vccd1 net1794 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08702__A _02912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10951__B _01663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold457 datapath.rf.registers\[13\]\[15\] vssd1 vssd1 vccd1 vccd1 net1805 sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 datapath.rf.registers\[29\]\[12\] vssd1 vssd1 vccd1 vccd1 net1816 sky130_fd_sc_hd__dlygate4sd3_1
X_09942_ _04776_ _04777_ vssd1 vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__nand2b_1
Xhold479 datapath.rf.registers\[23\]\[5\] vssd1 vssd1 vccd1 vccd1 net1827 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout904 _01620_ vssd1 vssd1 vccd1 vccd1 net904 sky130_fd_sc_hd__clkbuf_4
XFILLER_131_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout915 net916 vssd1 vssd1 vccd1 vccd1 net915 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout926 _01739_ vssd1 vssd1 vccd1 vccd1 net926 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09873_ net623 _04706_ _04707_ _04708_ vssd1 vssd1 vccd1 vccd1 _04709_ sky130_fd_sc_hd__o211a_1
Xfanout937 _01720_ vssd1 vssd1 vccd1 vccd1 net937 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout948 _01714_ vssd1 vssd1 vccd1 vccd1 net948 sky130_fd_sc_hd__buf_2
XANTENNA_fanout294_A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout959 net960 vssd1 vssd1 vccd1 vccd1 net959 sky130_fd_sc_hd__clkbuf_4
X_08824_ net456 _03659_ vssd1 vssd1 vccd1 vccd1 _03660_ sky130_fd_sc_hd__nor2_1
Xhold1102 datapath.rf.registers\[11\]\[19\] vssd1 vssd1 vccd1 vccd1 net2450 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1113 datapath.rf.registers\[27\]\[14\] vssd1 vssd1 vccd1 vccd1 net2461 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07037__B net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1124 datapath.rf.registers\[31\]\[16\] vssd1 vssd1 vccd1 vccd1 net2472 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1135 datapath.rf.registers\[20\]\[19\] vssd1 vssd1 vccd1 vccd1 net2483 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1146 datapath.rf.registers\[27\]\[19\] vssd1 vssd1 vccd1 vccd1 net2494 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09533__A net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1157 datapath.rf.registers\[14\]\[25\] vssd1 vssd1 vccd1 vccd1 net2505 sky130_fd_sc_hd__dlygate4sd3_1
X_08755_ _03497_ _03499_ _03588_ _03495_ _03493_ vssd1 vssd1 vccd1 vccd1 _03591_ sky130_fd_sc_hd__a311o_1
Xhold1168 datapath.rf.registers\[5\]\[25\] vssd1 vssd1 vccd1 vccd1 net2516 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1179 datapath.rf.registers\[0\]\[9\] vssd1 vssd1 vccd1 vccd1 net2527 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout559_A _03320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11274__S net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10089__A2 _03914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07706_ datapath.rf.registers\[0\]\[17\] net785 _02536_ _02541_ vssd1 vssd1 vccd1
+ vccd1 _02542_ sky130_fd_sc_hd__o22a_4
X_08686_ _02660_ _02681_ vssd1 vssd1 vccd1 vccd1 _03522_ sky130_fd_sc_hd__and2_1
X_07637_ datapath.rf.registers\[9\]\[18\] net702 net675 datapath.rf.registers\[29\]\[18\]
+ _02472_ vssd1 vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__a221o_1
XFILLER_54_887 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout726_A _01812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout347_X net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06892__A _01707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07568_ datapath.rf.registers\[14\]\[19\] net985 net919 vssd1 vssd1 vccd1 vccd1 _02404_
+ sky130_fd_sc_hd__and3_1
X_09307_ net904 _04119_ _04142_ net317 _04141_ vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout514_X net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07499_ datapath.rf.registers\[15\]\[20\] net982 net915 vssd1 vssd1 vccd1 vccd1 _02335_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09651__A1 _03008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10797__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09238_ net647 _04073_ _03770_ vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__o21a_1
XFILLER_5_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08206__A2 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09169_ _03791_ _03794_ net450 vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__mux2_1
XANTENNA__09403__A1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12833__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11200_ net192 net2157 net422 vssd1 vssd1 vccd1 vccd1 _00252_ sky130_fd_sc_hd__mux2_1
XFILLER_108_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07414__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12180_ net1270 _06164_ _06172_ screen.counter.ct\[18\] vssd1 vssd1 vccd1 vccd1 _06199_
+ sky130_fd_sc_hd__a31o_1
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout883_X net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11449__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11131_ net200 net2118 net427 vssd1 vssd1 vccd1 vccd1 _00186_ sky130_fd_sc_hd__mux2_1
XFILLER_150_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12134__A _06168_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold980 datapath.rf.registers\[24\]\[0\] vssd1 vssd1 vccd1 vccd1 net2328 sky130_fd_sc_hd__dlygate4sd3_1
Xhold991 datapath.rf.registers\[9\]\[23\] vssd1 vssd1 vccd1 vccd1 net2339 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10580__C _02522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11062_ net200 net2293 net431 vssd1 vssd1 vccd1 vccd1 _00122_ sky130_fd_sc_hd__mux2_1
XFILLER_150_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08050__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10013_ _04763_ _04764_ vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__nand2_1
XANTENNA__07193__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08390__A1 datapath.rf.registers\[0\]\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input22_A DAT_I[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08985__C _03779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11184__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06786__B net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14752_ net1291 vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__clkbuf_1
XFILLER_45_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11964_ net1001 _06002_ _06008_ _06009_ vssd1 vssd1 vccd1 vccd1 _06010_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_86_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13703_ clknet_leaf_142_clk _00513_ net1086 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10915_ _05658_ _05657_ net652 _01503_ vssd1 vssd1 vccd1 vccd1 _05659_ sky130_fd_sc_hd__o2bb2a_4
XFILLER_45_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14683_ clknet_leaf_38_clk _01388_ net1145 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_11895_ net134 _05960_ _05959_ vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__o21ai_1
XFILLER_60_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_143_Left_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13634_ clknet_leaf_151_clk _00444_ net1052 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10846_ net245 net2015 net542 vssd1 vssd1 vccd1 vccd1 _00018_ sky130_fd_sc_hd__mux2_1
X_13565_ clknet_leaf_149_clk _00375_ net1060 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10777_ _01486_ net619 _05539_ _05540_ vssd1 vssd1 vccd1 vccd1 _05541_ sky130_fd_sc_hd__a22o_2
XANTENNA__08445__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12516_ datapath.mulitply_result\[0\] datapath.multiplication_module.multiplicand_i\[0\]
+ _06376_ vssd1 vssd1 vccd1 vccd1 _06377_ sky130_fd_sc_hd__and3_1
X_13496_ clknet_leaf_4_clk _00306_ net1076 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_12447_ net167 _05942_ net129 screen.register.currentXbus\[3\] vssd1 vssd1 vccd1
+ vccd1 _00849_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_117_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12743__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11867__B screen.counter.ack vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12378_ net656 net156 vssd1 vssd1 vccd1 vccd1 _06336_ sky130_fd_sc_hd__and2_1
XANTENNA__06759__A2 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11359__S net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14117_ clknet_leaf_78_clk datapath.multiplication_module.zero_multi net1246 vssd1
+ vssd1 vccd1 vccd1 datapath.ru.zero_multi1 sky130_fd_sc_hd__dfrtp_1
X_11329_ net1633 net231 net414 vssd1 vssd1 vccd1 vccd1 _00374_ sky130_fd_sc_hd__mux2_1
XFILLER_141_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08241__B _01784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10490__C _05314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14048_ clknet_leaf_100_clk _00815_ net1228 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06870_ _01579_ _01703_ vssd1 vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__nand2_4
XANTENNA__07184__A2 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13871__Q datapath.ru.latched_instruction\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06696__B net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11094__S net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06931__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08540_ datapath.rf.registers\[22\]\[0\] net823 _01772_ datapath.rf.registers\[15\]\[0\]
+ _03363_ vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__a221o_1
X_08471_ datapath.rf.registers\[25\]\[1\] net843 net803 datapath.rf.registers\[3\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03307_ sky130_fd_sc_hd__a22o_1
XANTENNA__12918__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07422_ datapath.rf.registers\[16\]\[22\] net860 net841 datapath.rf.registers\[25\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__a22o_1
XFILLER_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07353_ _02179_ _02185_ _02188_ net784 datapath.rf.registers\[0\]\[24\] vssd1 vssd1
+ vccd1 vccd1 _02189_ sky130_fd_sc_hd__o32a_4
X_07284_ datapath.rf.registers\[17\]\[25\] net851 net847 datapath.rf.registers\[1\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_150_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09023_ _03857_ _03858_ net319 vssd1 vssd1 vccd1 vccd1 _03859_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_150_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1049_A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold210 datapath.rf.registers\[31\]\[2\] vssd1 vssd1 vccd1 vccd1 net1558 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold221 datapath.rf.registers\[5\]\[0\] vssd1 vssd1 vccd1 vccd1 net1569 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold232 datapath.rf.registers\[16\]\[8\] vssd1 vssd1 vccd1 vccd1 net1580 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11269__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold243 datapath.rf.registers\[10\]\[2\] vssd1 vssd1 vccd1 vccd1 net1591 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold254 datapath.rf.registers\[9\]\[22\] vssd1 vssd1 vccd1 vccd1 net1602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 datapath.rf.registers\[10\]\[3\] vssd1 vssd1 vccd1 vccd1 net1613 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold276 datapath.rf.registers\[21\]\[28\] vssd1 vssd1 vccd1 vccd1 net1624 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1216_A net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold287 datapath.rf.registers\[29\]\[20\] vssd1 vssd1 vccd1 vccd1 net1635 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08151__B net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout701 _01821_ vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__clkbuf_4
Xfanout712 net713 vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__buf_4
Xhold298 datapath.rf.registers\[2\]\[3\] vssd1 vssd1 vccd1 vccd1 net1646 sky130_fd_sc_hd__dlygate4sd3_1
X_09925_ _04758_ _04760_ vssd1 vssd1 vccd1 vccd1 _04761_ sky130_fd_sc_hd__nand2_1
Xfanout723 net725 vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__buf_2
Xfanout734 net737 vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__buf_4
XANTENNA_fanout297_X net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout676_A net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout745 _01807_ vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__clkbuf_4
Xfanout756 net757 vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__buf_4
XANTENNA__10901__S net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout767 net769 vssd1 vssd1 vccd1 vccd1 net767 sky130_fd_sc_hd__clkbuf_4
X_09856_ _04668_ _04691_ _01910_ _03473_ vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__o211a_1
Xfanout778 _01794_ vssd1 vssd1 vccd1 vccd1 net778 sky130_fd_sc_hd__buf_4
XANTENNA__06887__A _01707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07175__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout789 _01790_ vssd1 vssd1 vccd1 vccd1 net789 sky130_fd_sc_hd__buf_2
XFILLER_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08807_ net647 _03642_ vssd1 vssd1 vccd1 vccd1 _03643_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_29_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09787_ net609 _04608_ _04622_ net605 vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__a211oi_1
XANTENNA_fanout464_X net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06999_ net970 _01831_ vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout843_A net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08738_ _03524_ _03525_ _03573_ vssd1 vssd1 vccd1 vccd1 _03574_ sky130_fd_sc_hd__and3_1
XANTENNA__09321__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08124__B2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08669_ _02364_ _02386_ vssd1 vssd1 vccd1 vccd1 _03505_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_101_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout631_X net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12828__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09872__A1 _03669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout729_X net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10700_ net1395 _03123_ net570 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i_n\[5\]
+ sky130_fd_sc_hd__mux2_1
X_11680_ _05116_ net152 net151 net1417 vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__a22o_1
XANTENNA__07883__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10631_ _05450_ vssd1 vssd1 vccd1 vccd1 _05451_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_81_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10575__C net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07635__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13350_ clknet_leaf_11_clk _00160_ net1083 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10562_ screen.register.currentXbus\[29\] screen.register.currentXbus\[28\] screen.register.currentXbus\[31\]
+ screen.register.currentXbus\[30\] vssd1 vssd1 vccd1 vccd1 _05386_ sky130_fd_sc_hd__or4_1
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12301_ _06279_ _06281_ net1266 net308 vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_154_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11982__A2 _05773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13281_ clknet_leaf_45_clk _00091_ net1147 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10493_ screen.controlBus\[3\] _05314_ _05322_ screen.controlBus\[2\] vssd1 vssd1
+ vccd1 vccd1 _05323_ sky130_fd_sc_hd__and4b_1
XANTENNA__09388__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12232_ screen.counter.currentCt\[14\] _06228_ screen.counter.currentCt\[15\] vssd1
+ vssd1 vccd1 vccd1 _06231_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10591__B _02283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11179__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12163_ net1275 _06161_ net601 vssd1 vssd1 vccd1 vccd1 _06189_ sky130_fd_sc_hd__and3_1
XANTENNA__08061__B net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11114_ net284 net2416 net429 vssd1 vssd1 vccd1 vccd1 _00169_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_112_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12094_ _06132_ net1479 _06017_ vssd1 vssd1 vccd1 vccd1 _00733_ sky130_fd_sc_hd__mux2_1
XFILLER_77_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11045_ net283 net2133 net432 vssd1 vssd1 vccd1 vccd1 _00105_ sky130_fd_sc_hd__mux2_1
XFILLER_76_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10170__A1 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07405__B _02240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12996_ net1981 net260 net392 vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__mux2_1
X_11947_ screen.register.currentYbus\[30\] net160 vssd1 vssd1 vccd1 vccd1 _05995_
+ sky130_fd_sc_hd__nand2_1
XFILLER_18_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07124__C net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12738__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07874__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14666_ clknet_leaf_58_clk _01371_ net1167 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11878_ net2518 net161 vssd1 vssd1 vccd1 vccd1 _05949_ sky130_fd_sc_hd__nand2_1
XANTENNA__08076__X _02912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13617_ clknet_leaf_35_clk _00427_ net1127 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10829_ _05583_ _05584_ vssd1 vssd1 vccd1 vccd1 _05585_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_119_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14597_ clknet_leaf_119_clk _01302_ net1191 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08418__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07626__B1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13548_ clknet_leaf_14_clk _00358_ net1103 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08969__A3 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13479_ clknet_leaf_142_clk _00289_ net1086 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09379__B1 _02660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11089__S net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11725__A2 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07971_ datapath.rf.registers\[1\]\[11\] net764 net662 datapath.rf.registers\[5\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__a22o_1
XFILLER_99_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09710_ net328 _04387_ vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__nand2_1
X_06922_ net940 net931 vssd1 vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__and2_2
XFILLER_68_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07157__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09641_ net459 _04307_ _04308_ net349 vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__a211o_1
X_06853_ datapath.ru.latched_instruction\[17\] _01629_ _01682_ _01687_ _01688_ vssd1
+ vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07315__B net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09572_ net362 _04377_ _04404_ net371 vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__o211a_1
X_06784_ _01611_ net904 vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__nor2_1
X_08523_ net610 _03357_ _03324_ vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__o21ai_2
XANTENNA__09811__A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout257_A _05582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06668__B2 datapath.ru.latched_instruction\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_24_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07865__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08454_ _03275_ _03276_ _03277_ _03278_ vssd1 vssd1 vccd1 vccd1 _03290_ sky130_fd_sc_hd__or4_1
XFILLER_11_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07405_ _02218_ _02240_ vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__nand2_1
X_08385_ datapath.rf.registers\[3\]\[3\] net773 net721 datapath.rf.registers\[20\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout424_A net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1166_A net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07336_ datapath.rf.registers\[24\]\[24\] net767 net664 datapath.rf.registers\[15\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__a22o_1
XANTENNA__07617__B1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07267_ datapath.rf.registers\[6\]\[25\] net953 net935 vssd1 vssd1 vccd1 vccd1 _02103_
+ sky130_fd_sc_hd__and3_1
X_09006_ net456 _03840_ _03841_ vssd1 vssd1 vccd1 vccd1 _03842_ sky130_fd_sc_hd__and3_1
XANTENNA__06840__B2 datapath.ru.latched_instruction\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_3_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07198_ datapath.rf.registers\[26\]\[27\] net779 net688 datapath.rf.registers\[31\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02034_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout793_A net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1121_X net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07396__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout520 net521 vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06888__Y _01724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout679_X net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout531 net533 vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__clkbuf_8
Xfanout542 net545 vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__clkbuf_8
XFILLER_59_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09908_ _01611_ _03670_ net604 vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__a21o_1
Xfanout553 _03653_ vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__clkbuf_2
Xfanout564 _01786_ vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__buf_4
XANTENNA__09542__A0 _03009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07148__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout575 _03666_ vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__buf_2
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09839_ _03565_ _04518_ _04673_ _04674_ vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__or4_1
Xfanout597 net599 vssd1 vssd1 vccd1 vccd1 net597 sky130_fd_sc_hd__buf_2
XANTENNA__10152__A1 _04084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout846_X net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12850_ net232 net2017 net488 vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__mux2_1
XFILLER_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09891__B1_N _01593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_83_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ datapath.ru.latched_instruction\[7\] net333 net313 _01642_ vssd1 vssd1 vccd1
+ vccd1 _00667_ sky130_fd_sc_hd__a22o_1
X_12781_ net239 net2181 net496 vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11462__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14520_ clknet_leaf_7_clk _01225_ net1070 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11732_ net19 net1034 net1024 net1462 vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__o22a_1
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07856__B1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08337__A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07320__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10586__B _03292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14451_ clknet_leaf_36_clk _01156_ net1129 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11663_ keypad.apps.app_c\[0\] _05874_ vssd1 vssd1 vccd1 vccd1 _05881_ sky130_fd_sc_hd__and2_1
XFILLER_41_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_153_Right_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13402_ clknet_leaf_146_clk _00212_ net1065 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10614_ _05376_ _05377_ _05378_ vssd1 vssd1 vccd1 vccd1 _05434_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_12_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14382_ clknet_leaf_0_clk _01087_ net1057 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11594_ _05777_ _05783_ _05785_ vssd1 vssd1 vccd1 vccd1 _05818_ sky130_fd_sc_hd__and3_1
X_13333_ clknet_leaf_19_clk _00143_ net1116 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10545_ _05369_ _05370_ _05371_ _05372_ vssd1 vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__or4_1
XFILLER_6_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_130_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_130_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_114_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13264_ clknet_leaf_24_clk _00074_ net1160 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10476_ screen.controlBus\[9\] screen.controlBus\[8\] screen.controlBus\[11\] screen.controlBus\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05306_ sky130_fd_sc_hd__or4_1
XFILLER_136_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11707__A2 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12306__B _06253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12215_ net1986 _06217_ _06220_ vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__o21a_1
XANTENNA__08503__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08033__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13195_ clknet_leaf_58_clk _00005_ net1168 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_135_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12380__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12146_ _06001_ net601 _06176_ screen.counter.ct\[5\] vssd1 vssd1 vccd1 vccd1 _00740_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10391__A1 _03263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12077_ _05752_ _05766_ vssd1 vssd1 vccd1 vccd1 _06117_ sky130_fd_sc_hd__nand2_1
XFILLER_1_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07139__A2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11028_ net202 net1796 net539 vssd1 vssd1 vccd1 vccd1 _00090_ sky130_fd_sc_hd__mux2_1
XFILLER_37_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08887__A2 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14310__Q datapath.rf.registers\[0\]\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12979_ net240 net2522 net480 vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__mux2_1
XFILLER_80_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11372__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14649_ clknet_leaf_30_clk _01354_ net1131 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_120_Right_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_16 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08170_ _02986_ _02993_ _03004_ _03005_ vssd1 vssd1 vccd1 vccd1 _03006_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_31_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06990__A net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07121_ _01935_ _01956_ vssd1 vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_121_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_121_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08272__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07052_ datapath.rf.registers\[0\]\[30\] net870 _01887_ vssd1 vssd1 vccd1 vccd1 _01888_
+ sky130_fd_sc_hd__o21a_2
XFILLER_146_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput101 net101 vssd1 vssd1 vccd1 vccd1 DAT_O[6] sky130_fd_sc_hd__buf_2
Xoutput112 net112 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__buf_2
Xoutput123 net123 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
XANTENNA__08024__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12931__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06989__X _01825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07378__A2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12371__A2 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10382__A1 _03320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08710__A net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07029__C net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07954_ datapath.rf.registers\[1\]\[11\] net847 net843 datapath.rf.registers\[25\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__a22o_1
XFILLER_29_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06905_ datapath.rf.registers\[20\]\[31\] net958 net923 vssd1 vssd1 vccd1 vccd1 _01741_
+ sky130_fd_sc_hd__and3_1
XFILLER_96_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10134__A1 _03729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07885_ datapath.rf.registers\[14\]\[13\] net775 net766 datapath.rf.registers\[24\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02721_ sky130_fd_sc_hd__a22o_1
XFILLER_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09624_ net346 _04000_ _04456_ _04459_ vssd1 vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__a22o_1
X_06836_ _01455_ _01491_ _01508_ _01514_ vssd1 vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__or4_1
XFILLER_56_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07550__A2 _02385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09555_ _03549_ _03550_ vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__or2_1
X_06767_ net1046 net1016 net994 net1029 datapath.ru.latched_instruction\[25\] vssd1
+ vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__a32oi_4
XTAP_TAPCELL_ROW_65_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11282__S net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08506_ datapath.rf.registers\[18\]\[1\] net909 net907 vssd1 vssd1 vccd1 vccd1 _03342_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07838__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09486_ net557 net576 net546 _03204_ vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__o211ai_1
X_06698_ datapath.ru.latched_instruction\[9\] _01536_ vssd1 vssd1 vccd1 vccd1 _01537_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__07302__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08437_ datapath.rf.registers\[19\]\[2\] _01797_ net907 vssd1 vssd1 vccd1 vccd1 _03273_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout427_X net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout806_A _01768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08368_ datapath.rf.registers\[0\]\[3\] net869 _03203_ vssd1 vssd1 vccd1 vccd1 _03204_
+ sky130_fd_sc_hd__o21a_2
X_07319_ datapath.rf.registers\[30\]\[24\] net832 net796 datapath.rf.registers\[29\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__a22o_1
XANTENNA__08263__B1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_112_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_112_clk
+ sky130_fd_sc_hd__clkbuf_8
X_08299_ datapath.rf.registers\[19\]\[4\] net853 net808 datapath.rf.registers\[27\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03135_ sky130_fd_sc_hd__a22o_1
XANTENNA__10832__A1_N _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13002__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10330_ net223 _05165_ net1294 vssd1 vssd1 vccd1 vccd1 _05166_ sky130_fd_sc_hd__a21o_1
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout796_X net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10572__D _02750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08015__B1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10261_ net228 _05096_ vssd1 vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__nor2_1
XANTENNA__12841__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06899__X _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12000_ _05847_ _06043_ vssd1 vssd1 vccd1 vccd1 _06044_ sky130_fd_sc_hd__or2_1
XANTENNA__07369__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12362__A2 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13862__RESET_B net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10192_ _04864_ _04865_ _04867_ vssd1 vssd1 vccd1 vccd1 _05028_ sky130_fd_sc_hd__o21bai_1
XANTENNA__08620__A _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11457__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout350 _03650_ vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__clkbuf_2
Xfanout361 _03646_ vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__clkbuf_2
Xfanout372 net373 vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__buf_2
X_13951_ clknet_leaf_99_clk _00729_ net1228 vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__dfrtp_1
Xfanout383 net385 vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__buf_6
Xfanout394 _06555_ vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__buf_6
XFILLER_19_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12902_ net1658 net293 net482 vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__mux2_1
X_13882_ clknet_leaf_74_clk _00686_ net1242 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[26\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07541__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12833_ net303 net1738 net489 vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09818__A1 _01935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11192__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07829__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12764_ net208 net1616 net496 vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__mux2_1
X_11715_ net32 net1035 net1025 net2541 vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__a22o_1
X_14503_ clknet_leaf_143_clk _01208_ net1086 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10884__X _05632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12695_ net498 _06525_ _06526_ net502 net2537 vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__a32o_1
XFILLER_70_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11646_ _05844_ _05848_ _05865_ _05869_ vssd1 vssd1 vccd1 vccd1 _05870_ sky130_fd_sc_hd__and4_1
X_14434_ clknet_leaf_151_clk _01139_ net1053 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput14 DAT_I[20] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
Xinput25 DAT_I[30] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
X_14365_ clknet_leaf_144_clk _01070_ net1085 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08254__B1 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput36 gpio_in[6] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__buf_1
XFILLER_128_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_103_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_103_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11577_ _01424_ net1274 screen.counter.ct\[19\] screen.counter.ct\[18\] vssd1 vssd1
+ vccd1 vccd1 _05801_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_96_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13316_ clknet_leaf_22_clk _00126_ net1156 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10528_ _05315_ _05357_ vssd1 vssd1 vccd1 vccd1 _05358_ sky130_fd_sc_hd__nor2_2
Xhold809 datapath.rf.registers\[10\]\[26\] vssd1 vssd1 vccd1 vccd1 net2157 sky130_fd_sc_hd__dlygate4sd3_1
X_14296_ clknet_leaf_4_clk _01001_ net1077 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[16\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13247_ clknet_leaf_3_clk _00057_ net1077 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10459_ keypad.decode.sticky\[2\] net1483 net1022 vssd1 vssd1 vccd1 vccd1 keypad.decode.sticky_n\[1\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12751__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06602__X _01441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11875__B net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13178_ net1531 vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11367__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06969__B net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12129_ screen.counter.ct\[19\] screen.counter.ct\[20\] _06165_ vssd1 vssd1 vccd1
+ vccd1 _06166_ sky130_fd_sc_hd__and3_1
XFILLER_111_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09506__B1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07780__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11891__A _02824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07670_ datapath.rf.registers\[2\]\[17\] net984 net949 vssd1 vssd1 vccd1 vccd1 _02506_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07532__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06621_ net1286 net1281 mmio.memload_or_instruction\[3\] vssd1 vssd1 vccd1 vccd1
+ _01460_ sky130_fd_sc_hd__or3_1
XFILLER_53_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09809__A1 _01706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09340_ net609 _04147_ _04175_ net605 vssd1 vssd1 vccd1 vccd1 _04176_ sky130_fd_sc_hd__a211oi_1
XANTENNA__09080__B _03914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08408__C _01712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09271_ net356 _04104_ _04105_ _04099_ vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__o31a_1
XANTENNA__12926__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08222_ datapath.rf.registers\[11\]\[6\] net710 net664 datapath.rf.registers\[15\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03058_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_43_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08705__A net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10954__B _01663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08153_ datapath.rf.registers\[22\]\[7\] net952 net925 vssd1 vssd1 vccd1 vccd1 _02989_
+ sky130_fd_sc_hd__and3_1
XFILLER_107_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07104_ datapath.rf.registers\[4\]\[29\] net714 net680 datapath.rf.registers\[6\]\[29\]
+ _01938_ vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__a221o_1
XANTENNA__07599__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08084_ datapath.rf.registers\[26\]\[9\] net780 net728 datapath.rf.registers\[25\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02920_ sky130_fd_sc_hd__a22o_1
X_07035_ datapath.rf.registers\[31\]\[30\] net973 net916 vssd1 vssd1 vccd1 vccd1 _01871_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1031_A net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_902 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07205__D1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08548__B2 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout491_A _06551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11277__S net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06879__B _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08986_ _03758_ _03821_ net630 vssd1 vssd1 vccd1 vccd1 _03822_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07771__A2 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07937_ _02750_ _02772_ vssd1 vssd1 vccd1 vccd1 _02773_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout756_A net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11855__A1 _04909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07868_ net589 net587 datapath.rf.registers\[0\]\[13\] net870 vssd1 vssd1 vccd1 vccd1
+ _02704_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_84_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07523__A2 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09607_ net370 _04440_ _04442_ net327 vssd1 vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__a211o_1
X_06819_ net1002 net1018 _01654_ vssd1 vssd1 vccd1 vccd1 _01655_ sky130_fd_sc_hd__and3_1
XFILLER_28_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout923_A _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07799_ net610 _02633_ _01787_ vssd1 vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout544_X net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09538_ _04229_ _04373_ net373 vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__mux2_1
XANTENNA__07503__B net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout711_X net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09469_ _02856_ net554 net550 vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__or3_1
XANTENNA__12836__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout809_X net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11500_ net213 net2232 net510 vssd1 vssd1 vccd1 vccd1 _00536_ sky130_fd_sc_hd__mux2_1
X_12480_ net289 net1558 net508 vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__mux2_1
XFILLER_132_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11431_ net214 net1997 net514 vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__mux2_1
XANTENNA__08236__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12032__B2 _05335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09433__C1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10583__C _02725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14150_ clknet_leaf_116_clk _00907_ net1187 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11362_ net237 net2483 net520 vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__mux2_1
X_13101_ net290 net2597 net470 vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__mux2_1
XANTENNA__08053__C net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10313_ net468 _04474_ vssd1 vssd1 vccd1 vccd1 _05149_ sky130_fd_sc_hd__nand2_1
X_14081_ clknet_leaf_97_clk _00847_ net1231 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_125_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11293_ net235 net2159 net524 vssd1 vssd1 vccd1 vccd1 _00341_ sky130_fd_sc_hd__mux2_1
XFILLER_153_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12335__A2 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13032_ net303 net1570 net476 vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10244_ _01417_ net466 net1039 _05079_ vssd1 vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__o211a_1
XANTENNA__07892__C _01744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11187__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1101 net1120 vssd1 vssd1 vccd1 vccd1 net1101 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07211__A1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1112 net1115 vssd1 vssd1 vccd1 vccd1 net1112 sky130_fd_sc_hd__clkbuf_4
X_10175_ net1264 _01701_ net1041 vssd1 vssd1 vccd1 vccd1 _05011_ sky130_fd_sc_hd__o21ai_1
Xfanout1123 net1126 vssd1 vssd1 vccd1 vccd1 net1123 sky130_fd_sc_hd__clkbuf_4
Xfanout1134 net1139 vssd1 vssd1 vccd1 vccd1 net1134 sky130_fd_sc_hd__buf_2
XFILLER_121_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07762__A2 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1145 net1148 vssd1 vssd1 vccd1 vccd1 net1145 sky130_fd_sc_hd__clkbuf_4
Xfanout1156 net1162 vssd1 vssd1 vccd1 vccd1 net1156 sky130_fd_sc_hd__clkbuf_4
XFILLER_66_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1167 net1170 vssd1 vssd1 vccd1 vccd1 net1167 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10879__X _05628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1178 net1185 vssd1 vssd1 vccd1 vccd1 net1178 sky130_fd_sc_hd__clkbuf_2
XFILLER_19_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout191 _06252_ vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__clkbuf_2
Xfanout1189 net1204 vssd1 vssd1 vccd1 vccd1 net1189 sky130_fd_sc_hd__clkbuf_4
XFILLER_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13934_ clknet_leaf_122_clk _00712_ net1203 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07514__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13865_ clknet_leaf_71_clk _00669_ net1244 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_122_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12816_ net2308 net236 net492 vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__mux2_1
XFILLER_90_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13796_ clknet_leaf_52_clk _00605_ net1184 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08475__B1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12747_ net1797 net245 net402 vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__mux2_1
XANTENNA__12746__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12678_ datapath.mulitply_result\[28\] datapath.multiplication_module.multiplicand_i\[28\]
+ vssd1 vssd1 vccd1 vccd1 _06512_ sky130_fd_sc_hd__nand2_1
XANTENNA__08525__A net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14417_ clknet_leaf_41_clk _01122_ net1142 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11629_ screen.counter.ct\[4\] _01423_ _05800_ _05850_ vssd1 vssd1 vccd1 vccd1 _05853_
+ sky130_fd_sc_hd__or4_2
XFILLER_8_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08227__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14348_ clknet_leaf_15_clk _01053_ net1105 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire581 _03291_ vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__clkbuf_2
Xhold606 datapath.rf.registers\[18\]\[3\] vssd1 vssd1 vccd1 vccd1 net1954 sky130_fd_sc_hd__dlygate4sd3_1
Xhold617 datapath.rf.registers\[21\]\[17\] vssd1 vssd1 vccd1 vccd1 net1965 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold628 datapath.rf.registers\[21\]\[22\] vssd1 vssd1 vccd1 vccd1 net1976 sky130_fd_sc_hd__dlygate4sd3_1
Xhold639 datapath.rf.registers\[9\]\[21\] vssd1 vssd1 vccd1 vccd1 net1987 sky130_fd_sc_hd__dlygate4sd3_1
X_14279_ clknet_leaf_143_clk _00984_ net1086 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12481__S net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07428__X _02264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11097__S net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08840_ _03296_ _03671_ _03675_ vssd1 vssd1 vccd1 vccd1 _03676_ sky130_fd_sc_hd__o21a_1
XFILLER_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1306 screen.register.currentXbus\[8\] vssd1 vssd1 vccd1 vccd1 net2654 sky130_fd_sc_hd__dlygate4sd3_1
X_08771_ net651 net643 _03601_ vssd1 vssd1 vccd1 vccd1 _03607_ sky130_fd_sc_hd__and3_2
X_07722_ datapath.rf.registers\[11\]\[16\] net882 net841 datapath.rf.registers\[25\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_4_7_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07653_ _02467_ _02488_ vssd1 vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__nor2_1
XFILLER_25_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06604_ mmio.key_data\[2\] net1048 _01442_ vssd1 vssd1 vccd1 vccd1 _01443_ sky130_fd_sc_hd__o21a_2
XFILLER_92_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07584_ datapath.rf.registers\[1\]\[19\] net764 net728 datapath.rf.registers\[25\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__a22o_1
XFILLER_22_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09323_ net552 net548 _02567_ vssd1 vssd1 vccd1 vccd1 _04159_ sky130_fd_sc_hd__a21o_1
XFILLER_34_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10273__B1 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1079_A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09254_ _02365_ _03761_ _04089_ vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__a21oi_1
X_08205_ datapath.rf.registers\[8\]\[6\] net876 _03035_ _03036_ _03039_ vssd1 vssd1
+ vccd1 vccd1 _03041_ sky130_fd_sc_hd__a2111o_1
XFILLER_138_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08218__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09185_ net317 _04020_ _04015_ _04013_ _04003_ vssd1 vssd1 vccd1 vccd1 _04021_ sky130_fd_sc_hd__o2111a_1
XANTENNA_fanout504_A net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08154__B net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1246_A net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08136_ datapath.rf.registers\[19\]\[8\] net733 net717 datapath.rf.registers\[4\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02972_ sky130_fd_sc_hd__a22o_1
XFILLER_147_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07993__B net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08067_ datapath.rf.registers\[17\]\[9\] net851 net809 datapath.rf.registers\[27\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02903_ sky130_fd_sc_hd__a22o_1
X_07018_ datapath.rf.registers\[0\]\[31\] net784 _01839_ _01853_ vssd1 vssd1 vccd1
+ vccd1 _01854_ sky130_fd_sc_hd__o22ai_4
XTAP_TAPCELL_ROW_73_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout494_X net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout873_A _01723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09194__A1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07744__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout661_X net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08969_ _03082_ _03103_ net447 _03804_ vssd1 vssd1 vccd1 vccd1 _03805_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout759_X net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11980_ _05324_ _06003_ vssd1 vssd1 vccd1 vccd1 _06025_ sky130_fd_sc_hd__and2_1
XFILLER_57_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10931_ datapath.PC\[29\] _05665_ vssd1 vssd1 vccd1 vccd1 _05672_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout926_X net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10578__C _01981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10862_ _05611_ _05612_ vssd1 vssd1 vccd1 vccd1 _05613_ sky130_fd_sc_hd__nor2_1
X_13650_ clknet_leaf_30_clk _00460_ net1132 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_27_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08048__C net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12601_ _06446_ _06447_ vssd1 vssd1 vccd1 vccd1 _06448_ sky130_fd_sc_hd__or2_1
XFILLER_140_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13581_ clknet_leaf_132_clk _00391_ net1113 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10793_ net280 net2100 net543 vssd1 vssd1 vccd1 vccd1 _00010_ sky130_fd_sc_hd__mux2_1
XANTENNA__11470__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12532_ datapath.mulitply_result\[4\] datapath.multiplication_module.multiplicand_i\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06390_ sky130_fd_sc_hd__and2_1
XFILLER_12_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12463_ net166 _05974_ net128 screen.register.currentXbus\[19\] vssd1 vssd1 vccd1
+ vccd1 _00865_ sky130_fd_sc_hd__a2bb2o_1
X_11414_ net298 net2037 net514 vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__mux2_1
X_14202_ clknet_leaf_69_clk datapath.multiplication_module.multiplicand_i_n\[13\]
+ net1245 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_126_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12394_ screen.controlBus\[7\] net133 _06344_ vssd1 vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_73_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14133_ clknet_leaf_93_clk _00890_ net1210 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_126_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11345_ net286 net2068 net521 vssd1 vssd1 vccd1 vccd1 _00388_ sky130_fd_sc_hd__mux2_1
XANTENNA__12308__A2 _06246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07983__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14064_ clknet_leaf_122_clk _00831_ net1200 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_11276_ net286 net1847 net525 vssd1 vssd1 vccd1 vccd1 _00324_ sky130_fd_sc_hd__mux2_1
X_13015_ net1696 net231 net391 vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__mux2_1
X_10227_ datapath.PC\[28\] net468 net1042 vssd1 vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__o21a_1
XANTENNA__07408__B net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_88_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07196__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07735__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10158_ _04834_ _04873_ vssd1 vssd1 vccd1 vccd1 _04994_ sky130_fd_sc_hd__and2b_1
XFILLER_67_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_131_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold3 mmio.WEN1 vssd1 vssd1 vccd1 vccd1 net1351 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10089_ _03868_ _03914_ _01702_ vssd1 vssd1 vccd1 vccd1 _04925_ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_11_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13917_ clknet_leaf_101_clk _00695_ net1227 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_866 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08160__A2 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_146_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13848_ clknet_leaf_78_clk WEN net1245 vssd1 vssd1 vccd1 vccd1 mmio.WEN1 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08448__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_26_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13779_ clknet_leaf_51_clk _00588_ net1181 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11380__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08999__A1 _02025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07120__B1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_4_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_4_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_135_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold403 datapath.rf.registers\[26\]\[23\] vssd1 vssd1 vccd1 vccd1 net1751 sky130_fd_sc_hd__dlygate4sd3_1
Xhold414 datapath.rf.registers\[4\]\[8\] vssd1 vssd1 vccd1 vccd1 net1762 sky130_fd_sc_hd__dlygate4sd3_1
Xhold425 datapath.rf.registers\[26\]\[30\] vssd1 vssd1 vccd1 vccd1 net1773 sky130_fd_sc_hd__dlygate4sd3_1
Xhold436 datapath.rf.registers\[14\]\[4\] vssd1 vssd1 vccd1 vccd1 net1784 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13100__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold447 datapath.rf.registers\[28\]\[5\] vssd1 vssd1 vccd1 vccd1 net1795 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07974__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold458 datapath.rf.registers\[9\]\[9\] vssd1 vssd1 vccd1 vccd1 net1806 sky130_fd_sc_hd__dlygate4sd3_1
Xhold469 mmio.memload_or_instruction\[21\] vssd1 vssd1 vccd1 vccd1 net1817 sky130_fd_sc_hd__dlygate4sd3_1
X_09941_ datapath.PC\[3\] _03206_ vssd1 vssd1 vccd1 vccd1 _04777_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_55_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout905 _01619_ vssd1 vssd1 vccd1 vccd1 net905 sky130_fd_sc_hd__buf_2
Xfanout916 _01771_ vssd1 vssd1 vccd1 vccd1 net916 sky130_fd_sc_hd__clkbuf_4
Xfanout927 _01732_ vssd1 vssd1 vccd1 vccd1 net927 sky130_fd_sc_hd__buf_4
X_09872_ net642 _03669_ _04682_ vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_5_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout938 net939 vssd1 vssd1 vccd1 vccd1 net938 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07726__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout949 net951 vssd1 vssd1 vccd1 vccd1 net949 sky130_fd_sc_hd__buf_4
XANTENNA__08384__C1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1103 datapath.rf.registers\[28\]\[29\] vssd1 vssd1 vccd1 vccd1 net2451 sky130_fd_sc_hd__dlygate4sd3_1
X_08823_ net551 net547 net566 vssd1 vssd1 vccd1 vccd1 _03659_ sky130_fd_sc_hd__a21o_1
Xhold1114 datapath.rf.registers\[20\]\[14\] vssd1 vssd1 vccd1 vccd1 net2462 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07037__C net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06934__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1125 datapath.rf.registers\[11\]\[14\] vssd1 vssd1 vccd1 vccd1 net2473 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1136 datapath.rf.registers\[29\]\[4\] vssd1 vssd1 vccd1 vccd1 net2484 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1147 datapath.rf.registers\[28\]\[16\] vssd1 vssd1 vccd1 vccd1 net2495 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08754_ _03497_ _03499_ _03588_ _03495_ vssd1 vssd1 vccd1 vccd1 _03590_ sky130_fd_sc_hd__a31o_1
Xhold1158 datapath.rf.registers\[22\]\[25\] vssd1 vssd1 vccd1 vccd1 net2506 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1169 datapath.rf.registers\[28\]\[14\] vssd1 vssd1 vccd1 vccd1 net2517 sky130_fd_sc_hd__dlygate4sd3_1
X_07705_ _02531_ _02532_ _02540_ vssd1 vssd1 vccd1 vccd1 _02541_ sky130_fd_sc_hd__or3_1
XFILLER_26_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08685_ _02612_ _02635_ vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__or2_2
Xclkbuf_leaf_92_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_92_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08149__B net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1196_A net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07636_ datapath.rf.registers\[26\]\[18\] net778 net730 datapath.rf.registers\[19\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__a22o_1
XFILLER_54_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08439__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07567_ datapath.rf.registers\[13\]\[19\] net985 net918 vssd1 vssd1 vccd1 vccd1 _02403_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_24_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11290__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06892__B net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout719_A net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09306_ net319 _03908_ vssd1 vssd1 vccd1 vccd1 _04142_ sky130_fd_sc_hd__or2_1
XANTENNA__10246__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07498_ datapath.rf.registers\[25\]\[20\] net973 net943 vssd1 vssd1 vccd1 vccd1 _02334_
+ sky130_fd_sc_hd__and3_1
XFILLER_10_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09237_ net348 _04072_ vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__nor2_1
XANTENNA__07500__C net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout507_X net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1249_X net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09168_ _03781_ _03790_ net450 vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__mux2_1
XFILLER_108_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout990_A _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08119_ datapath.rf.registers\[20\]\[8\] net840 net823 datapath.rf.registers\[22\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__a22o_1
XFILLER_79_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09099_ net574 _03933_ _03934_ _03925_ vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_135_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13010__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11130_ net204 net2339 net426 vssd1 vssd1 vccd1 vccd1 _00185_ sky130_fd_sc_hd__mux2_1
XANTENNA__07965__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold970 datapath.mulitply_result\[27\] vssd1 vssd1 vccd1 vccd1 net2318 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12134__B net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout876_X net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09167__A1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold981 datapath.rf.registers\[26\]\[3\] vssd1 vssd1 vccd1 vccd1 net2329 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10580__D _02567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11061_ net205 net2046 net430 vssd1 vssd1 vccd1 vccd1 _00121_ sky130_fd_sc_hd__mux2_1
Xhold992 datapath.rf.registers\[21\]\[0\] vssd1 vssd1 vccd1 vccd1 net2340 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07178__B1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07717__A2 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10012_ _04846_ _04847_ vssd1 vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__nor2_1
XANTENNA__10721__A1 _03008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06925__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11465__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08390__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10589__B _01908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06786__C net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input15_A DAT_I[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11963_ _05794_ _05797_ net1010 vssd1 vssd1 vccd1 vccd1 _06009_ sky130_fd_sc_hd__a21boi_1
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_83_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_86_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08142__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13702_ clknet_leaf_11_clk _00512_ net1082 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10914_ datapath.mulitply_result\[26\] net597 net618 vssd1 vssd1 vccd1 vccd1 _05658_
+ sky130_fd_sc_hd__a21oi_1
X_11894_ _02771_ net657 vssd1 vssd1 vccd1 vccd1 _05960_ sky130_fd_sc_hd__nand2_1
X_14682_ clknet_leaf_136_clk _01387_ net1091 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07350__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10845_ _05597_ _05598_ _01523_ net617 vssd1 vssd1 vccd1 vccd1 _05599_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_60_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13633_ clknet_leaf_46_clk _00443_ net1171 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10809__S net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13564_ clknet_leaf_7_clk _00374_ net1073 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10776_ datapath.mulitply_result\[6\] net615 net654 vssd1 vssd1 vccd1 vccd1 _05540_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__07102__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11985__B1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08506__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12515_ datapath.mulitply_result\[1\] datapath.multiplication_module.multiplicand_i\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06376_ sky130_fd_sc_hd__xor2_1
X_13495_ clknet_leaf_127_clk _00305_ net1209 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_12446_ net167 _05940_ net129 net2650 vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09458__X _04294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12377_ _04909_ _05073_ _05285_ _05931_ vssd1 vssd1 vccd1 vccd1 _06335_ sky130_fd_sc_hd__or4b_4
XTAP_TAPCELL_ROW_10_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06759__A3 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07956__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14116_ clknet_leaf_78_clk datapath.ack_mul net1245 vssd1 vssd1 vccd1 vccd1 datapath.ru.ack_mul_reg
+ sky130_fd_sc_hd__dfrtp_1
X_11328_ net1852 net238 net417 vssd1 vssd1 vccd1 vccd1 _00373_ sky130_fd_sc_hd__mux2_1
XANTENNA__07419__A net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11259_ net218 net2399 net418 vssd1 vssd1 vccd1 vccd1 _00308_ sky130_fd_sc_hd__mux2_1
X_14047_ clknet_leaf_101_clk _00814_ net1228 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07169__B1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07706__X _02542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10712__A1 _03321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06977__B net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08381__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_74_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08133__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08470_ datapath.rf.registers\[11\]\[1\] net884 net847 datapath.rf.registers\[1\]\[1\]
+ _03305_ vssd1 vssd1 vccd1 vccd1 _03306_ sky130_fd_sc_hd__a221o_1
XANTENNA__07341__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07421_ datapath.rf.registers\[2\]\[22\] net887 net845 datapath.rf.registers\[1\]\[22\]
+ _02256_ vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__a221o_1
X_07352_ _02171_ _02172_ _02186_ _02187_ vssd1 vssd1 vccd1 vccd1 _02188_ sky130_fd_sc_hd__or4_1
XFILLER_148_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07283_ _02115_ _02116_ _02117_ _02118_ vssd1 vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__or4_1
XANTENNA__12934__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09022_ net340 _03713_ vssd1 vssd1 vccd1 vccd1 _03858_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_150_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold200 datapath.rf.registers\[15\]\[0\] vssd1 vssd1 vccd1 vccd1 net1548 sky130_fd_sc_hd__dlygate4sd3_1
Xhold211 columns.count\[1\] vssd1 vssd1 vccd1 vccd1 net1559 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout202_A _05646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08432__B net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold222 datapath.rf.registers\[21\]\[3\] vssd1 vssd1 vccd1 vccd1 net1570 sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 datapath.rf.registers\[25\]\[30\] vssd1 vssd1 vccd1 vccd1 net1581 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 datapath.rf.registers\[22\]\[20\] vssd1 vssd1 vccd1 vccd1 net1592 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 datapath.rf.registers\[4\]\[25\] vssd1 vssd1 vccd1 vccd1 net1603 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold266 datapath.rf.registers\[6\]\[18\] vssd1 vssd1 vccd1 vccd1 net1614 sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 datapath.rf.registers\[13\]\[24\] vssd1 vssd1 vccd1 vccd1 net1625 sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 datapath.rf.registers\[5\]\[29\] vssd1 vssd1 vccd1 vccd1 net1636 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout702 net705 vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__buf_4
Xhold299 datapath.rf.registers\[11\]\[11\] vssd1 vssd1 vccd1 vccd1 net1647 sky130_fd_sc_hd__dlygate4sd3_1
X_09924_ datapath.PC\[10\] _02877_ vssd1 vssd1 vccd1 vccd1 _04760_ sky130_fd_sc_hd__or2_1
Xfanout713 _01817_ vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__clkbuf_4
Xfanout724 net725 vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__buf_4
Xfanout735 net737 vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__clkbuf_4
Xfanout746 net749 vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__buf_4
XANTENNA_input7_A DAT_I[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout757 _01803_ vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__buf_4
X_09855_ _02048_ _02094_ _02049_ vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__o21a_1
XANTENNA__10703__A1 _02980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout571_A _05367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout768 net769 vssd1 vssd1 vccd1 vccd1 net768 sky130_fd_sc_hd__buf_4
Xfanout779 _01794_ vssd1 vssd1 vccd1 vccd1 net779 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11285__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06887__B net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout669_A _01832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08372__A2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08806_ _03601_ _03611_ vssd1 vssd1 vccd1 vccd1 _03642_ sky130_fd_sc_hd__or2_4
XANTENNA__13231__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09786_ _04621_ _04619_ _04615_ vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__and3b_1
X_06998_ net971 _01825_ vssd1 vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_29_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_134_Right_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08737_ _03530_ _03531_ _03570_ _03527_ _03526_ vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__a311o_1
XFILLER_27_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout836_A _01743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_65_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_68_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_68_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08668_ _02312_ _02332_ vssd1 vssd1 vccd1 vccd1 _03504_ sky130_fd_sc_hd__nand2_1
XANTENNA__13887__RESET_B net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07619_ datapath.rf.registers\[23\]\[18\] net813 net799 datapath.rf.registers\[15\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__a22o_1
XANTENNA__09609__C1 _03613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08599_ _02937_ _03434_ _03432_ vssd1 vssd1 vccd1 vccd1 _03435_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout624_X net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13005__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10630_ net122 net123 net124 net121 vssd1 vssd1 vccd1 vccd1 _05450_ sky130_fd_sc_hd__or4b_4
XANTENNA__07511__B net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10575__D net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10561_ screen.register.currentXbus\[25\] screen.register.currentXbus\[24\] screen.register.currentXbus\[27\]
+ screen.register.currentXbus\[26\] vssd1 vssd1 vccd1 vccd1 _05385_ sky130_fd_sc_hd__or4_1
XANTENNA__12844__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08832__B1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12300_ _05571_ _06254_ _06280_ net190 vssd1 vssd1 vccd1 vccd1 _06281_ sky130_fd_sc_hd__o22a_1
XFILLER_139_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13280_ clknet_leaf_133_clk _00090_ net1112 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10492_ screen.controlBus\[0\] screen.controlBus\[1\] _05317_ vssd1 vssd1 vccd1 vccd1
+ _05322_ sky130_fd_sc_hd__nor3_1
XFILLER_108_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12231_ net1518 _06228_ _06230_ vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09388__A1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07399__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10591__C _02331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08342__B net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12162_ _06187_ _06188_ vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__and2_1
XANTENNA__10942__A1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08061__C net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11113_ net292 net1855 net426 vssd1 vssd1 vccd1 vccd1 _00168_ sky130_fd_sc_hd__mux2_1
XFILLER_146_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12093_ _05846_ _05854_ _06124_ _06131_ vssd1 vssd1 vccd1 vccd1 _06132_ sky130_fd_sc_hd__o22a_1
XANTENNA_clkbuf_4_15_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11044_ net292 net2030 net430 vssd1 vssd1 vccd1 vccd1 _00104_ sky130_fd_sc_hd__mux2_1
XANTENNA__11195__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08363__A2 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07571__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12995_ net1578 net207 net392 vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_56_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_18_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08115__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11946_ net134 _05994_ _05993_ vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__o21ai_1
XFILLER_44_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06677__A2 _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14665_ clknet_leaf_62_clk _01370_ net1234 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11877_ net135 _05948_ _05947_ vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__o21ai_1
XFILLER_60_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13616_ clknet_leaf_24_clk _00426_ net1155 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10828_ datapath.PC\[14\] _05576_ vssd1 vssd1 vccd1 vccd1 _05584_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_119_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14596_ clknet_leaf_18_clk _01301_ net1109 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13547_ clknet_leaf_47_clk _00357_ net1171 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12754__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08823__B1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10759_ net1269 datapath.PC\[3\] datapath.PC\[4\] vssd1 vssd1 vccd1 vccd1 _05525_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_146_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11878__B net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13478_ clknet_leaf_17_clk _00288_ net1106 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_132_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12429_ _05986_ net159 vssd1 vssd1 vccd1 vccd1 _06362_ sky130_fd_sc_hd__nor2_1
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07929__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11894__A _02771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07970_ datapath.rf.registers\[10\]\[11\] net708 net693 datapath.rf.registers\[13\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__a22o_1
XANTENNA__06988__A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06921_ datapath.rf.registers\[22\]\[31\] net821 net819 datapath.rf.registers\[5\]\[31\]
+ _01754_ vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_147_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07011__C1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06852_ datapath.ru.latched_instruction\[31\] _01593_ _01648_ datapath.ru.latched_instruction\[10\]
+ _01679_ vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__a221o_1
X_09640_ net359 _04184_ _04190_ vssd1 vssd1 vccd1 vccd1 _04476_ sky130_fd_sc_hd__or3_1
X_09571_ _04154_ _04406_ net372 vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__mux2_1
XFILLER_83_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06783_ _01614_ _01618_ vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__nand2_2
XANTENNA__10797__X _05558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07315__C net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12929__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_47_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_clk sky130_fd_sc_hd__clkbuf_8
X_08522_ net610 _03357_ _03324_ vssd1 vssd1 vccd1 vccd1 _03358_ sky130_fd_sc_hd__o21a_2
XFILLER_51_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08708__A _03205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08453_ datapath.rf.registers\[17\]\[2\] net749 net724 datapath.rf.registers\[18\]\[2\]
+ _03288_ vssd1 vssd1 vccd1 vccd1 _03289_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout152_A net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07404_ net610 net465 _01787_ vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__o21ai_2
X_08384_ datapath.rf.registers\[14\]\[3\] net776 _03219_ net788 vssd1 vssd1 vccd1
+ vccd1 _03220_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_63_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07335_ datapath.rf.registers\[26\]\[24\] net779 net688 datapath.rf.registers\[31\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_63_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout417_A _05726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1159_A net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07093__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07266_ datapath.rf.registers\[7\]\[25\] net941 net934 vssd1 vssd1 vccd1 vccd1 _02102_
+ sky130_fd_sc_hd__and3_1
X_09005_ net551 net547 _01934_ vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__a21o_1
X_07197_ datapath.rf.registers\[16\]\[27\] net739 net672 datapath.rf.registers\[7\]\[27\]
+ _02032_ vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__a221o_1
XFILLER_151_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout786_A net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout510 _05735_ vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__buf_6
Xfanout521 _05728_ vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14015__RESET_B net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09907_ datapath.PC\[15\] net604 _04741_ vssd1 vssd1 vccd1 vccd1 _04743_ sky130_fd_sc_hd__or3_1
Xfanout532 net533 vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__buf_6
XFILLER_99_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout543 net544 vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__buf_4
XFILLER_59_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout554 _03653_ vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout953_A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout565 _01786_ vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09542__A1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout576 _03616_ vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07506__B net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09838_ _03536_ _04273_ vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__nand2b_1
Xfanout598 net599 vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__buf_2
X_09769_ _03978_ _04604_ vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout741_X net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12839__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout839_X net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_38_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_8
X_11800_ datapath.ru.latched_instruction\[6\] net333 net313 _01578_ vssd1 vssd1 vccd1
+ vccd1 _00666_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_83_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ net243 net2207 net494 vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__mux2_1
XFILLER_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07305__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11731_ net18 net1036 _05889_ net2626 vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__a22o_1
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10586__C _03357_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14450_ clknet_leaf_33_clk _01155_ net1124 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11662_ net2326 _05875_ _05880_ vssd1 vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__a21bo_1
XFILLER_30_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13401_ clknet_leaf_9_clk _00211_ net1073 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08056__C net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10613_ net36 _05379_ _05382_ net35 vssd1 vssd1 vccd1 vccd1 _05433_ sky130_fd_sc_hd__and4b_2
X_11593_ screen.counter.ct\[21\] screen.counter.ct\[22\] screen.counter.ct\[20\] vssd1
+ vssd1 vccd1 vccd1 _05817_ sky130_fd_sc_hd__nor3b_1
XTAP_TAPCELL_ROW_12_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14381_ clknet_leaf_125_clk _01086_ net1207 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10544_ datapath.multiplication_module.multiplier_i\[13\] datapath.multiplication_module.multiplier_i\[12\]
+ datapath.multiplication_module.multiplier_i\[15\] datapath.multiplication_module.multiplier_i\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05372_ sky130_fd_sc_hd__or4_1
X_13332_ clknet_leaf_128_clk _00142_ net1209 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10475_ screen.controlBus\[13\] screen.controlBus\[12\] screen.controlBus\[15\] screen.controlBus\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05305_ sky130_fd_sc_hd__or4_1
X_13263_ clknet_leaf_27_clk _00073_ net1131 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12214_ _06168_ _06219_ vssd1 vssd1 vccd1 vccd1 _06220_ sky130_fd_sc_hd__nor2_1
X_13194_ net2601 vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10915__B2 _01503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12145_ net1280 _06177_ _06176_ vssd1 vssd1 vccd1 vccd1 _00739_ sky130_fd_sc_hd__o21a_1
XFILLER_96_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08800__B _01607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07792__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12076_ net1011 _06111_ _06115_ _05330_ _06106_ vssd1 vssd1 vccd1 vccd1 _06116_ sky130_fd_sc_hd__a221o_1
XFILLER_49_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11027_ net204 net1940 net538 vssd1 vssd1 vccd1 vccd1 _00089_ sky130_fd_sc_hd__mux2_1
XANTENNA__07544__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06898__A2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12749__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_29_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_8
X_12978_ net243 net1961 net478 vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_125_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11929_ net2543 net162 vssd1 vssd1 vccd1 vccd1 _05983_ sky130_fd_sc_hd__nand2_1
XANTENNA__08247__B net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14648_ clknet_leaf_6_clk _01353_ net1075 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09049__B1 _02125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13320__RESET_B net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_17 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12484__S net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14579_ clknet_leaf_34_clk _01284_ net1128 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06990__B _01825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07120_ net614 _01954_ net565 vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__a21o_1
XANTENNA__13877__Q datapath.ru.latched_instruction\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07051_ _01875_ _01881_ _01886_ vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__nand3b_4
XFILLER_127_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput102 net102 vssd1 vssd1 vccd1 vccd1 DAT_O[7] sky130_fd_sc_hd__buf_2
Xoutput113 net113 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__buf_2
Xoutput124 net124 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_149_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08575__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12513__A datapath.multiplication_module.multiplier_i\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07783__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10382__A2 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07953_ datapath.rf.registers\[28\]\[11\] net929 net920 vssd1 vssd1 vccd1 vccd1 _02789_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08327__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06904_ net957 net921 vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__and2_2
X_07884_ datapath.rf.registers\[18\]\[13\] net725 net667 datapath.rf.registers\[15\]\[13\]
+ _02719_ vssd1 vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__a221o_1
XFILLER_29_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07535__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09623_ net360 _04457_ _04458_ net345 vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__a31oi_1
X_06835_ _01487_ _01515_ net1015 vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__a21boi_1
XFILLER_56_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout367_A net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09288__A0 _02467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09554_ _03770_ _04364_ _04369_ _04389_ vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__a211o_1
X_06766_ _01466_ _01568_ net1030 datapath.ru.latched_instruction\[30\] vssd1 vssd1
+ vccd1 vccd1 _01603_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_102_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_65_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06884__C _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08505_ _03328_ _03332_ _03336_ _03340_ vssd1 vssd1 vccd1 vccd1 _03341_ sky130_fd_sc_hd__or4_1
X_06697_ net1289 net1282 mmio.memload_or_instruction\[9\] vssd1 vssd1 vccd1 vccd1
+ _01536_ sky130_fd_sc_hd__nor3b_2
X_09485_ _04318_ _04320_ net373 vssd1 vssd1 vccd1 vccd1 _04321_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout155_X net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout534_A net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08436_ datapath.rf.registers\[13\]\[2\] net969 _01823_ vssd1 vssd1 vccd1 vccd1 _03272_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07996__B _01707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08367_ net874 _03197_ _03199_ _03202_ vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__or4_4
X_07318_ datapath.rf.registers\[9\]\[24\] net885 net877 datapath.rf.registers\[8\]\[24\]
+ _02153_ vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__a221o_1
XANTENNA__07066__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08298_ _03131_ _03133_ vssd1 vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__or2_1
XANTENNA__09460__B1 _04294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12407__B net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07249_ datapath.rf.registers\[17\]\[26\] net746 net738 datapath.rf.registers\[16\]\[26\]
+ _02084_ vssd1 vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__a221o_1
XFILLER_137_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1231_X net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10260_ _04857_ _04859_ vssd1 vssd1 vccd1 vccd1 _05096_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08460__X _03296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout691_X net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10358__C1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout789_X net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09763__A1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10191_ _04999_ _05026_ _05023_ net228 vssd1 vssd1 vccd1 vccd1 _05027_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_76_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09763__B2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07517__A net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout340 net343 vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__buf_2
XFILLER_94_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout956_X net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08318__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout351 _03650_ vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__buf_2
Xfanout362 net365 vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__buf_2
X_13950_ clknet_leaf_103_clk _00728_ net1225 vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__dfrtp_1
Xfanout373 _03625_ vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__buf_2
Xfanout384 net385 vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__buf_6
XFILLER_87_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout395 _06555_ vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__buf_4
X_12901_ net2455 net296 net482 vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__mux2_1
XFILLER_101_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13881_ clknet_leaf_72_clk _00685_ net1242 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[25\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11473__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12832_ net289 net2609 net489 vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ _05518_ _05691_ vssd1 vssd1 vccd1 vccd1 _06550_ sky130_fd_sc_hd__or2_4
XFILLER_15_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14502_ clknet_leaf_23_clk _01207_ net1154 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11714_ net31 net1033 net1023 net1496 vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__o22a_1
X_12694_ _06518_ _06524_ _06523_ _06522_ vssd1 vssd1 vccd1 vccd1 _06526_ sky130_fd_sc_hd__o211ai_1
X_14433_ clknet_leaf_46_clk _01138_ net1172 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11645_ _05788_ _05866_ _05868_ vssd1 vssd1 vccd1 vccd1 _05869_ sky130_fd_sc_hd__or3b_1
XFILLER_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput15 DAT_I[21] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
X_14364_ clknet_leaf_8_clk _01069_ net1071 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07057__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput26 DAT_I[31] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
X_11576_ net1278 net1279 vssd1 vssd1 vccd1 vccd1 _05800_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_96_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput37 gpio_in[7] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__buf_1
XFILLER_155_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13315_ clknet_leaf_121_clk _00125_ net1192 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08514__C _01825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10527_ screen.controlBus\[6\] _05316_ _05326_ screen.controlBus\[7\] vssd1 vssd1
+ vccd1 vccd1 _05357_ sky130_fd_sc_hd__or4b_1
X_14295_ clknet_leaf_124_clk _01000_ net1208 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10458_ _01405_ _05291_ _05290_ vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__a21bo_1
X_13246_ clknet_leaf_1_clk _00056_ net1056 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_124_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13177_ net2134 vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__clkbuf_1
X_10389_ _05223_ _05224_ _01607_ vssd1 vssd1 vccd1 vccd1 _05225_ sky130_fd_sc_hd__a21oi_1
XFILLER_112_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07765__B1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06969__C net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08863__A_N _03669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12128_ net1270 screen.counter.ct\[18\] _06164_ vssd1 vssd1 vccd1 vccd1 _06165_ sky130_fd_sc_hd__and3_1
XANTENNA__08309__A2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12059_ screen.register.currentYbus\[28\] _05757_ _05769_ screen.register.currentXbus\[20\]
+ vssd1 vssd1 vccd1 vccd1 _06100_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_127_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11891__B net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14418__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12479__S net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11383__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08190__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06620_ net1286 net1281 mmio.key_data\[3\] vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_36_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09270_ _04104_ _04105_ vssd1 vssd1 vccd1 vccd1 _04106_ sky130_fd_sc_hd__or2_1
XANTENNA__07296__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08221_ datapath.rf.registers\[0\]\[6\] net866 _03045_ _03056_ vssd1 vssd1 vccd1
+ vccd1 _03057_ sky130_fd_sc_hd__a2bb2o_4
XTAP_TAPCELL_ROW_60_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10727__S _05367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13103__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08152_ datapath.rf.registers\[10\]\[7\] net987 _01720_ vssd1 vssd1 vccd1 vccd1 _02988_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07048__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12041__A2 _05773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07103_ datapath.rf.registers\[8\]\[29\] net695 net665 datapath.rf.registers\[15\]\[29\]
+ _01936_ vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__a221o_1
XFILLER_9_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_3_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08083_ _02917_ _02918_ vssd1 vssd1 vccd1 vccd1 _02919_ sky130_fd_sc_hd__or2_1
XANTENNA__12942__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_9_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_8
X_07034_ datapath.rf.registers\[14\]\[30\] net830 net800 datapath.rf.registers\[15\]\[30\]
+ _01869_ vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__a221o_1
XFILLER_103_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07756__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07220__A2 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08985_ _03819_ _03820_ _03779_ _03799_ vssd1 vssd1 vccd1 vccd1 _03821_ sky130_fd_sc_hd__and4b_1
XANTENNA_fanout484_A net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07936_ net613 _02771_ net564 vssd1 vssd1 vccd1 vccd1 _02772_ sky130_fd_sc_hd__a21oi_2
XFILLER_29_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07867_ _02693_ _02697_ _02699_ _02702_ vssd1 vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__nor4_1
XFILLER_84_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11855__A2 _05073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11293__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08181__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09606_ net362 _04325_ _04441_ net373 vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__o211a_1
X_06818_ datapath.ru.latched_instruction\[16\] _01523_ net1014 vssd1 vssd1 vccd1 vccd1
+ _01654_ sky130_fd_sc_hd__mux2_2
X_07798_ _02633_ vssd1 vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__inv_2
XFILLER_25_920 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09537_ net366 _04370_ _04372_ vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__o21a_1
X_06749_ _01585_ _01587_ _01582_ _01583_ vssd1 vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__or4bb_2
XANTENNA__07503__C net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout537_X net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10815__A0 _04580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09468_ net552 net548 _03205_ vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__a21o_1
XFILLER_12_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07800__A _02613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08419_ datapath.rf.registers\[4\]\[2\] net865 _03236_ _03237_ _03241_ vssd1 vssd1
+ vccd1 vccd1 _03255_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout704_X net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09399_ _03523_ net623 _03524_ net906 vssd1 vssd1 vccd1 vccd1 _04235_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__13013__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11430_ net233 net2246 net514 vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__mux2_1
XFILLER_138_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09433__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10583__D _02771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11361_ net220 net2050 net518 vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__mux2_1
XFILLER_138_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12852__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10594__A2 _05416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14030__RESET_B net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13100_ net296 net1795 net470 vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__mux2_1
X_10312_ _04475_ _05147_ vssd1 vssd1 vccd1 vccd1 _05148_ sky130_fd_sc_hd__nand2_1
X_11292_ net218 net2365 net522 vssd1 vssd1 vccd1 vccd1 _00340_ sky130_fd_sc_hd__mux2_1
X_14080_ clknet_leaf_101_clk _00846_ net1227 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_138_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11468__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08539__A2 _01716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13031_ net287 net2402 net477 vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__mux2_1
X_10243_ net466 _04428_ vssd1 vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_91_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07747__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08350__B net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10174_ _03947_ _03949_ _01702_ vssd1 vssd1 vccd1 vccd1 _05010_ sky130_fd_sc_hd__a21oi_1
Xfanout1102 net1110 vssd1 vssd1 vccd1 vccd1 net1102 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07211__A2 _02045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1113 net1115 vssd1 vssd1 vccd1 vccd1 net1113 sky130_fd_sc_hd__clkbuf_4
XFILLER_79_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1124 net1126 vssd1 vssd1 vccd1 vccd1 net1124 sky130_fd_sc_hd__clkbuf_4
XFILLER_120_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1135 net1139 vssd1 vssd1 vccd1 vccd1 net1135 sky130_fd_sc_hd__clkbuf_4
Xfanout1146 net1148 vssd1 vssd1 vccd1 vccd1 net1146 sky130_fd_sc_hd__buf_2
XFILLER_93_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1157 net1162 vssd1 vssd1 vccd1 vccd1 net1157 sky130_fd_sc_hd__clkbuf_2
Xfanout170 net171 vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_109_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1168 net1170 vssd1 vssd1 vccd1 vccd1 net1168 sky130_fd_sc_hd__clkbuf_2
Xfanout1179 net1180 vssd1 vssd1 vccd1 vccd1 net1179 sky130_fd_sc_hd__clkbuf_4
Xfanout181 net182 vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__clkbuf_2
Xfanout192 _05659_ vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__clkbuf_2
X_13933_ clknet_leaf_110_clk _00711_ net1222 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_75_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13864_ clknet_leaf_72_clk _00668_ net1243 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_75_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_122_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12815_ net1677 net218 net490 vssd1 vssd1 vccd1 vccd1 _01067_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_122_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13795_ clknet_leaf_52_clk _00604_ net1184 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12746_ net1881 net248 net403 vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__mux2_1
XANTENNA__08806__A _03601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14189__RESET_B net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12677_ net499 _06510_ _06511_ net503 net2318 vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__a32o_1
XANTENNA__08525__B _03358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14416_ clknet_leaf_24_clk _01121_ net1157 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11628_ _05800_ _05806_ _05850_ vssd1 vssd1 vccd1 vccd1 _05852_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_100_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12762__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14347_ clknet_leaf_56_clk _01052_ net1171 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11559_ _05754_ _05774_ vssd1 vssd1 vccd1 vccd1 _05783_ sky130_fd_sc_hd__or2_2
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold607 datapath.rf.registers\[22\]\[0\] vssd1 vssd1 vccd1 vccd1 net1955 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07986__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire593 _01933_ vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__clkbuf_1
Xhold618 datapath.rf.registers\[1\]\[15\] vssd1 vssd1 vccd1 vccd1 net1966 sky130_fd_sc_hd__dlygate4sd3_1
Xhold629 datapath.rf.registers\[4\]\[9\] vssd1 vssd1 vccd1 vccd1 net1977 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14278_ clknet_leaf_11_clk _00983_ net1083 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11378__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13229_ clknet_leaf_131_clk _00039_ net1113 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07738__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07202__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1307 keypad.apps.app_c\[0\] vssd1 vssd1 vccd1 vccd1 net2655 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08770_ _01859_ _03481_ _03598_ vssd1 vssd1 vccd1 vccd1 _03606_ sky130_fd_sc_hd__or3_1
XFILLER_78_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07721_ net872 _02552_ _02554_ _02556_ vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__or4_2
XFILLER_66_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07652_ net613 _02487_ net565 vssd1 vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__a21o_1
XFILLER_81_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06603_ net1286 net1281 mmio.memload_or_instruction\[2\] vssd1 vssd1 vccd1 vccd1
+ _01442_ sky130_fd_sc_hd__or3_1
XFILLER_25_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07583_ datapath.rf.registers\[0\]\[19\] net868 _02417_ vssd1 vssd1 vccd1 vccd1 _02419_
+ sky130_fd_sc_hd__o21ai_4
XANTENNA__12937__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09322_ _02419_ _02467_ net453 vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__mux2_1
X_09253_ net557 net577 net546 _02419_ vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__o211a_1
XANTENNA__08772__C_N _03601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08435__B net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08204_ datapath.rf.registers\[4\]\[6\] net957 net931 vssd1 vssd1 vccd1 vccd1 _03040_
+ sky130_fd_sc_hd__and3_1
X_09184_ net337 _04019_ vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__nand2_1
XANTENNA__08154__C net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08135_ datapath.rf.registers\[17\]\[8\] net749 net725 datapath.rf.registers\[18\]\[8\]
+ _02970_ vssd1 vssd1 vccd1 vccd1 _02971_ sky130_fd_sc_hd__a221o_1
XFILLER_134_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07977__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08066_ datapath.rf.registers\[30\]\[9\] net834 net802 datapath.rf.registers\[3\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__a22o_1
XANTENNA__07441__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07993__C net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07017_ _01841_ _01844_ _01845_ _01852_ vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__or4_2
XANTENNA__11288__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout699_A net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07729__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08926__C1 _01889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09194__A2 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout866_A net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout487_X net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08968_ net560 net447 vssd1 vssd1 vccd1 vccd1 _03804_ sky130_fd_sc_hd__nor2_1
XANTENNA__07354__X _02190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07919_ datapath.rf.registers\[16\]\[12\] net741 net725 datapath.rf.registers\[18\]\[12\]
+ _02753_ vssd1 vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__a221o_1
XFILLER_84_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout654_X net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08899_ net1268 datapath.PC\[7\] _03734_ vssd1 vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__or3_1
XFILLER_84_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_3_Left_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13008__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10930_ datapath.PC\[29\] _05665_ vssd1 vssd1 vccd1 vccd1 _05671_ sky130_fd_sc_hd__and2_1
XFILLER_57_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10861_ datapath.PC\[18\] _05600_ datapath.PC\[19\] vssd1 vssd1 vccd1 vccd1 _05612_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout821_X net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12847__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09103__C1 _03673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout919_X net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12600_ datapath.mulitply_result\[15\] datapath.multiplication_module.multiplicand_i\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06447_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_27_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13580_ clknet_leaf_133_clk _00390_ net1111 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10792_ _01467_ net620 _05552_ _05553_ vssd1 vssd1 vccd1 vccd1 _05554_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__14282__RESET_B net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12531_ net2538 net504 net500 _06389_ vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__a22o_1
XFILLER_149_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08345__B net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14211__RESET_B net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12462_ net166 _05972_ net128 screen.register.currentXbus\[18\] vssd1 vssd1 vccd1
+ vccd1 _00864_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09406__B1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07680__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14201_ clknet_leaf_67_clk datapath.multiplication_module.multiplicand_i_n\[12\]
+ net1240 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11413_ net303 net1846 net516 vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__mux2_1
X_12393_ _05950_ net157 vssd1 vssd1 vccd1 vccd1 _06344_ sky130_fd_sc_hd__nor2_1
XANTENNA__07968__B1 _02803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11764__B2 _02189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14132_ clknet_leaf_33_clk _00889_ net1128 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07432__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11344_ net259 net2257 net520 vssd1 vssd1 vccd1 vccd1 _00387_ sky130_fd_sc_hd__mux2_1
XFILLER_126_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11198__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14063_ clknet_leaf_122_clk _00830_ net1200 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11275_ net261 net2633 net525 vssd1 vssd1 vccd1 vccd1 _00323_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_148_Right_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09744__X _04580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13014_ net1629 net236 net392 vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__mux2_1
X_10226_ _03822_ _03826_ _01702_ vssd1 vssd1 vccd1 vccd1 _05062_ sky130_fd_sc_hd__a21o_1
XANTENNA__07408__C net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10157_ _04992_ _04603_ net640 _04991_ vssd1 vssd1 vccd1 vccd1 _04993_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__10830__S net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold4 screen.screenEdge.enable1 vssd1 vssd1 vccd1 vccd1 net1352 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_121_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11819__A2 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10088_ datapath.PC\[25\] _01702_ net1043 vssd1 vssd1 vccd1 vccd1 _04924_ sky130_fd_sc_hd__a21o_1
XFILLER_75_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13916_ clknet_leaf_101_clk _00694_ net1227 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_63_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13847_ clknet_leaf_77_clk net1353 net1246 vssd1 vssd1 vccd1 vccd1 mmio.key_en2 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12757__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09645__B1 _03770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13778_ clknet_leaf_85_clk _00587_ net1258 vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__dfrtp_1
X_12729_ _05893_ _06548_ _06530_ vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__a21o_1
XANTENNA__07120__A1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11897__A _02725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12492__S net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_152_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11755__B2 _02634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold404 datapath.rf.registers\[23\]\[25\] vssd1 vssd1 vccd1 vccd1 net1752 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold415 datapath.rf.registers\[6\]\[31\] vssd1 vssd1 vccd1 vccd1 net1763 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07423__A2 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13885__Q datapath.ru.latched_instruction\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold426 datapath.rf.registers\[8\]\[2\] vssd1 vssd1 vccd1 vccd1 net1774 sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 datapath.rf.registers\[7\]\[17\] vssd1 vssd1 vccd1 vccd1 net1785 sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 datapath.rf.registers\[27\]\[24\] vssd1 vssd1 vccd1 vccd1 net1796 sky130_fd_sc_hd__dlygate4sd3_1
Xhold459 datapath.rf.registers\[0\]\[23\] vssd1 vssd1 vccd1 vccd1 net1807 sky130_fd_sc_hd__dlygate4sd3_1
X_09940_ datapath.PC\[3\] _03206_ vssd1 vssd1 vccd1 vccd1 _04776_ sky130_fd_sc_hd__and2_1
XFILLER_132_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout906 _01619_ vssd1 vssd1 vccd1 vccd1 net906 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_115_Right_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout917 _01764_ vssd1 vssd1 vccd1 vccd1 net917 sky130_fd_sc_hd__buf_4
X_09871_ net626 _04706_ vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__nand2_1
Xfanout928 _01732_ vssd1 vssd1 vccd1 vccd1 net928 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout939 _01718_ vssd1 vssd1 vccd1 vccd1 net939 sky130_fd_sc_hd__buf_4
X_08822_ net552 net548 vssd1 vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__nand2_1
Xhold1104 datapath.rf.registers\[2\]\[23\] vssd1 vssd1 vccd1 vccd1 net2452 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1115 datapath.rf.registers\[18\]\[22\] vssd1 vssd1 vccd1 vccd1 net2463 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07592__D1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1126 datapath.rf.registers\[18\]\[25\] vssd1 vssd1 vccd1 vccd1 net2474 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1137 datapath.rf.registers\[30\]\[22\] vssd1 vssd1 vccd1 vccd1 net2485 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08753_ _03497_ _03499_ _03588_ vssd1 vssd1 vccd1 vccd1 _03589_ sky130_fd_sc_hd__and3_1
Xhold1148 datapath.rf.registers\[3\]\[21\] vssd1 vssd1 vccd1 vccd1 net2496 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1159 screen.controlBus\[6\] vssd1 vssd1 vccd1 vccd1 net2507 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08136__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07704_ _02526_ _02527_ _02538_ _02539_ vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__or4_1
XFILLER_66_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08684_ _03519_ vssd1 vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__inv_2
XANTENNA__08149__C net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09830__A _01610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07635_ datapath.rf.registers\[27\]\[18\] net683 net660 datapath.rf.registers\[5\]\[18\]
+ _02470_ vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__a221o_1
XFILLER_54_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1091_A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1189_A net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07566_ datapath.rf.registers\[28\]\[19\] net929 net920 vssd1 vssd1 vccd1 vccd1 _02402_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_24_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09305_ _03515_ net626 net625 _03514_ net643 vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__a221oi_1
XFILLER_110_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10246__A1 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07497_ _02311_ _02332_ vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__and2_1
XFILLER_139_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09236_ _03775_ _04071_ net361 vssd1 vssd1 vccd1 vccd1 _04072_ sky130_fd_sc_hd__mux2_1
XFILLER_155_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_30_clk_X clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12255__X _06246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout402_X net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09167_ net575 _04001_ _04002_ _03990_ vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__a22o_1
XFILLER_107_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11746__B2 _03076_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08118_ datapath.rf.registers\[4\]\[8\] net864 net816 datapath.rf.registers\[21\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02954_ sky130_fd_sc_hd__a22o_1
XFILLER_119_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07414__A2 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09098_ net649 _03933_ net438 vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout983_A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08049_ datapath.rf.registers\[11\]\[9\] net986 net938 vssd1 vssd1 vccd1 vccd1 _02885_
+ sky130_fd_sc_hd__and3_1
XFILLER_123_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold960 datapath.rf.registers\[1\]\[19\] vssd1 vssd1 vccd1 vccd1 net2308 sky130_fd_sc_hd__dlygate4sd3_1
Xhold971 mmio.key_data\[6\] vssd1 vssd1 vccd1 vccd1 net2319 sky130_fd_sc_hd__dlygate4sd3_1
Xhold982 datapath.rf.registers\[25\]\[14\] vssd1 vssd1 vccd1 vccd1 net2330 sky130_fd_sc_hd__dlygate4sd3_1
X_11060_ net211 net2171 net430 vssd1 vssd1 vccd1 vccd1 _00120_ sky130_fd_sc_hd__mux2_1
Xhold993 datapath.rf.registers\[19\]\[29\] vssd1 vssd1 vccd1 vccd1 net2341 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout771_X net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08375__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10011_ _04794_ _04796_ vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__xnor2_1
XFILLER_131_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_48_Left_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08127__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10589__C _01954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11962_ _05999_ _06007_ vssd1 vssd1 vccd1 vccd1 _06008_ sky130_fd_sc_hd__or2_1
XFILLER_151_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13701_ clknet_leaf_115_clk _00511_ net1188 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_86_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09740__A net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08059__C net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10913_ _04624_ _05656_ net901 vssd1 vssd1 vccd1 vccd1 _05657_ sky130_fd_sc_hd__mux2_2
X_14681_ clknet_leaf_31_clk _01386_ net1122 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_11893_ net2476 net160 vssd1 vssd1 vccd1 vccd1 _05959_ sky130_fd_sc_hd__nand2_1
XFILLER_60_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11481__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13632_ clknet_leaf_134_clk _00442_ net1112 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10844_ datapath.mulitply_result\[16\] net615 net653 vssd1 vssd1 vccd1 vccd1 _05598_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_4_11_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13563_ clknet_leaf_45_clk _00373_ net1146 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10775_ net901 _04474_ _05538_ vssd1 vssd1 vccd1 vccd1 _05539_ sky130_fd_sc_hd__o21ai_2
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09739__X _04575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12514_ datapath.multiplication_module.multiplier_i\[0\] _05368_ vssd1 vssd1 vccd1
+ vccd1 _06375_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_57_Left_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10892__Y _05639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13494_ clknet_leaf_139_clk _00304_ net1099 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_12445_ net167 _05938_ net129 net2585 vssd1 vssd1 vccd1 vccd1 _00847_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_117_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12376_ net1363 _01428_ _06334_ screen.counter.currentEnable vssd1 vssd1 vccd1 vccd1
+ _00813_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_10_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14115_ clknet_leaf_75_clk net622 net1246 vssd1 vssd1 vccd1 vccd1 datapath.ru.n_memread
+ sky130_fd_sc_hd__dfrtp_1
X_11327_ net1689 net219 net414 vssd1 vssd1 vccd1 vccd1 _00372_ sky130_fd_sc_hd__mux2_1
XFILLER_114_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14046_ clknet_leaf_99_clk net1350 net1229 vssd1 vssd1 vccd1 vccd1 screen.register.xFill2
+ sky130_fd_sc_hd__dfrtp_1
X_11258_ net240 net1911 net420 vssd1 vssd1 vccd1 vccd1 _00307_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10209_ net1041 _05042_ _05044_ net640 vssd1 vssd1 vccd1 vccd1 _05045_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_66_Left_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11189_ net248 net2252 net423 vssd1 vssd1 vccd1 vccd1 _00241_ sky130_fd_sc_hd__mux2_1
XFILLER_94_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08118__B1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09315__C1 _02466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08965__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11673__B1 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12487__S net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11391__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06993__B _01823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07420_ datapath.rf.registers\[14\]\[22\] net829 net796 datapath.rf.registers\[29\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__a22o_1
XFILLER_23_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07351_ datapath.rf.registers\[3\]\[24\] net771 net763 datapath.rf.registers\[1\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_75_Left_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07282_ datapath.rf.registers\[5\]\[25\] net820 _02101_ _02103_ _02105_ vssd1 vssd1
+ vccd1 vccd1 _02118_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07644__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08841__A1 _03296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09021_ _03856_ vssd1 vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__inv_2
XANTENNA__13111__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09097__A net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold201 datapath.multiplication_module.multiplicand_i\[22\] vssd1 vssd1 vccd1 vccd1
+ net1549 sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 datapath.rf.registers\[11\]\[24\] vssd1 vssd1 vccd1 vccd1 net1560 sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 datapath.rf.registers\[5\]\[23\] vssd1 vssd1 vccd1 vccd1 net1571 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08432__C _01816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold234 datapath.rf.registers\[16\]\[28\] vssd1 vssd1 vccd1 vccd1 net1582 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12950__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold245 datapath.rf.registers\[2\]\[17\] vssd1 vssd1 vccd1 vccd1 net1593 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold256 datapath.rf.registers\[13\]\[2\] vssd1 vssd1 vccd1 vccd1 net1604 sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 datapath.rf.registers\[7\]\[21\] vssd1 vssd1 vccd1 vccd1 net1615 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold278 datapath.rf.registers\[5\]\[12\] vssd1 vssd1 vccd1 vccd1 net1626 sky130_fd_sc_hd__dlygate4sd3_1
X_09923_ _04758_ vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__inv_2
Xhold289 datapath.rf.registers\[14\]\[18\] vssd1 vssd1 vccd1 vccd1 net1637 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout703 net705 vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__buf_4
Xfanout714 net717 vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_84_Left_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06801__X _01637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08357__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout725 _01813_ vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout397_A _06555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout736 net737 vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__clkbuf_8
Xfanout747 net749 vssd1 vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__buf_2
X_09854_ _02242_ _02285_ _04688_ _04689_ _02241_ vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__o2111a_1
Xfanout758 _01802_ vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__clkbuf_8
XFILLER_113_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1104_A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout769 _01799_ vssd1 vssd1 vccd1 vccd1 net769 sky130_fd_sc_hd__clkbuf_4
X_08805_ _03637_ _03640_ vssd1 vssd1 vccd1 vccd1 _03641_ sky130_fd_sc_hd__and2_2
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09785_ net905 _03492_ _03700_ _04555_ _04620_ vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__a221o_1
X_06997_ datapath.rf.registers\[7\]\[31\] net671 net669 datapath.rf.registers\[21\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__a22o_1
XANTENNA__08109__B1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout564_A _01786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08736_ _03530_ _03531_ _03570_ _03527_ vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__a31o_1
XFILLER_26_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_72_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout731_A _01811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08667_ _02312_ _02332_ vssd1 vssd1 vccd1 vccd1 _03503_ sky130_fd_sc_hd__nor2_1
XANTENNA__07999__B net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout829_A net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07618_ datapath.rf.registers\[5\]\[18\] net819 _02445_ _02446_ _02448_ vssd1 vssd1
+ vccd1 vccd1 _02454_ sky130_fd_sc_hd__a2111o_1
XFILLER_81_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07883__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_93_Left_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08598_ _03433_ vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__inv_2
X_07549_ datapath.rf.registers\[0\]\[20\] net783 _02384_ vssd1 vssd1 vccd1 vccd1 _02385_
+ sky130_fd_sc_hd__o21a_4
XANTENNA_fanout1261_X net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_87_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10560_ screen.register.currentXbus\[17\] screen.register.currentXbus\[16\] screen.register.currentXbus\[19\]
+ screen.register.currentXbus\[18\] vssd1 vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__or4_1
XANTENNA__07635__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08832__A1 _03661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13856__RESET_B net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_130_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09219_ _04046_ _04050_ _04054_ vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__and3_1
XFILLER_148_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10491_ _05319_ _05320_ vssd1 vssd1 vccd1 vccd1 _05321_ sky130_fd_sc_hd__or2_1
XFILLER_154_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13021__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12230_ screen.counter.currentCt\[14\] _06228_ net602 vssd1 vssd1 vccd1 vccd1 _06230_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_leaf_10_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout986_X net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08342__C net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10591__D _02385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12161_ _06161_ _06172_ net1275 vssd1 vssd1 vccd1 vccd1 _06188_ sky130_fd_sc_hd__a21o_1
XANTENNA__12860__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_145_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11112_ net294 net2026 net426 vssd1 vssd1 vccd1 vccd1 _00167_ sky130_fd_sc_hd__mux2_1
XFILLER_150_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12092_ net1001 _06128_ _06130_ net1011 vssd1 vssd1 vccd1 vccd1 _06131_ sky130_fd_sc_hd__a22o_1
XFILLER_104_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold790 datapath.rf.registers\[13\]\[14\] vssd1 vssd1 vccd1 vccd1 net2138 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_25_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11043_ net297 net2644 net431 vssd1 vssd1 vccd1 vccd1 _00103_ sky130_fd_sc_hd__mux2_1
XANTENNA__07020__B1 _01787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_3_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_3_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_92_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12994_ _05696_ _05727_ vssd1 vssd1 vccd1 vccd1 _06557_ sky130_fd_sc_hd__nor2_1
XFILLER_45_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11945_ _01954_ net656 vssd1 vssd1 vccd1 vccd1 _05994_ sky130_fd_sc_hd__nand2_1
XFILLER_91_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14664_ clknet_leaf_65_clk _01369_ net1235 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11876_ _03076_ net656 vssd1 vssd1 vccd1 vccd1 _05948_ sky130_fd_sc_hd__nand2_1
XANTENNA__07874__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13615_ clknet_leaf_26_clk _00425_ net1135 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10827_ datapath.PC\[14\] _05576_ vssd1 vssd1 vccd1 vccd1 _05583_ sky130_fd_sc_hd__and2_1
XANTENNA__09076__A1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14595_ clknet_leaf_139_clk _01300_ net1099 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_119_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07087__B1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13546_ clknet_leaf_61_clk _00356_ net1164 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07626__A2 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10758_ net1269 datapath.PC\[3\] datapath.PC\[4\] vssd1 vssd1 vccd1 vccd1 _05524_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08833__C_N _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13477_ clknet_leaf_117_clk _00287_ net1190 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10689_ _05462_ _05482_ _05505_ _05428_ _01430_ vssd1 vssd1 vccd1 vccd1 _05506_ sky130_fd_sc_hd__o221a_1
XANTENNA__12336__A net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12428_ net1447 net132 _06361_ vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__a21o_1
XANTENNA__09784__C1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12770__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12359_ net229 _05673_ vssd1 vssd1 vccd1 vccd1 _06323_ sky130_fd_sc_hd__nand2_1
XFILLER_113_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11894__B net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06988__B _01823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11386__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14029_ clknet_leaf_82_clk _00798_ net1257 vssd1 vssd1 vccd1 vccd1 datapath.PC\[19\]
+ sky130_fd_sc_hd__dfrtp_2
X_06920_ net946 net932 vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__and2_2
XFILLER_68_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10290__S net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_842 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10697__A1 _03292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06851_ _01408_ _01582_ _01598_ datapath.ru.latched_instruction\[27\] vssd1 vssd1
+ vccd1 vccd1 _01687_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09570_ _04228_ _04370_ net366 vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__mux2_1
XANTENNA__12438__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06782_ _01614_ _01618_ vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__and2_1
XANTENNA__08548__X _03384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08521_ datapath.rf.registers\[0\]\[1\] net783 _03341_ _03356_ vssd1 vssd1 vccd1
+ vccd1 _03357_ sky130_fd_sc_hd__o22a_4
XFILLER_82_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08708__B _03228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08511__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13106__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07612__B net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08452_ datapath.rf.registers\[12\]\[2\] net757 net701 datapath.rf.registers\[23\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__a22o_1
XANTENNA__07865__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07403_ net465 vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__inv_2
XANTENNA__12945__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08383_ datapath.rf.registers\[11\]\[3\] net713 net709 datapath.rf.registers\[10\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03219_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout145_A net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07334_ datapath.rf.registers\[0\]\[24\] net871 _02159_ _02168_ vssd1 vssd1 vccd1
+ vccd1 _02170_ sky130_fd_sc_hd__o22ai_4
XTAP_TAPCELL_ROW_63_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07617__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08724__A _03057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07265_ datapath.rf.registers\[20\]\[25\] net959 net924 vssd1 vssd1 vccd1 vccd1 _02101_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1054_A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09004_ _01888_ net553 net549 vssd1 vssd1 vccd1 vccd1 _03840_ sky130_fd_sc_hd__or3_1
X_07196_ datapath.rf.registers\[4\]\[27\] net715 net702 datapath.rf.registers\[9\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02032_ sky130_fd_sc_hd__a22o_1
XFILLER_151_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1221_A net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07250__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout681_A _01828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout500 net501 vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__buf_2
Xfanout511 _05735_ vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11296__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout779_A _01794_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09906_ net604 _04741_ datapath.PC\[15\] vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__o21a_1
Xfanout522 _05723_ vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__buf_6
Xfanout533 _05718_ vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__clkbuf_4
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout544 net545 vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__buf_4
XFILLER_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout555 _03609_ vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07002__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout566 _01779_ vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07075__A _01889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout577 _03616_ vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__dlymetal6s2s_1
X_09837_ _03524_ _03530_ _04179_ _04240_ vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__or4bb_1
Xfanout599 net600 vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout946_A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09768_ _04023_ _04057_ _04603_ vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__or3_2
XANTENNA__08458__X _03294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08719_ _03552_ _03553_ _03544_ vssd1 vssd1 vccd1 vccd1 _03555_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout734_X net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ _04529_ _04531_ _04532_ _04533_ net609 vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__a32o_1
XANTENNA__13016__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11730_ net17 net1033 net1023 net1532 vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__o22a_1
XANTENNA__07856__A2 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10586__D _03417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11661_ button\[4\] _05874_ vssd1 vssd1 vccd1 vccd1 _05880_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout901_X net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12855__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13400_ clknet_leaf_7_clk _00210_ net1070 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10612_ button\[0\] net1022 vssd1 vssd1 vccd1 vccd1 _05432_ sky130_fd_sc_hd__nand2_1
X_14380_ clknet_leaf_18_clk _01085_ net1108 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11592_ net1280 screen.counter.ct\[5\] net1279 net1278 vssd1 vssd1 vccd1 vccd1 _05816_
+ sky130_fd_sc_hd__or4b_1
XFILLER_128_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13331_ clknet_leaf_33_clk _00141_ net1128 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10543_ datapath.multiplication_module.multiplier_i\[9\] datapath.multiplication_module.multiplier_i\[8\]
+ datapath.multiplication_module.multiplier_i\[11\] datapath.multiplication_module.multiplier_i\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05371_ sky130_fd_sc_hd__or4_1
XANTENNA__08281__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08353__B net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13262_ clknet_leaf_3_clk _00072_ net1076 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10474_ _05303_ vssd1 vssd1 vccd1 vccd1 _05304_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_114_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12213_ screen.counter.currentCt\[8\] _06217_ vssd1 vssd1 vccd1 vccd1 _06219_ sky130_fd_sc_hd__and2_1
XANTENNA__12365__B2 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12443__X _06369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13193_ datapath.rf.registers\[0\]\[30\] vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08033__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10376__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07241__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12144_ _05780_ _06171_ vssd1 vssd1 vccd1 vccd1 _06177_ sky130_fd_sc_hd__nor2_1
XFILLER_2_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09465__A _03423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12075_ _06076_ _06113_ _06114_ vssd1 vssd1 vccd1 vccd1 _06115_ sky130_fd_sc_hd__or3_1
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11026_ net210 net2106 net538 vssd1 vssd1 vccd1 vccd1 _00088_ sky130_fd_sc_hd__mux2_1
XANTENNA__08368__X _03204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08809__A _01647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12977_ net250 net1729 net479 vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_125_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11928_ net135 _05982_ _05981_ vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__o21ai_1
XFILLER_32_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08247__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14647_ clknet_leaf_126_clk _01352_ net1206 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11859_ net137 _05936_ _05935_ vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12765__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11522__X _05747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_18 clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14578_ clknet_leaf_32_clk _01283_ net1122 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11800__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13529_ clknet_leaf_31_clk _00339_ net1122 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08272__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07050_ _01882_ _01883_ _01884_ _01885_ vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__nor4_1
XANTENNA__07480__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08831__X _03667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 DAT_O[8] sky130_fd_sc_hd__buf_2
Xoutput114 net114 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__buf_2
XANTENNA__08024__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09221__A1 _01706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput125 net125 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__buf_2
XANTENNA__09221__B2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06999__A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07447__X _02283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_775 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07952_ datapath.rf.registers\[15\]\[11\] net985 net915 vssd1 vssd1 vccd1 vccd1 _02788_
+ sky130_fd_sc_hd__and3_1
XFILLER_96_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06903_ _01630_ _01638_ net979 vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__and3_2
X_07883_ datapath.rf.registers\[17\]\[13\] net749 net690 datapath.rf.registers\[31\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02719_ sky130_fd_sc_hd__a22o_1
X_09622_ net457 _04340_ _04343_ net351 vssd1 vssd1 vccd1 vccd1 _04458_ sky130_fd_sc_hd__a211o_1
XFILLER_95_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06834_ datapath.ru.n_memwrite2 datapath.ru.n_memread2 vssd1 vssd1 vccd1 vccd1 _01670_
+ sky130_fd_sc_hd__nor2_1
X_09553_ _03619_ _04388_ _04383_ _03613_ vssd1 vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_39_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09288__A1 _02523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06765_ datapath.ru.latched_instruction\[30\] net1029 _01568_ _01466_ vssd1 vssd1
+ vccd1 vccd1 _01602_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout262_A _05575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08438__B net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08504_ datapath.rf.registers\[9\]\[1\] net705 _03337_ _03338_ _03339_ vssd1 vssd1
+ vccd1 vccd1 _03340_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07299__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06884__D _01656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07838__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09484_ _02961_ net440 _04319_ net362 vssd1 vssd1 vccd1 vccd1 _04320_ sky130_fd_sc_hd__a211o_1
X_06696_ datapath.ru.latched_instruction\[28\] net1045 vssd1 vssd1 vccd1 vccd1 _01535_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_51_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08435_ datapath.rf.registers\[3\]\[2\] net914 _01797_ vssd1 vssd1 vccd1 vccd1 _03271_
+ sky130_fd_sc_hd__and3_1
XFILLER_24_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1171_A net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout527_A _05721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09187__A1_N net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12044__B1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08366_ _03185_ _03192_ _03200_ _03201_ vssd1 vssd1 vccd1 vccd1 _03202_ sky130_fd_sc_hd__or4_1
XANTENNA__07996__C net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07317_ datapath.rf.registers\[11\]\[24\] net983 net939 vssd1 vssd1 vccd1 vccd1 _02153_
+ sky130_fd_sc_hd__and3_1
XFILLER_109_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08263__A2 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08297_ datapath.rf.registers\[9\]\[4\] net886 net846 datapath.rf.registers\[1\]\[4\]
+ _03132_ vssd1 vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__a221o_1
XANTENNA__09460__A1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07471__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07248_ datapath.rf.registers\[27\]\[26\] net683 _02083_ net786 vssd1 vssd1 vccd1
+ vccd1 _02084_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_12_Left_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08015__A2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07179_ datapath.rf.registers\[5\]\[27\] net819 net813 datapath.rf.registers\[23\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__a22o_1
XFILLER_118_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10190_ _05021_ _05025_ _05024_ vssd1 vssd1 vccd1 vccd1 _05026_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_76_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout684_X net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout330 _03619_ vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__buf_2
Xfanout341 net343 vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08665__A_N net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout352 _03650_ vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__clkbuf_2
Xfanout363 net365 vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout851_X net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout374 _03625_ vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__buf_2
XANTENNA_fanout949_X net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout385 _06562_ vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__clkbuf_4
X_12900_ net1713 net298 net482 vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__mux2_1
Xfanout396 _06555_ vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__clkbuf_8
X_13880_ clknet_leaf_53_clk _00684_ net1183 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_21_Left_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12831_ net260 net1818 net489 vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__mux2_1
XANTENNA__09279__A1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08348__B net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12762_ net2589 net168 net403 vssd1 vssd1 vccd1 vccd1 _00984_ sky130_fd_sc_hd__mux2_1
XANTENNA__07829__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14501_ clknet_leaf_116_clk _01206_ net1187 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11713_ net30 net1033 net1023 net1377 vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__o22a_1
XFILLER_15_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12693_ _06522_ _06523_ _06524_ _06518_ vssd1 vssd1 vccd1 vccd1 _06525_ sky130_fd_sc_hd__a211o_1
XFILLER_14_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14432_ clknet_leaf_132_clk _01137_ net1112 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_11644_ _05349_ net998 _05824_ vssd1 vssd1 vccd1 vccd1 _05868_ sky130_fd_sc_hd__nor3_1
XANTENNA__12035__B1 _06018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14363_ clknet_leaf_37_clk _01068_ net1136 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput16 DAT_I[22] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
X_11575_ _05798_ vssd1 vssd1 vccd1 vccd1 _05799_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_30_Left_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08254__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput27 DAT_I[3] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_96_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput38 gpio_in[8] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__buf_1
X_13314_ clknet_leaf_151_clk _00124_ net1052 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_96_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10526_ screen.counter.ct\[1\] net1278 _05355_ _05354_ vssd1 vssd1 vccd1 vccd1 _05356_
+ sky130_fd_sc_hd__a31o_1
XFILLER_6_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14294_ clknet_leaf_139_clk _00999_ net1099 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13394__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13245_ clknet_leaf_136_clk _00055_ net1091 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10457_ _04909_ _05073_ _05285_ _05286_ mmio.wishbone.curr_state\[0\] vssd1 vssd1
+ vccd1 vccd1 _05291_ sky130_fd_sc_hd__o311a_2
XANTENNA__10833__S net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07214__B1 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07708__A _02522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13176_ net1512 vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__clkbuf_1
X_10388_ _01610_ _05215_ _05217_ vssd1 vssd1 vccd1 vccd1 _05224_ sky130_fd_sc_hd__a21oi_1
X_12127_ net1273 _06153_ _06163_ vssd1 vssd1 vccd1 vccd1 _06164_ sky130_fd_sc_hd__and3_1
XFILLER_97_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12058_ _06095_ _06096_ _06097_ _06098_ vssd1 vssd1 vccd1 vccd1 _06099_ sky130_fd_sc_hd__or4_1
XFILLER_77_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12510__A1 datapath.multiplication_module.multiplier_i\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11009_ net294 net1984 net539 vssd1 vssd1 vccd1 vccd1 _00071_ sky130_fd_sc_hd__mux2_1
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08098__X _02934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10285__C1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12495__S net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08220_ _03047_ _03051_ _03053_ _03055_ vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__nor4_1
XANTENNA__13180__A datapath.rf.registers\[0\]\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08151_ datapath.rf.registers\[3\]\[7\] net803 vssd1 vssd1 vccd1 vccd1 _02987_ sky130_fd_sc_hd__nand2_1
XFILLER_146_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07102_ datapath.rf.registers\[14\]\[29\] net775 net711 datapath.rf.registers\[11\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_155_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08082_ datapath.rf.registers\[1\]\[9\] net764 net720 datapath.rf.registers\[20\]\[9\]
+ _02916_ vssd1 vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__a221o_1
X_07033_ datapath.rf.registers\[20\]\[30\] net959 net925 vssd1 vssd1 vccd1 vccd1 _01869_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_58_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08953__A0 _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08984_ net905 _03487_ net318 _03818_ vssd1 vssd1 vccd1 vccd1 _03820_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_114_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07935_ datapath.rf.registers\[0\]\[12\] net783 _02760_ _02770_ vssd1 vssd1 vccd1
+ vccd1 _02771_ sky130_fd_sc_hd__o22a_4
X_07866_ _02685_ _02687_ _02700_ _02701_ vssd1 vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__or4_1
X_09605_ _02961_ net440 _04319_ net366 vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__a211o_1
X_06817_ _01411_ _01575_ _01573_ vssd1 vssd1 vccd1 vccd1 _01653_ sky130_fd_sc_hd__o21a_1
XFILLER_56_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07797_ datapath.rf.registers\[0\]\[15\] net784 _02618_ _02632_ vssd1 vssd1 vccd1
+ vccd1 _02633_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_73_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09536_ _02805_ net440 _04371_ net362 vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__a211o_1
X_06748_ _01443_ net1005 net1021 net1029 datapath.ru.latched_instruction\[2\] vssd1
+ vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__a32o_1
XANTENNA__12265__B1 _06253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10276__C1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09467_ net560 net464 net452 vssd1 vssd1 vccd1 vccd1 _04303_ sky130_fd_sc_hd__mux2_1
X_06679_ datapath.ru.latched_instruction\[26\] _01504_ _01513_ datapath.ru.latched_instruction\[14\]
+ vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout811_A net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout432_X net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12017__B1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08418_ datapath.rf.registers\[21\]\[2\] net816 _03238_ _03239_ _03240_ vssd1 vssd1
+ vccd1 vccd1 _03254_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07692__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09398_ net574 _04223_ _04224_ _04233_ vssd1 vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_138_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08349_ datapath.rf.registers\[21\]\[3\] net948 _01739_ vssd1 vssd1 vccd1 vccd1 _03185_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08236__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_129_Right_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07444__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11360_ net239 net2348 net520 vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__mux2_1
XFILLER_138_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout899_X net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10311_ _04429_ _04455_ _04474_ vssd1 vssd1 vccd1 vccd1 _05147_ sky130_fd_sc_hd__a21o_1
XFILLER_152_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11291_ net239 net2380 net524 vssd1 vssd1 vccd1 vccd1 _00339_ sky130_fd_sc_hd__mux2_1
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13030_ net258 net2089 net476 vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__mux2_1
X_10242_ _04429_ _05077_ vssd1 vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08944__A0 _02169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08350__C _01744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10173_ _04977_ _04987_ _04997_ _05008_ vssd1 vssd1 vccd1 vccd1 _05009_ sky130_fd_sc_hd__or4_1
Xfanout1103 net1110 vssd1 vssd1 vccd1 vccd1 net1103 sky130_fd_sc_hd__buf_2
Xfanout1114 net1115 vssd1 vssd1 vccd1 vccd1 net1114 sky130_fd_sc_hd__clkbuf_2
XFILLER_121_756 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1125 net1126 vssd1 vssd1 vccd1 vccd1 net1125 sky130_fd_sc_hd__clkbuf_2
Xfanout1136 net1139 vssd1 vssd1 vccd1 vccd1 net1136 sky130_fd_sc_hd__buf_2
XANTENNA_input38_A gpio_in[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1147 net1148 vssd1 vssd1 vccd1 vccd1 net1147 sky130_fd_sc_hd__clkbuf_4
Xfanout160 net161 vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__buf_2
Xfanout1158 net1162 vssd1 vssd1 vccd1 vccd1 net1158 sky130_fd_sc_hd__clkbuf_4
Xfanout171 _05688_ vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__buf_1
XANTENNA__11484__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1169 net1170 vssd1 vssd1 vccd1 vccd1 net1169 sky130_fd_sc_hd__clkbuf_4
Xfanout182 net184 vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__clkbuf_2
Xfanout193 _05659_ vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__buf_1
X_13932_ clknet_leaf_122_clk _00710_ net1201 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_86_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08172__B2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13863_ clknet_leaf_71_clk _00667_ net1244 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_89_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12814_ net2228 net240 net492 vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_122_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13794_ clknet_leaf_52_clk _00603_ net1183 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12745_ net2398 net252 net402 vssd1 vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__mux2_1
XANTENNA__08475__A2 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07710__B net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12676_ _06508_ _06509_ _06507_ vssd1 vssd1 vccd1 vccd1 _06511_ sky130_fd_sc_hd__o21ai_1
X_14415_ clknet_leaf_28_clk _01120_ net1134 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11627_ _05800_ _05806_ _05850_ vssd1 vssd1 vccd1 vccd1 _05851_ sky130_fd_sc_hd__nor3_1
XANTENNA__08227__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07435__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14346_ clknet_leaf_58_clk _01051_ net1167 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09918__A _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11558_ _05779_ _05781_ vssd1 vssd1 vccd1 vccd1 _05782_ sky130_fd_sc_hd__or2_1
Xwire561 _02568_ vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__buf_4
Xhold608 datapath.rf.registers\[5\]\[17\] vssd1 vssd1 vccd1 vccd1 net1956 sky130_fd_sc_hd__dlygate4sd3_1
Xwire583 _03001_ vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__buf_1
X_10509_ screen.counter.ct\[2\] _01425_ net1276 vssd1 vssd1 vccd1 vccd1 _05339_ sky130_fd_sc_hd__a21o_1
X_14277_ clknet_leaf_116_clk _00982_ net1189 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold619 datapath.rf.registers\[30\]\[15\] vssd1 vssd1 vccd1 vccd1 net1967 sky130_fd_sc_hd__dlygate4sd3_1
X_11489_ net268 net1638 net512 vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__mux2_1
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13228_ clknet_leaf_134_clk _00038_ net1105 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13159_ net1763 net170 net382 vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__mux2_1
XFILLER_33_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1308 screen.register.currentXbus\[10\] vssd1 vssd1 vccd1 vccd1 net2656 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11394__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06996__B _01831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07720_ datapath.rf.registers\[24\]\[16\] net856 net799 datapath.rf.registers\[15\]\[16\]
+ _02555_ vssd1 vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__a221o_1
XANTENNA__10151__X _04987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07651_ datapath.rf.registers\[0\]\[18\] net782 _02486_ vssd1 vssd1 vccd1 vccd1 _02487_
+ sky130_fd_sc_hd__o21a_4
XTAP_TAPCELL_ROW_0_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06602_ mmio.memload_or_instruction\[5\] net1049 _01440_ vssd1 vssd1 vccd1 vccd1
+ _01441_ sky130_fd_sc_hd__a21o_2
X_07582_ datapath.rf.registers\[0\]\[19\] net868 _02417_ vssd1 vssd1 vccd1 vccd1 _02418_
+ sky130_fd_sc_hd__o21a_2
X_09321_ net330 _04156_ net311 vssd1 vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__a21o_1
XANTENNA__13114__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10273__A2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09252_ net607 _04086_ vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__or2_1
XANTENNA__07674__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08203_ datapath.rf.registers\[18\]\[6\] net974 net949 vssd1 vssd1 vccd1 vccd1 _03039_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08435__C _01797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08218__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09183_ _04016_ _04018_ net340 vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__mux2_1
XANTENNA__12953__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout225_A net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07426__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08134_ datapath.rf.registers\[27\]\[8\] net686 _02968_ _02969_ net789 vssd1 vssd1
+ vccd1 vccd1 _02970_ sky130_fd_sc_hd__a2111o_1
XFILLER_119_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08065_ net874 _02898_ _02899_ _02900_ vssd1 vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout1134_A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07016_ _01847_ _01849_ _01851_ vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__or3_1
XFILLER_115_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout594_A net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08926__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08967_ _02960_ _03008_ net447 vssd1 vssd1 vccd1 vccd1 _03803_ sky130_fd_sc_hd__mux2_1
XFILLER_124_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout382_X net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout761_A _01802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07918_ datapath.rf.registers\[20\]\[12\] net719 net703 datapath.rf.registers\[9\]\[12\]
+ _02752_ vssd1 vssd1 vccd1 vccd1 _02754_ sky130_fd_sc_hd__a221o_1
X_08898_ datapath.PC\[5\] _03733_ vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__or2_1
XFILLER_68_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07849_ datapath.rf.registers\[26\]\[13\] net837 net805 datapath.rf.registers\[28\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02685_ sky130_fd_sc_hd__a22o_1
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout647_X net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10860_ datapath.PC\[18\] datapath.PC\[19\] _05600_ vssd1 vssd1 vccd1 vccd1 _05611_
+ sky130_fd_sc_hd__and3_1
XFILLER_72_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09519_ net354 _04217_ _04354_ vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__o21a_1
XFILLER_140_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout814_X net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10791_ datapath.mulitply_result\[8\] net598 net620 vssd1 vssd1 vccd1 vccd1 _05553_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__13024__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12530_ _06387_ _06388_ vssd1 vssd1 vccd1 vccd1 _06389_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08345__C net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12461_ net166 _05970_ net128 screen.register.currentXbus\[17\] vssd1 vssd1 vccd1
+ vccd1 _00863_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08209__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12863__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14200_ clknet_leaf_66_clk datapath.multiplication_module.multiplicand_i_n\[11\]
+ net1236 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11412_ net288 net1701 net517 vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__mux2_1
XANTENNA__07417__B1 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12392_ net2507 net133 _06343_ vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__a21o_1
XFILLER_153_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11479__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14131_ clknet_leaf_30_clk _00888_ net1124 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11343_ net208 net1823 net520 vssd1 vssd1 vccd1 vccd1 _00386_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_104_Left_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08090__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07529__Y _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14062_ clknet_leaf_121_clk _00829_ net1200 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07258__A _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11274_ net209 net2167 net525 vssd1 vssd1 vccd1 vccd1 _00322_ sky130_fd_sc_hd__mux2_1
X_13013_ net1643 net218 net391 vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__mux2_1
XFILLER_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10225_ datapath.PC\[29\] net1293 _05058_ _05060_ vssd1 vssd1 vccd1 vccd1 _05061_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07196__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10156_ _04084_ _04602_ net894 vssd1 vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06943__A2 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold5 mmio.key_en1 vssd1 vssd1 vccd1 vccd1 net1353 sky130_fd_sc_hd__dlygate4sd3_1
X_10087_ net641 _03915_ _04606_ vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__and3_1
XANTENNA__10412__A net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13915_ clknet_leaf_104_clk _00693_ net1225 vssd1 vssd1 vccd1 vccd1 screen.csx sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_113_Left_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10131__B net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload3_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13846_ clknet_leaf_78_clk net1351 net1245 vssd1 vssd1 vccd1 vccd1 mmio.WEN2 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07721__A net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09645__A1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08448__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13777_ clknet_leaf_85_clk _00586_ net1258 vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__dfrtp_1
X_10989_ net2489 net231 net435 vssd1 vssd1 vccd1 vccd1 _00054_ sky130_fd_sc_hd__mux2_1
X_12728_ _01431_ _06538_ columns.count\[10\] vssd1 vssd1 vccd1 vccd1 _06548_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_139_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07120__A2 _01954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12659_ datapath.mulitply_result\[24\] net502 net498 _06496_ vssd1 vssd1 vccd1 vccd1
+ _00934_ sky130_fd_sc_hd__a22o_1
XFILLER_90_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12773__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11897__B net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09948__A2 _03384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11389__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14329_ clknet_leaf_8_clk _01034_ net1072 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold405 datapath.rf.registers\[1\]\[2\] vssd1 vssd1 vccd1 vccd1 net1753 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08081__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold416 datapath.rf.registers\[22\]\[22\] vssd1 vssd1 vccd1 vccd1 net1764 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold427 datapath.rf.registers\[16\]\[30\] vssd1 vssd1 vccd1 vccd1 net1775 sky130_fd_sc_hd__dlygate4sd3_1
Xhold438 mmio.memload_or_instruction\[27\] vssd1 vssd1 vccd1 vccd1 net1786 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07168__A _01981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold449 datapath.rf.registers\[15\]\[16\] vssd1 vssd1 vccd1 vccd1 net1797 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout907 _01805_ vssd1 vssd1 vccd1 vccd1 net907 sky130_fd_sc_hd__buf_2
X_09870_ _04685_ _04705_ _04683_ vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_55_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout918 _01764_ vssd1 vssd1 vccd1 vccd1 net918 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07187__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout929 _01727_ vssd1 vssd1 vccd1 vccd1 net929 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ net554 net550 vssd1 vssd1 vccd1 vccd1 _03657_ sky130_fd_sc_hd__nor2_1
XFILLER_100_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1105 screen.counter.currentCt\[13\] vssd1 vssd1 vccd1 vccd1 net2453 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06934__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13109__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1116 datapath.rf.registers\[27\]\[7\] vssd1 vssd1 vccd1 vccd1 net2464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1127 datapath.rf.registers\[23\]\[6\] vssd1 vssd1 vccd1 vccd1 net2475 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08752_ _03502_ _03504_ _03585_ _03500_ _03498_ vssd1 vssd1 vccd1 vccd1 _03588_ sky130_fd_sc_hd__a311o_1
Xhold1138 datapath.rf.registers\[20\]\[12\] vssd1 vssd1 vccd1 vccd1 net2486 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1149 datapath.multiplication_module.multiplicand_i\[3\] vssd1 vssd1 vccd1 vccd1
+ net2497 sky130_fd_sc_hd__dlygate4sd3_1
X_07703_ datapath.rf.registers\[12\]\[17\] net756 net740 datapath.rf.registers\[16\]\[17\]
+ _02528_ vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__a221o_1
X_08683_ _02612_ _02635_ vssd1 vssd1 vccd1 vccd1 _03519_ sky130_fd_sc_hd__nand2_1
XANTENNA__12948__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout175_A _05684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07634_ datapath.rf.registers\[1\]\[18\] net762 net746 datapath.rf.registers\[17\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__a22o_1
XANTENNA__07895__B1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09830__B net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07631__A _02466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07565_ datapath.rf.registers\[31\]\[19\] net977 net916 vssd1 vssd1 vccd1 vccd1 _02401_
+ sky130_fd_sc_hd__and3_1
XFILLER_81_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08439__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1084_A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09304_ net319 _03906_ _04139_ net324 vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__a211o_1
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07647__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07496_ net613 _02331_ net565 vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13305__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09235_ _03930_ _04070_ net354 vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1251_A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout607_A _03608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09166_ net649 _04001_ net439 vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__a21o_1
XANTENNA__08462__A _03262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11299__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08117_ datapath.rf.registers\[5\]\[8\] net820 net814 datapath.rf.registers\[23\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02953_ sky130_fd_sc_hd__a22o_1
XANTENNA__08072__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09097_ net347 _03932_ vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__or2_1
X_08048_ datapath.rf.registers\[29\]\[9\] net977 net918 vssd1 vssd1 vccd1 vccd1 _02884_
+ sky130_fd_sc_hd__and3_1
XFILLER_123_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold950 datapath.rf.registers\[2\]\[29\] vssd1 vssd1 vccd1 vccd1 net2298 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07509__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold961 datapath.rf.registers\[27\]\[12\] vssd1 vssd1 vccd1 vccd1 net2309 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout976_A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold972 datapath.rf.registers\[23\]\[9\] vssd1 vssd1 vccd1 vccd1 net2320 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold983 datapath.rf.registers\[28\]\[8\] vssd1 vssd1 vccd1 vccd1 net2331 sky130_fd_sc_hd__dlygate4sd3_1
Xhold994 datapath.rf.registers\[22\]\[9\] vssd1 vssd1 vccd1 vccd1 net2342 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07178__A2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10010_ _04844_ _04845_ vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__nand2_1
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10182__A1 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout764_X net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09999_ _04762_ _04799_ vssd1 vssd1 vccd1 vccd1 _04835_ sky130_fd_sc_hd__xnor2_2
XFILLER_131_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13019__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06925__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11961_ _05323_ _06003_ _06006_ screen.controlBus\[7\] vssd1 vssd1 vccd1 vccd1 _06007_
+ sky130_fd_sc_hd__a22o_1
XFILLER_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout931_X net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12858__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10912_ _05654_ _05655_ vssd1 vssd1 vccd1 vccd1 _05656_ sky130_fd_sc_hd__or2_1
XFILLER_72_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13700_ clknet_leaf_23_clk _00510_ net1154 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_14680_ clknet_leaf_6_clk _01385_ net1067 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[6\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07886__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09740__B _03818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11892_ net136 _05958_ _05957_ vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07350__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13631_ clknet_leaf_11_clk _00441_ net1081 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10843_ net900 _04177_ _05596_ net616 vssd1 vssd1 vccd1 vccd1 _05597_ sky130_fd_sc_hd__o211a_1
XANTENNA__07638__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13562_ clknet_leaf_2_clk _00372_ net1078 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10774_ net898 _05537_ net616 vssd1 vssd1 vccd1 vccd1 _05538_ sky130_fd_sc_hd__o21a_1
XANTENNA__07102__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11985__A2 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12513_ datapath.multiplication_module.multiplier_i\[0\] net572 vssd1 vssd1 vccd1
+ vccd1 _06374_ sky130_fd_sc_hd__nor2_1
X_13493_ clknet_leaf_20_clk _00303_ net1117 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_12444_ net167 _05936_ net129 net2551 vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_67_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12375_ screen.counter.ack3 screen.counter.ack2 vssd1 vssd1 vccd1 vccd1 _06334_ sky130_fd_sc_hd__nand2b_1
XFILLER_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14114_ clknet_leaf_100_clk screen.register.controlFill net1228 vssd1 vssd1 vccd1
+ vccd1 screen.register.cFill1 sky130_fd_sc_hd__dfrtp_1
X_11326_ net1994 net241 net416 vssd1 vssd1 vccd1 vccd1 _00371_ sky130_fd_sc_hd__mux2_1
XFILLER_141_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14045_ clknet_leaf_107_clk _00813_ net1220 vssd1 vssd1 vccd1 vccd1 screen.counter.currentEnable
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_130_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11257_ net245 net2390 net418 vssd1 vssd1 vccd1 vccd1 _00306_ sky130_fd_sc_hd__mux2_1
XANTENNA__07169__A2 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10208_ _03743_ _05043_ net1041 vssd1 vssd1 vccd1 vccd1 _05044_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10845__A1_N _05597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11188_ net252 net1912 net422 vssd1 vssd1 vccd1 vccd1 _00240_ sky130_fd_sc_hd__mux2_1
XFILLER_68_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10139_ _04833_ _04877_ vssd1 vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__xnor2_1
XFILLER_83_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09315__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12768__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11673__A1 _05211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07877__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07341__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13829_ clknet_leaf_113_clk _00638_ net1197 vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09618__B2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07170__B net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07350_ datapath.rf.registers\[14\]\[24\] net775 net742 datapath.rf.registers\[2\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__a22o_1
X_07281_ datapath.rf.registers\[22\]\[25\] net823 _02099_ _02102_ _02104_ vssd1 vssd1
+ vccd1 vccd1 _02117_ sky130_fd_sc_hd__a2111o_1
XFILLER_148_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_151_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_151_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09020_ net344 _03710_ _03855_ vssd1 vssd1 vccd1 vccd1 _03856_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09378__A _02612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11728__A2 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold202 datapath.rf.registers\[19\]\[1\] vssd1 vssd1 vccd1 vccd1 net1550 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10936__B1 _05675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold213 datapath.multiplication_module.multiplicand_i\[19\] vssd1 vssd1 vccd1 vccd1
+ net1561 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold224 datapath.multiplication_module.multiplicand_i\[17\] vssd1 vssd1 vccd1 vccd1
+ net1572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 datapath.rf.registers\[18\]\[20\] vssd1 vssd1 vccd1 vccd1 net1583 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold246 datapath.rf.registers\[8\]\[3\] vssd1 vssd1 vccd1 vccd1 net1594 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold257 datapath.rf.registers\[12\]\[7\] vssd1 vssd1 vccd1 vccd1 net1605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 datapath.rf.registers\[23\]\[0\] vssd1 vssd1 vccd1 vccd1 net1616 sky130_fd_sc_hd__dlygate4sd3_1
Xhold279 datapath.rf.registers\[22\]\[7\] vssd1 vssd1 vccd1 vccd1 net1627 sky130_fd_sc_hd__dlygate4sd3_1
X_09922_ datapath.PC\[10\] _02877_ vssd1 vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__nand2_1
Xfanout704 net705 vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__clkbuf_8
Xfanout715 net717 vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__buf_4
Xfanout726 _01812_ vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__buf_4
XFILLER_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09853_ _03457_ _03502_ _03951_ vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__or3b_1
Xfanout737 _01810_ vssd1 vssd1 vccd1 vccd1 net737 sky130_fd_sc_hd__clkbuf_4
XFILLER_113_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10164__A1 _04177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout748 net749 vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__buf_4
Xfanout759 _01802_ vssd1 vssd1 vccd1 vccd1 net759 sky130_fd_sc_hd__buf_2
XFILLER_140_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08804_ _03611_ _03638_ vssd1 vssd1 vccd1 vccd1 _03640_ sky130_fd_sc_hd__or2_1
XFILLER_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09784_ _03490_ net627 net624 _03491_ net644 vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__a221o_1
X_06996_ net963 _01831_ vssd1 vssd1 vccd1 vccd1 _01832_ sky130_fd_sc_hd__and2_2
XFILLER_39_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08735_ _03530_ _03531_ _03570_ vssd1 vssd1 vccd1 vccd1 _03571_ sky130_fd_sc_hd__and3_1
XFILLER_73_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12310__C1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout557_A _03418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08666_ _02285_ _02286_ vssd1 vssd1 vccd1 vccd1 _03502_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_68_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07999__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08457__A net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07617_ datapath.rf.registers\[14\]\[18\] net829 net804 datapath.rf.registers\[28\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_101_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10198__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08597_ _02960_ _02983_ vssd1 vssd1 vccd1 vccd1 _03433_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout345_X net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout724_A net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07548_ _02376_ _02378_ _02383_ vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__or3_4
XANTENNA__08817__C1 _03384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08293__B1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07479_ datapath.rf.registers\[30\]\[21\] net758 net702 datapath.rf.registers\[9\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_142_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_142_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout512_X net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10926__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1254_X net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08832__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11611__A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09218_ _01620_ _04024_ _04053_ net318 _04051_ vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__o221a_1
XFILLER_10_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10490_ screen.controlBus\[0\] screen.controlBus\[1\] _05314_ _05318_ vssd1 vssd1
+ vccd1 vccd1 _05320_ sky130_fd_sc_hd__and4b_1
XANTENNA__06705__A datapath.ru.latched_instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09149_ _03765_ _03919_ net368 vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__mux2_1
XFILLER_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07399__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12160_ _06178_ _06186_ vssd1 vssd1 vccd1 vccd1 _06187_ sky130_fd_sc_hd__nor2_1
XANTENNA__12392__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout881_X net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11111_ net299 net1779 net427 vssd1 vssd1 vccd1 vccd1 _00166_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout979_X net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12091_ _06120_ _06125_ _06126_ _06129_ vssd1 vssd1 vccd1 vccd1 _06130_ sky130_fd_sc_hd__or4_1
Xhold780 datapath.rf.registers\[7\]\[15\] vssd1 vssd1 vccd1 vccd1 net2128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold791 datapath.rf.registers\[29\]\[30\] vssd1 vssd1 vccd1 vccd1 net2139 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_112_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09227__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11042_ net298 net1962 net430 vssd1 vssd1 vccd1 vccd1 _00102_ sky130_fd_sc_hd__mux2_1
XFILLER_131_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07020__A1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07571__A2 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input20_A DAT_I[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12993_ net168 net2529 net479 vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__mux2_1
XFILLER_92_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11492__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07859__B1 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11944_ screen.register.currentYbus\[29\] net160 vssd1 vssd1 vccd1 vccd1 _05993_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__08367__A net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11875_ screen.register.currentYbus\[6\] net161 vssd1 vssd1 vccd1 vccd1 _05947_ sky130_fd_sc_hd__nand2_1
X_14663_ clknet_leaf_143_clk _01368_ net1093 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13614_ clknet_leaf_5_clk _00424_ net1067 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10826_ net256 net1589 net544 vssd1 vssd1 vccd1 vccd1 _00015_ sky130_fd_sc_hd__mux2_1
X_14594_ clknet_leaf_152_clk _01299_ net1054 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_119_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08284__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13545_ clknet_leaf_62_clk _00355_ net1234 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10757_ net303 net2174 net544 vssd1 vssd1 vccd1 vccd1 _00005_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_133_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_133_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09481__C1 _02913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13476_ clknet_leaf_21_clk _00286_ net1163 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10688_ net1013 _05503_ _05476_ vssd1 vssd1 vccd1 vccd1 _05505_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_132_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12427_ _05984_ net158 vssd1 vssd1 vccd1 vccd1 _06361_ sky130_fd_sc_hd__nor2_1
XFILLER_142_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09784__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12358_ datapath.PC\[28\] net309 _06320_ _06322_ vssd1 vssd1 vccd1 vccd1 _00807_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08830__A _03636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11309_ net1547 net208 net417 vssd1 vssd1 vccd1 vccd1 _00354_ sky130_fd_sc_hd__mux2_1
XFILLER_141_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12289_ net636 _04534_ _04536_ net308 vssd1 vssd1 vccd1 vccd1 _06273_ sky130_fd_sc_hd__a31o_1
XFILLER_141_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14028_ clknet_leaf_80_clk _00797_ net1257 vssd1 vssd1 vccd1 vccd1 datapath.PC\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_68_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06850_ datapath.ru.latched_instruction\[26\] _01595_ net971 datapath.ru.latched_instruction\[24\]
+ _01685_ vssd1 vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__a221o_1
XFILLER_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_147_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06781_ datapath.ru.latched_instruction\[13\] net1031 net994 _01615_ vssd1 vssd1
+ vccd1 vccd1 _01618_ sky130_fd_sc_hd__a22oi_4
XANTENNA__12498__S net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08520_ _03345_ _03347_ _03351_ _03355_ vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__or4_1
X_08451_ _03284_ _03285_ _03286_ vssd1 vssd1 vccd1 vccd1 _03287_ sky130_fd_sc_hd__or3_1
XANTENNA__07612__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07402_ datapath.rf.registers\[0\]\[23\] net782 _02223_ _02237_ vssd1 vssd1 vccd1
+ vccd1 _02238_ sky130_fd_sc_hd__o22ai_2
X_08382_ datapath.rf.registers\[18\]\[3\] net725 net700 datapath.rf.registers\[23\]\[3\]
+ _03217_ vssd1 vssd1 vccd1 vccd1 _03218_ sky130_fd_sc_hd__a221o_1
XFILLER_149_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07333_ datapath.rf.registers\[0\]\[24\] net871 _02159_ _02168_ vssd1 vssd1 vccd1
+ vccd1 _02169_ sky130_fd_sc_hd__o22a_4
XTAP_TAPCELL_ROW_34_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08275__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_124_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_124_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_63_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13122__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout138_A net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07264_ datapath.rf.registers\[13\]\[25\] net986 net918 vssd1 vssd1 vccd1 vccd1 _02100_
+ sky130_fd_sc_hd__and3_1
XFILLER_137_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09003_ net331 _03838_ net312 vssd1 vssd1 vccd1 vccd1 _03839_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08027__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07195_ datapath.rf.registers\[24\]\[27\] net767 net751 datapath.rf.registers\[28\]\[27\]
+ _02029_ vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__a221o_1
XFILLER_133_902 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12262__A _05002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout501 _06375_ vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__buf_2
XFILLER_59_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09905_ _01585_ net900 _01678_ vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__and3_1
XFILLER_99_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout512 _05735_ vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__clkbuf_8
XFILLER_59_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout523 _05723_ vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__clkbuf_4
Xfanout534 net535 vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__buf_4
Xfanout545 _05519_ vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__buf_4
Xfanout556 _03609_ vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__clkbuf_2
Xfanout567 _06171_ vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__buf_2
X_09836_ _03513_ _03518_ _04085_ _04119_ vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__or4b_1
Xfanout578 net580 vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__buf_2
XFILLER_86_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09767_ _04084_ _04118_ _04586_ _04600_ vssd1 vssd1 vccd1 vccd1 _04603_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout841_A net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06979_ net968 net911 _01809_ vssd1 vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__and3_1
XFILLER_55_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07803__B net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08718_ _03544_ _03553_ vssd1 vssd1 vccd1 vccd1 _03554_ sky130_fd_sc_hd__nand2b_1
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09698_ net630 _04533_ vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_83_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07305__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14095__RESET_B net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08649_ _01980_ _02003_ vssd1 vssd1 vccd1 vccd1 _03485_ sky130_fd_sc_hd__and2_1
XFILLER_15_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout727_X net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11660_ net1454 _05875_ _05879_ vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__a21o_1
XFILLER_148_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10611_ button\[0\] _01435_ vssd1 vssd1 vccd1 vccd1 _05431_ sky130_fd_sc_hd__and2_1
X_11591_ screen.counter.ct\[16\] _05296_ _05814_ net1270 vssd1 vssd1 vccd1 vccd1 _05815_
+ sky130_fd_sc_hd__or4b_1
Xclkbuf_leaf_115_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_115_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_12_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13032__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13330_ clknet_leaf_32_clk _00140_ net1122 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10542_ datapath.multiplication_module.multiplier_i\[1\] datapath.multiplication_module.multiplier_i\[0\]
+ datapath.multiplication_module.multiplier_i\[3\] datapath.multiplication_module.multiplier_i\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05370_ sky130_fd_sc_hd__or4_1
XANTENNA__08353__C _01712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13261_ clknet_leaf_132_clk _00071_ net1113 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_98_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10473_ _05294_ _05302_ vssd1 vssd1 vccd1 vccd1 _05303_ sky130_fd_sc_hd__or2_1
XANTENNA__09215__C1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12871__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12212_ _06217_ _06218_ vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__nor2_1
XANTENNA__12365__A2 _06254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13192_ datapath.rf.registers\[0\]\[29\] vssd1 vssd1 vccd1 vccd1 _01014_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08650__A _01980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10376__A1 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11487__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12143_ _06000_ net1012 net567 vssd1 vssd1 vccd1 vccd1 _06176_ sky130_fd_sc_hd__a21o_1
XFILLER_2_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07792__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12074_ screen.register.currentXbus\[13\] _05768_ _06019_ screen.register.currentYbus\[13\]
+ _06104_ vssd1 vssd1 vccd1 vccd1 _06114_ sky130_fd_sc_hd__a221o_1
X_11025_ net214 net2460 net538 vssd1 vssd1 vccd1 vccd1 _00087_ sky130_fd_sc_hd__mux2_1
XFILLER_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10898__Y _05644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07544__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07713__B net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12976_ net251 net2510 net479 vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__mux2_1
XFILLER_73_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_142_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11927_ net465 screen.counter.ack vssd1 vssd1 vccd1 vccd1 _05982_ sky130_fd_sc_hd__or2_1
X_14646_ clknet_leaf_141_clk _01351_ net1095 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_11858_ _03417_ net658 vssd1 vssd1 vccd1 vccd1 _05936_ sky130_fd_sc_hd__nand2_1
XFILLER_14_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10809_ _04300_ _05567_ net899 vssd1 vssd1 vccd1 vccd1 _05568_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_106_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_106_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_19 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11789_ net1291 _05747_ _05900_ vssd1 vssd1 vccd1 vccd1 _05901_ sky130_fd_sc_hd__mux2_1
XFILLER_14_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14577_ clknet_leaf_40_clk _01282_ net1140 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13528_ clknet_leaf_3_clk _00338_ net1076 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_119_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13747__RESET_B net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12781__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13459_ clknet_leaf_34_clk _00269_ net1127 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_115_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 DAT_O[9] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_71_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput115 net115 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__buf_2
XANTENNA__11397__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06999__B _01831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09509__A0 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07783__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07951_ datapath.rf.registers\[19\]\[11\] net977 net928 vssd1 vssd1 vccd1 vccd1 _02787_
+ sky130_fd_sc_hd__and3_1
XFILLER_101_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06902_ net976 net944 vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__and2_1
X_07882_ datapath.rf.registers\[26\]\[13\] net779 _02717_ net787 vssd1 vssd1 vccd1
+ vccd1 _02718_ sky130_fd_sc_hd__a211o_1
XANTENNA_clkbuf_leaf_86_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07535__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06833_ datapath.ru.latched_instruction\[25\] net1046 net1016 net993 vssd1 vssd1
+ vccd1 vccd1 _01669_ sky130_fd_sc_hd__and4b_1
XFILLER_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09621_ net460 _04353_ _04352_ net354 vssd1 vssd1 vccd1 vccd1 _04457_ sky130_fd_sc_hd__a211o_1
XANTENNA__07904__A net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13117__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09552_ _04385_ _04387_ net378 vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__mux2_1
X_06764_ _01593_ _01594_ _01599_ _01600_ vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_65_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08503_ datapath.rf.registers\[17\]\[1\] _01800_ net907 vssd1 vssd1 vccd1 vccd1 _03339_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_65_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08438__C _01816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09483_ net557 net576 net546 _03009_ vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__o211a_1
X_06695_ net1287 net1284 mmio.memload_or_instruction\[28\] vssd1 vssd1 vccd1 vccd1
+ _01534_ sky130_fd_sc_hd__nor3b_1
XANTENNA__12956__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_144_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08434_ datapath.rf.registers\[10\]\[2\] net969 net909 net908 vssd1 vssd1 vccd1 vccd1
+ _03270_ sky130_fd_sc_hd__and4_1
XFILLER_51_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08365_ datapath.rf.registers\[19\]\[3\] net854 _01753_ datapath.rf.registers\[6\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_24_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout422_A net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07316_ datapath.rf.registers\[4\]\[24\] net958 net933 vssd1 vssd1 vccd1 vccd1 _02152_
+ sky130_fd_sc_hd__and3_1
XFILLER_20_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08296_ datapath.rf.registers\[10\]\[4\] net880 net798 datapath.rf.registers\[29\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__a22o_1
XANTENNA__09460__A2 _03859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07247_ datapath.rf.registers\[10\]\[26\] net706 net691 datapath.rf.registers\[13\]\[26\]
+ _02082_ vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__a221o_1
Xclkbuf_4_2_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_2_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout308_X net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_39_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07178_ datapath.rf.registers\[20\]\[27\] net839 net824 datapath.rf.registers\[6\]\[27\]
+ _02013_ vssd1 vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__a221o_1
XANTENNA__12263__Y _06253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout791_A net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10358__A1 net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout889_A _01713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10505__A _05315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06702__B datapath.ru.latched_instruction\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11100__S net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1217_X net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout320 _03684_ vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__buf_2
XANTENNA_fanout677_X net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout331 _03619_ vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__buf_2
Xfanout342 net343 vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__clkbuf_2
Xfanout353 net355 vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__buf_2
Xfanout364 net365 vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__buf_2
Xfanout375 _03625_ vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__clkbuf_2
XFILLER_143_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout386 net389 vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__clkbuf_8
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09819_ _04654_ _03783_ net450 vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__mux2_1
Xfanout397 _06555_ vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__buf_2
XANTENNA_fanout844_X net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14205__RESET_B net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12830_ net209 net2563 net489 vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08348__C net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ net1844 net172 net404 vssd1 vssd1 vccd1 vccd1 _00983_ sky130_fd_sc_hd__mux2_1
XANTENNA__12866__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14500_ clknet_leaf_22_clk _01205_ net1156 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11712_ net29 net1035 net1025 net2442 vssd1 vssd1 vccd1 vccd1 _00593_ sky130_fd_sc_hd__a22o_1
X_12692_ _06517_ _06519_ vssd1 vssd1 vccd1 vccd1 _06524_ sky130_fd_sc_hd__nor2_1
XANTENNA__08645__A _01888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11643_ _05788_ _05866_ vssd1 vssd1 vccd1 vccd1 _05867_ sky130_fd_sc_hd__or2_1
X_14431_ clknet_leaf_10_clk _01136_ net1080 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11574_ net1008 _05783_ _05787_ net1007 _05797_ vssd1 vssd1 vccd1 vccd1 _05798_ sky130_fd_sc_hd__o221a_1
X_14362_ clknet_leaf_2_clk _01067_ net1063 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput17 DAT_I[23] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
Xinput28 DAT_I[4] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11794__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput39 nrst vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_1
X_10525_ screen.counter.ct\[5\] _05349_ vssd1 vssd1 vccd1 vccd1 _05355_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_96_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13313_ clknet_leaf_46_clk _00123_ net1147 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_14293_ clknet_leaf_94_clk _00998_ net1217 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12338__A2 _03978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13244_ clknet_leaf_7_clk _00054_ net1071 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07548__X _02384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09739__B1 _03667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10456_ _01419_ _05289_ vssd1 vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__or2_1
XFILLER_6_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13175_ net2586 vssd1 vssd1 vccd1 vccd1 _00997_ sky130_fd_sc_hd__clkbuf_1
X_10387_ net381 _04156_ _05222_ _03614_ vssd1 vssd1 vccd1 vccd1 _05223_ sky130_fd_sc_hd__a211o_1
XANTENNA__11010__S net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12126_ _06162_ vssd1 vssd1 vccd1 vccd1 _06163_ sky130_fd_sc_hd__inv_2
XANTENNA__07765__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12057_ screen.register.currentYbus\[12\] _05776_ net996 screen.register.currentXbus\[28\]
+ vssd1 vssd1 vccd1 vccd1 _06098_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_127_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11008_ net301 net2286 net539 vssd1 vssd1 vccd1 vccd1 _00070_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_144_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08190__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08478__B1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12776__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12959_ net174 net1901 net396 vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__mux2_1
XANTENNA__06627__X _01466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14629_ clknet_leaf_117_clk _01334_ net1188 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12026__B2 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09427__C1 _03613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08150_ datapath.rf.registers\[11\]\[7\] net987 net938 vssd1 vssd1 vccd1 vccd1 _02986_
+ sky130_fd_sc_hd__and3_1
XFILLER_119_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07101_ datapath.rf.registers\[16\]\[29\] net739 net698 datapath.rf.registers\[23\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__a22o_1
X_08081_ datapath.rf.registers\[29\]\[9\] net677 net662 datapath.rf.registers\[5\]\[9\]
+ _02915_ vssd1 vssd1 vccd1 vccd1 _02917_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_155_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12329__A2 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07032_ datapath.rf.registers\[17\]\[30\] net851 _01865_ _01866_ _01867_ vssd1 vssd1
+ vccd1 vccd1 _01868_ sky130_fd_sc_hd__a2111o_1
XFILLER_142_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07756__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08953__A1 _02419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08983_ _03485_ net628 net624 _03486_ net644 vssd1 vssd1 vccd1 vccd1 _03819_ sky130_fd_sc_hd__a221o_1
XFILLER_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07934_ _02756_ _02766_ _02768_ _02769_ vssd1 vssd1 vccd1 vccd1 _02770_ sky130_fd_sc_hd__or4_1
XFILLER_84_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07865_ datapath.rf.registers\[23\]\[13\] net814 net801 datapath.rf.registers\[3\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02701_ sky130_fd_sc_hd__a22o_1
XFILLER_96_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09604_ net367 _04289_ _04439_ vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__o21a_1
XANTENNA__08181__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06816_ _01616_ _01617_ datapath.ru.latched_instruction\[13\] vssd1 vssd1 vccd1 vccd1
+ _01652_ sky130_fd_sc_hd__mux2_1
X_07796_ _02620_ _02625_ _02629_ _02631_ vssd1 vssd1 vccd1 vccd1 _02632_ sky130_fd_sc_hd__and4b_1
XFILLER_83_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06747_ _01585_ vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__inv_2
XFILLER_37_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09535_ net557 net576 net546 _02857_ vssd1 vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__o211a_1
XANTENNA__08469__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12265__A1 _05002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout637_A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09466_ net631 _04301_ vssd1 vssd1 vccd1 vccd1 _04302_ sky130_fd_sc_hd__nand2_1
X_06678_ datapath.ru.latched_instruction\[8\] _01467_ _01470_ datapath.ru.latched_instruction\[19\]
+ vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__a22o_1
XANTENNA__07141__B1 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08417_ datapath.rf.registers\[2\]\[2\] net889 net848 datapath.rf.registers\[1\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__a22o_1
XFILLER_11_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09397_ net332 _04225_ _04232_ _03613_ vssd1 vssd1 vccd1 vccd1 _04233_ sky130_fd_sc_hd__o211a_1
XFILLER_12_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout804_A net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout425_X net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08348_ datapath.rf.registers\[7\]\[3\] net942 net936 vssd1 vssd1 vccd1 vccd1 _03184_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09433__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08279_ datapath.rf.registers\[10\]\[5\] net707 net692 datapath.rf.registers\[13\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03115_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_78_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10310_ net1266 net1249 _05142_ _05145_ vssd1 vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__o22a_1
XFILLER_137_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11290_ net245 net2192 net522 vssd1 vssd1 vccd1 vccd1 _00338_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout794_X net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10241_ _04396_ _04428_ vssd1 vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_91_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10200__B1 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07747__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08944__A1 _02217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10172_ datapath.PC\[16\] net1294 _05000_ _05007_ vssd1 vssd1 vccd1 vccd1 _05008_
+ sky130_fd_sc_hd__a22o_1
XFILLER_121_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1104 net1110 vssd1 vssd1 vccd1 vccd1 net1104 sky130_fd_sc_hd__clkbuf_4
Xfanout1115 net1120 vssd1 vssd1 vccd1 vccd1 net1115 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1126 net1153 vssd1 vssd1 vccd1 vccd1 net1126 sky130_fd_sc_hd__clkbuf_2
XFILLER_121_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1137 net1139 vssd1 vssd1 vccd1 vccd1 net1137 sky130_fd_sc_hd__clkbuf_4
Xfanout150 net151 vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__clkbuf_4
Xfanout1148 net1152 vssd1 vssd1 vccd1 vccd1 net1148 sky130_fd_sc_hd__clkbuf_2
Xfanout161 _05933_ vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__clkbuf_2
Xfanout1159 net1162 vssd1 vssd1 vccd1 vccd1 net1159 sky130_fd_sc_hd__buf_2
XFILLER_59_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout172 _05684_ vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_109_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13931_ clknet_leaf_110_clk _00709_ net1222 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout183 net184 vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__clkbuf_2
Xfanout194 net195 vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__clkbuf_2
XFILLER_75_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11700__B1 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07263__B net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13862_ clknet_leaf_71_clk _00666_ net1244 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_16_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12813_ net1673 net244 net490 vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_122_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13793_ clknet_leaf_74_clk _00602_ net1247 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12744_ net1536 net255 net405 vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__mux2_1
XANTENNA__07132__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12675_ _06507_ _06508_ _06509_ vssd1 vssd1 vccd1 vccd1 _06510_ sky130_fd_sc_hd__or3_1
XANTENNA__07710__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11005__S net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14414_ clknet_leaf_1_clk _01119_ net1057 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_42_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11626_ _05803_ _05804_ _05805_ vssd1 vssd1 vccd1 vccd1 _05850_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_100_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14345_ clknet_leaf_92_clk _01050_ net1232 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11557_ net1008 _05780_ vssd1 vssd1 vccd1 vccd1 _05781_ sky130_fd_sc_hd__nor2_1
XANTENNA__09918__B net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire562 _02437_ vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07986__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10508_ net1277 screen.counter.ct\[11\] screen.counter.ct\[19\] vssd1 vssd1 vccd1
+ vccd1 _05338_ sky130_fd_sc_hd__nor3_1
Xhold609 datapath.rf.registers\[14\]\[28\] vssd1 vssd1 vccd1 vccd1 net1957 sky130_fd_sc_hd__dlygate4sd3_1
Xwire584 _02959_ vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__clkbuf_1
X_14276_ clknet_leaf_22_clk _00981_ net1154 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11488_ net270 net1910 net512 vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__mux2_1
X_13227_ clknet_leaf_56_clk _00037_ net1158 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10439_ _01702_ _04338_ _05274_ net1039 vssd1 vssd1 vccd1 vccd1 _05275_ sky130_fd_sc_hd__o211a_1
XANTENNA__07199__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07738__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13158_ net1648 net172 net383 vssd1 vssd1 vccd1 vccd1 _01399_ sky130_fd_sc_hd__mux2_1
XFILLER_112_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12109_ screen.counter.currentCt\[0\] screen.counter.currentCt\[3\] screen.counter.currentCt\[2\]
+ screen.counter.currentCt\[1\] vssd1 vssd1 vccd1 vccd1 _06146_ sky130_fd_sc_hd__or4b_1
X_13089_ net1715 net185 net387 vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__mux2_1
XFILLER_26_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09360__A1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08163__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07650_ _02476_ _02485_ vssd1 vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_0_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06601_ net1286 net1281 mmio.key_data\[5\] vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__o21a_1
XFILLER_93_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07581_ _02410_ _02414_ _02416_ vssd1 vssd1 vccd1 vccd1 _02417_ sky130_fd_sc_hd__or3_4
XFILLER_80_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_730 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09320_ _03923_ _04155_ net377 vssd1 vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__mux2_1
XANTENNA__10258__B1 net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13762__RESET_B net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06827__A1_N _01467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09251_ _03581_ _04085_ vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__xnor2_1
X_08202_ datapath.rf.registers\[6\]\[6\] net954 net931 vssd1 vssd1 vccd1 vccd1 _03038_
+ sky130_fd_sc_hd__and3_1
XFILLER_138_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09182_ _04017_ vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__inv_2
X_08133_ datapath.rf.registers\[28\]\[8\] net752 net737 datapath.rf.registers\[22\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__a22o_1
XANTENNA__13130__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07977__A2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08064_ datapath.rf.registers\[12\]\[9\] _01749_ _02892_ _02895_ _02897_ vssd1 vssd1
+ vccd1 vccd1 _02900_ sky130_fd_sc_hd__a2111o_1
XFILLER_146_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07015_ datapath.rf.registers\[8\]\[31\] net694 net679 datapath.rf.registers\[6\]\[31\]
+ _01850_ vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__a221o_1
XANTENNA__09179__A1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07729__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08926__A1 _03418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06820__X _01656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08966_ _03800_ _03801_ net448 vssd1 vssd1 vccd1 vccd1 _03802_ sky130_fd_sc_hd__mux2_1
XFILLER_57_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08098__B1_N _02933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07917_ datapath.rf.registers\[14\]\[12\] net777 net713 datapath.rf.registers\[11\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout754_A net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08897_ net1269 datapath.PC\[3\] datapath.PC\[4\] vssd1 vssd1 vccd1 vccd1 _03733_
+ sky130_fd_sc_hd__or3_1
XFILLER_124_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_95_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_95_clk sky130_fd_sc_hd__clkbuf_8
X_07848_ datapath.rf.registers\[15\]\[13\] net983 net916 vssd1 vssd1 vccd1 vccd1 _02684_
+ sky130_fd_sc_hd__and3_1
XFILLER_16_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07651__X _02487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07901__A2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout542_X net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout921_A net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10929__S net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07779_ datapath.rf.registers\[14\]\[15\] net775 net743 datapath.rf.registers\[2\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02615_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_104_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09518_ net460 _04353_ _04352_ net351 vssd1 vssd1 vccd1 vccd1 _04354_ sky130_fd_sc_hd__a211o_1
X_10790_ _04515_ _05551_ net899 vssd1 vssd1 vccd1 vccd1 _05552_ sky130_fd_sc_hd__mux2_1
XANTENNA__07114__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08195__A _03009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12429__B net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09449_ net325 _03847_ _04284_ vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout807_X net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12460_ net166 _05968_ net128 screen.register.currentXbus\[16\] vssd1 vssd1 vccd1
+ vccd1 _00862_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_130_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08923__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11749__B1 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11411_ net258 net1656 net517 vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__mux2_1
X_12391_ _05948_ net157 vssd1 vssd1 vccd1 vccd1 _06343_ sky130_fd_sc_hd__nor2_1
XANTENNA__13040__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07098__X _01934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10421__A0 _03262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14130_ clknet_leaf_35_clk _00887_ net1127 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11342_ _05518_ _05727_ vssd1 vssd1 vccd1 vccd1 _05728_ sky130_fd_sc_hd__or2_1
XFILLER_125_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14061_ clknet_leaf_121_clk _00828_ net1199 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07258__B _02091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11273_ _05517_ _05715_ vssd1 vssd1 vccd1 vccd1 _05723_ sky130_fd_sc_hd__nand2_4
X_13012_ net1748 net240 net392 vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__mux2_1
X_10224_ net229 _04899_ _05059_ net1258 vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__o31a_1
XFILLER_140_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10724__A1 _02856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11495__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10155_ net1041 _04988_ _04990_ vssd1 vssd1 vccd1 vccd1 _04991_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_7_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10086_ net1043 _03748_ vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__nand2_1
Xhold6 screen.counter.ack1 vssd1 vssd1 vccd1 vccd1 net1354 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_86_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_86_clk sky130_fd_sc_hd__clkbuf_8
X_13914_ clknet_leaf_43_clk _00003_ net1150 vssd1 vssd1 vccd1 vccd1 keypad.debounce.debounce\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07353__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13845_ clknet_leaf_51_clk net1281 net1182 vssd1 vssd1 vccd1 vccd1 mmio.key_en3 sky130_fd_sc_hd__dfrtp_1
XFILLER_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07105__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13776_ clknet_leaf_85_clk _00585_ net1258 vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__dfrtp_1
X_10988_ net1733 net237 net436 vssd1 vssd1 vccd1 vccd1 _00053_ sky130_fd_sc_hd__mux2_1
XFILLER_31_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12727_ _05893_ _06546_ _06547_ _06530_ vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__a31o_1
XFILLER_31_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_139_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12658_ _06493_ _06495_ vssd1 vssd1 vccd1 vccd1 _06496_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08392__X _03228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08833__A _01611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11609_ net998 net996 net995 _05793_ vssd1 vssd1 vccd1 vccd1 _05833_ sky130_fd_sc_hd__or4_1
X_12589_ _06436_ _06437_ vssd1 vssd1 vccd1 vccd1 _06438_ sky130_fd_sc_hd__nand2_1
XFILLER_144_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_10_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_152_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14328_ clknet_leaf_6_clk _01033_ net1068 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07449__A net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold406 datapath.rf.registers\[25\]\[22\] vssd1 vssd1 vccd1 vccd1 net1754 sky130_fd_sc_hd__dlygate4sd3_1
Xhold417 datapath.rf.registers\[19\]\[25\] vssd1 vssd1 vccd1 vccd1 net1765 sky130_fd_sc_hd__dlygate4sd3_1
Xhold428 datapath.rf.registers\[10\]\[25\] vssd1 vssd1 vccd1 vccd1 net1776 sky130_fd_sc_hd__dlygate4sd3_1
Xhold439 datapath.rf.registers\[26\]\[16\] vssd1 vssd1 vccd1 vccd1 net1787 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14259_ clknet_leaf_41_clk _00964_ net1141 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_55_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout908 _01793_ vssd1 vssd1 vccd1 vccd1 net908 sky130_fd_sc_hd__clkbuf_2
XFILLER_98_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout919 _01745_ vssd1 vssd1 vccd1 vccd1 net919 sky130_fd_sc_hd__buf_4
XFILLER_124_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08384__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08820_ net991 _03643_ vssd1 vssd1 vccd1 vccd1 _03656_ sky130_fd_sc_hd__or2_1
XFILLER_58_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1106 datapath.rf.registers\[1\]\[20\] vssd1 vssd1 vccd1 vccd1 net2454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1117 datapath.rf.registers\[30\]\[21\] vssd1 vssd1 vccd1 vccd1 net2465 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1128 screen.register.currentYbus\[12\] vssd1 vssd1 vccd1 vccd1 net2476 sky130_fd_sc_hd__dlygate4sd3_1
X_08751_ _03502_ _03504_ _03585_ _03500_ vssd1 vssd1 vccd1 vccd1 _03587_ sky130_fd_sc_hd__a31o_1
XFILLER_112_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_77_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_clk sky130_fd_sc_hd__clkbuf_8
Xhold1139 screen.register.currentYbus\[8\] vssd1 vssd1 vccd1 vccd1 net2487 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08136__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07702_ datapath.rf.registers\[2\]\[17\] net744 net685 datapath.rf.registers\[27\]\[17\]
+ _02537_ vssd1 vssd1 vccd1 vccd1 _02538_ sky130_fd_sc_hd__a221o_1
X_08682_ _02589_ _02590_ vssd1 vssd1 vccd1 vccd1 _03518_ sky130_fd_sc_hd__or2_2
XANTENNA__07344__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07633_ datapath.rf.registers\[12\]\[18\] net754 net698 datapath.rf.registers\[23\]\[18\]
+ _02468_ vssd1 vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__a221o_1
XFILLER_81_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13125__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06766__A1_N _01466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07564_ datapath.rf.registers\[15\]\[19\] net985 net916 vssd1 vssd1 vccd1 vccd1 _02400_
+ sky130_fd_sc_hd__and3_1
XFILLER_81_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09303_ net321 _03899_ vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_24_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07495_ _02321_ _02326_ _02330_ net782 datapath.rf.registers\[0\]\[21\] vssd1 vssd1
+ vccd1 vccd1 _02331_ sky130_fd_sc_hd__o32a_4
XANTENNA__12964__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1077_A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09234_ _03996_ _04069_ net459 vssd1 vssd1 vccd1 vccd1 _04070_ sky130_fd_sc_hd__mux2_1
XFILLER_22_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09165_ net345 _04000_ vssd1 vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__or2_1
XFILLER_147_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1244_A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08116_ datapath.rf.registers\[19\]\[8\] net854 net794 datapath.rf.registers\[31\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__a22o_1
X_09096_ net356 _03931_ vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__or2_1
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08047_ datapath.rf.registers\[10\]\[9\] net986 net937 vssd1 vssd1 vccd1 vccd1 _02883_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07078__B net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1032_X net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold940 datapath.rf.registers\[11\]\[31\] vssd1 vssd1 vccd1 vccd1 net2288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold951 datapath.rf.registers\[20\]\[8\] vssd1 vssd1 vccd1 vccd1 net2299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold962 datapath.rf.registers\[8\]\[12\] vssd1 vssd1 vccd1 vccd1 net2310 sky130_fd_sc_hd__dlygate4sd3_1
Xhold973 datapath.rf.registers\[5\]\[16\] vssd1 vssd1 vccd1 vccd1 net2321 sky130_fd_sc_hd__dlygate4sd3_1
Xhold984 datapath.rf.registers\[11\]\[29\] vssd1 vssd1 vccd1 vccd1 net2332 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09631__A1_N net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10706__A1 _02824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout871_A _01724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold995 datapath.rf.registers\[17\]\[0\] vssd1 vssd1 vccd1 vccd1 net2343 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout492_X net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout969_A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08375__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09998_ _04726_ _04813_ vssd1 vssd1 vccd1 vccd1 _04834_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07583__B1 _02417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08949_ _03784_ vssd1 vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__inv_2
XANTENNA__09324__A1 _02522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout757_X net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08127__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_68_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_clk sky130_fd_sc_hd__clkbuf_8
X_11960_ _05787_ _05852_ _05853_ _05783_ _05791_ vssd1 vssd1 vccd1 vccd1 _06006_ sky130_fd_sc_hd__o221a_1
XANTENNA__07335__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07381__X _02217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10911_ net1263 _05647_ vssd1 vssd1 vccd1 vccd1 _05655_ sky130_fd_sc_hd__nor2_1
XFILLER_45_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11891_ _02824_ net658 vssd1 vssd1 vccd1 vccd1 _05958_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_86_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout924_X net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13035__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13630_ clknet_leaf_148_clk _00440_ net1060 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10842_ net897 _05595_ vssd1 vssd1 vccd1 vccd1 _05596_ sky130_fd_sc_hd__or2_1
XFILLER_72_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12874__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13561_ clknet_leaf_9_clk _00371_ net1074 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07260__C net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10773_ net1268 _05530_ vssd1 vssd1 vccd1 vccd1 _05537_ sky130_fd_sc_hd__xnor2_1
X_12512_ _06372_ _06373_ vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__nor2_1
XANTENNA__09749__A _04178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13492_ clknet_leaf_93_clk _00302_ net1211 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08653__A _02025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12443_ net165 _05746_ vssd1 vssd1 vccd1 vccd1 _06369_ sky130_fd_sc_hd__and2_2
XFILLER_12_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06861__A2 _01604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12374_ _06333_ datapath.PC\[1\] net190 vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__mux2_1
X_14113_ clknet_leaf_100_clk screen.register.xFill net1228 vssd1 vssd1 vccd1 vccd1
+ screen.register.xFill1 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_10_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11325_ net1742 net246 net414 vssd1 vssd1 vccd1 vccd1 _00370_ sky130_fd_sc_hd__mux2_1
XFILLER_114_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14044_ clknet_leaf_99_clk net1372 net1229 vssd1 vssd1 vccd1 vccd1 screen.register.cFill3
+ sky130_fd_sc_hd__dfrtp_1
X_11256_ net248 net1931 net419 vssd1 vssd1 vccd1 vccd1 _00305_ sky130_fd_sc_hd__mux2_1
XFILLER_79_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09563__A1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10207_ datapath.PC\[17\] _03742_ datapath.PC\[18\] vssd1 vssd1 vccd1 vccd1 _05043_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__09563__B2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11187_ net255 net1783 net423 vssd1 vssd1 vccd1 vccd1 _00239_ sky130_fd_sc_hd__mux2_1
XFILLER_95_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10138_ net230 _04970_ _04973_ vssd1 vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__and3_1
XFILLER_94_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_59_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_76_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08118__A2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10069_ datapath.PC\[31\] net595 vssd1 vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07326__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13828_ clknet_leaf_116_clk _00637_ net1187 vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__dfrtp_1
XFILLER_90_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07170__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08826__A0 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13759_ clknet_leaf_76_clk _00568_ net1248 vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__dfrtp_1
XFILLER_149_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12784__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07280_ datapath.rf.registers\[8\]\[25\] net878 net838 datapath.rf.registers\[26\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__a22o_1
XANTENNA__06852__A2 _01593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold203 datapath.rf.registers\[15\]\[1\] vssd1 vssd1 vccd1 vccd1 net1551 sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 datapath.rf.registers\[4\]\[14\] vssd1 vssd1 vccd1 vccd1 net1562 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10936__B2 _05676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold225 datapath.rf.registers\[20\]\[31\] vssd1 vssd1 vccd1 vccd1 net1573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 datapath.rf.registers\[27\]\[18\] vssd1 vssd1 vccd1 vccd1 net1584 sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 datapath.rf.registers\[13\]\[1\] vssd1 vssd1 vccd1 vccd1 net1595 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 screen.counter.ct\[6\] vssd1 vssd1 vccd1 vccd1 net1606 sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ datapath.PC\[11\] _01786_ _04754_ _04755_ vssd1 vssd1 vccd1 vccd1 _04757_
+ sky130_fd_sc_hd__or4_2
Xhold269 datapath.rf.registers\[3\]\[2\] vssd1 vssd1 vccd1 vccd1 net1617 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout705 _01819_ vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09554__A1 _03770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08357__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout716 net717 vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__clkbuf_8
Xfanout727 _01812_ vssd1 vssd1 vccd1 vccd1 net727 sky130_fd_sc_hd__clkbuf_4
X_09852_ _02441_ _04686_ _04687_ _04671_ vssd1 vssd1 vccd1 vccd1 _04688_ sky130_fd_sc_hd__a31o_1
Xfanout738 net741 vssd1 vssd1 vccd1 vccd1 net738 sky130_fd_sc_hd__buf_4
Xfanout749 _01806_ vssd1 vssd1 vccd1 vccd1 net749 sky130_fd_sc_hd__clkbuf_4
XFILLER_58_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08803_ _03638_ vssd1 vssd1 vccd1 vccd1 _03639_ sky130_fd_sc_hd__inv_2
X_09783_ net320 _04593_ _04618_ net322 vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__a211o_1
XANTENNA__12959__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06995_ net991 _01637_ net990 net972 vssd1 vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__and4_2
XANTENNA__08109__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout285_A _05547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08734_ _03536_ _03537_ _03567_ _03534_ _03533_ vssd1 vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__a311o_1
X_08665_ net563 _02284_ vssd1 vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_68_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1194_A net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07616_ datapath.rf.registers\[26\]\[18\] net836 net815 datapath.rf.registers\[21\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__a22o_1
XANTENNA__07361__B net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08596_ _02913_ _02936_ vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__nand2_1
XFILLER_35_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_132_Left_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07547_ _02369_ _02370_ _02382_ vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_81_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07478_ datapath.rf.registers\[28\]\[21\] net750 net691 datapath.rf.registers\[13\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__a22o_1
XANTENNA__08473__A net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09217_ net320 _04052_ vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout505_X net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11103__S net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09148_ net375 _03982_ _03627_ net378 vssd1 vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__a211oi_1
XFILLER_136_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09242__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09079_ _03868_ _03914_ vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__and2_1
X_11110_ net304 net1640 net428 vssd1 vssd1 vccd1 vccd1 _00165_ sky130_fd_sc_hd__mux2_1
X_12090_ screen.register.currentYbus\[30\] _05786_ net999 screen.register.currentXbus\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06129_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_141_Left_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold770 datapath.rf.registers\[9\]\[24\] vssd1 vssd1 vccd1 vccd1 net2118 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout874_X net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold781 datapath.rf.registers\[5\]\[11\] vssd1 vssd1 vccd1 vccd1 net2129 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_112_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold792 datapath.rf.registers\[31\]\[15\] vssd1 vssd1 vccd1 vccd1 net2140 sky130_fd_sc_hd__dlygate4sd3_1
X_11041_ net302 net1594 net432 vssd1 vssd1 vccd1 vccd1 _00101_ sky130_fd_sc_hd__mux2_1
XANTENNA__10243__A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13865__RESET_B net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07020__A2 _01854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12869__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12992_ net174 net2139 net480 vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__mux2_1
XANTENNA__08648__A _01935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input13_A DAT_I[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11943_ net134 _05992_ _05991_ vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__o21ai_1
XFILLER_91_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10863__A0 _04118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07271__B net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14662_ clknet_leaf_11_clk _01367_ net1083 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11874_ net135 _05946_ _05945_ vssd1 vssd1 vccd1 vccd1 _00699_ sky130_fd_sc_hd__o21ai_1
X_13613_ clknet_leaf_132_clk _00423_ net1112 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10825_ _01446_ net655 _05580_ _05581_ vssd1 vssd1 vccd1 vccd1 _05582_ sky130_fd_sc_hd__o22a_2
XFILLER_32_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14593_ clknet_leaf_37_clk _01298_ net1138 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_119_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07087__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13544_ clknet_leaf_64_clk _00354_ net1235 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_41_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09481__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10756_ _01461_ net654 _05522_ vssd1 vssd1 vccd1 vccd1 _05523_ sky130_fd_sc_hd__o21a_1
X_13475_ clknet_leaf_118_clk _00285_ net1192 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10687_ _05433_ _05464_ _05503_ _05502_ _05501_ vssd1 vssd1 vccd1 vccd1 _05504_ sky130_fd_sc_hd__o32a_1
XANTENNA__11013__S net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12426_ net1394 net130 _06360_ vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__a21o_1
XANTENNA__09233__A0 _02312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12357_ _05002_ net306 _06321_ _06253_ _05667_ vssd1 vssd1 vccd1 vccd1 _06322_ sky130_fd_sc_hd__a32o_1
XFILLER_142_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07795__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11308_ _05696_ _05725_ vssd1 vssd1 vccd1 vccd1 _05726_ sky130_fd_sc_hd__nor2_4
X_12288_ net222 _05555_ _06271_ net891 vssd1 vssd1 vccd1 vccd1 _06272_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_52_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09536__A1 _02805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14027_ clknet_leaf_80_clk _00796_ net1257 vssd1 vssd1 vccd1 vccd1 datapath.PC\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_141_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11239_ net169 net2345 net527 vssd1 vssd1 vccd1 vccd1 _00289_ sky130_fd_sc_hd__mux2_1
XFILLER_68_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07011__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12779__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06780_ net1030 _01616_ vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__nor2_1
XFILLER_67_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10299__S net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08511__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08450_ datapath.rf.registers\[1\]\[2\] net764 net741 datapath.rf.registers\[16\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__a22o_1
X_07401_ _02225_ _02228_ _02229_ _02236_ vssd1 vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__or4_1
X_08381_ datapath.rf.registers\[1\]\[3\] net765 net697 datapath.rf.registers\[8\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03217_ sky130_fd_sc_hd__a22o_1
X_07332_ _02161_ _02163_ _02165_ _02167_ vssd1 vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_63_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06806__A _01438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07263_ datapath.rf.registers\[4\]\[25\] net959 net935 vssd1 vssd1 vccd1 vccd1 _02099_
+ sky130_fd_sc_hd__and3_1
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06838__A_N datapath.ru.latched_instruction\[29\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09002_ _03623_ _03837_ vssd1 vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__nand2_1
XFILLER_136_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07194_ datapath.rf.registers\[8\]\[27\] net695 net661 datapath.rf.registers\[5\]\[27\]
+ _02028_ vssd1 vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__a221o_1
XANTENNA__09224__B1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11826__D_N _05874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07786__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08983__C1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07250__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12262__B net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09904_ datapath.PC\[16\] _04738_ vssd1 vssd1 vccd1 vccd1 _04740_ sky130_fd_sc_hd__xor2_2
Xfanout502 net503 vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__buf_2
Xfanout513 _05735_ vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__buf_4
Xfanout524 _05723_ vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07538__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1207_A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout535 net537 vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__buf_4
XANTENNA__12531__B1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout546 _03759_ vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__clkbuf_4
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input5_A DAT_I[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07002__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout557 _03418_ vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__clkbuf_4
X_09835_ _03502_ _03507_ _03951_ _04024_ vssd1 vssd1 vccd1 vccd1 _04671_ sky130_fd_sc_hd__or4bb_1
Xfanout568 net569 vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__clkbuf_2
Xfanout579 net580 vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__buf_1
XANTENNA_fanout190_X net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09399__A2_N net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09766_ _04118_ _04586_ _04600_ vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__or3_1
XFILLER_101_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06978_ net963 net911 _01809_ vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__and3_1
XFILLER_67_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08717_ _03205_ _03228_ vssd1 vssd1 vccd1 vccd1 _03553_ sky130_fd_sc_hd__nand2_1
XANTENNA__07803__C net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout834_A net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09697_ _03436_ _04518_ vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_83_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08648_ _01935_ _01955_ vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__nand2_1
XFILLER_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10937__S net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08579_ datapath.rf.registers\[10\]\[0\] net708 _03412_ _03413_ _03414_ vssd1 vssd1
+ vccd1 vccd1 _03415_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12598__B1 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10610_ _05429_ vssd1 vssd1 vccd1 vccd1 _05430_ sky130_fd_sc_hd__inv_2
XFILLER_23_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11590_ net1273 net1274 _05802_ vssd1 vssd1 vccd1 vccd1 _05814_ sky130_fd_sc_hd__or3b_1
XANTENNA__12437__B net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10541_ datapath.multiplication_module.multiplier_i\[5\] datapath.multiplication_module.multiplier_i\[4\]
+ datapath.multiplication_module.multiplier_i\[7\] datapath.multiplication_module.multiplier_i\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05369_ sky130_fd_sc_hd__or4_1
XANTENNA__10238__A _04909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13260_ clknet_leaf_16_clk _00070_ net1108 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_98_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10472_ net1280 _01423_ _05301_ vssd1 vssd1 vccd1 vccd1 _05302_ sky130_fd_sc_hd__or3_2
XANTENNA_fanout991_X net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09215__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12211_ net2377 _06215_ net603 vssd1 vssd1 vccd1 vccd1 _06218_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08569__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09746__B _04580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13191_ net2219 vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__clkbuf_1
XFILLER_135_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10376__A2 net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12142_ _05771_ net601 _06174_ screen.counter.ct\[3\] vssd1 vssd1 vccd1 vccd1 _00738_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07241__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07266__B net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12073_ screen.register.currentXbus\[21\] _05769_ _05772_ screen.register.currentXbus\[29\]
+ _06112_ vssd1 vssd1 vccd1 vccd1 _06113_ sky130_fd_sc_hd__a221o_1
XANTENNA__07529__B1 _02363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11024_ net233 net2149 net538 vssd1 vssd1 vccd1 vccd1 _00086_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11516__B _05314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07713__C net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12975_ net254 net2389 net479 vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__mux2_1
XANTENNA__11008__S net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11926_ net2403 net160 vssd1 vssd1 vccd1 vccd1 _05981_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_142_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07701__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14645_ clknet_leaf_18_clk _01350_ net1108 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11857_ net2123 net163 vssd1 vssd1 vccd1 vccd1 _05935_ sky130_fd_sc_hd__nand2_1
XFILLER_32_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10808_ _05565_ _05566_ vssd1 vssd1 vccd1 vccd1 _05567_ sky130_fd_sc_hd__nor2_1
X_14576_ clknet_leaf_24_clk _01281_ net1157 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11788_ datapath.pc_module.i_ack1 datapath.i_ack vssd1 vssd1 vccd1 vccd1 _05900_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_45_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13527_ clknet_leaf_127_clk _00337_ net1211 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10739_ net1514 net568 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[25\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__11800__A2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07480__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13458_ clknet_leaf_30_clk _00268_ net1131 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06913__X _01749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12409_ _05966_ net157 vssd1 vssd1 vccd1 vccd1 _06352_ sky130_fd_sc_hd__nor2_1
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 SEL_O[0] sky130_fd_sc_hd__buf_2
X_13389_ clknet_leaf_124_clk _00199_ net1207 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13787__RESET_B net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput116 net116 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__buf_2
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07768__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09509__A1 _03149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07950_ datapath.rf.registers\[4\]\[11\] net959 net934 vssd1 vssd1 vccd1 vccd1 _02786_
+ sky130_fd_sc_hd__and3_1
X_06901_ net985 _01707_ net947 vssd1 vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__and3_4
X_07881_ datapath.rf.registers\[30\]\[13\] net759 net680 datapath.rf.registers\[6\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02717_ sky130_fd_sc_hd__a22o_1
X_09620_ net352 _04213_ _04218_ net360 vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__a211o_1
X_06832_ _01408_ net993 _01581_ _01667_ vssd1 vssd1 vccd1 vccd1 _01668_ sky130_fd_sc_hd__a31o_1
XFILLER_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08288__A _01604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09551_ net370 _03987_ _04386_ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__a21o_1
X_06763_ net1045 net1016 net994 net1029 datapath.ru.latched_instruction\[28\] vssd1
+ vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__a32oi_4
XFILLER_52_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08502_ datapath.rf.registers\[3\]\[1\] net914 _01797_ vssd1 vssd1 vccd1 vccd1 _03338_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_19_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06694_ datapath.ru.latched_instruction\[25\] net1046 vssd1 vssd1 vccd1 vccd1 _01533_
+ sky130_fd_sc_hd__xnor2_1
X_09482_ _02857_ net440 _04317_ net366 vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_65_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07299__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08433_ datapath.rf.registers\[4\]\[2\] net968 net911 _01809_ vssd1 vssd1 vccd1 vccd1
+ _03269_ sky130_fd_sc_hd__and4_1
XANTENNA__10757__S net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08775__C_N _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06807__Y _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13133__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout248_A net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08364_ datapath.rf.registers\[25\]\[3\] net844 net838 datapath.rf.registers\[26\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__a22o_1
XANTENNA__12257__B net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07315_ datapath.rf.registers\[20\]\[24\] net958 net923 vssd1 vssd1 vccd1 vccd1 _02151_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12972__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08295_ datapath.rf.registers\[13\]\[4\] net811 net805 datapath.rf.registers\[28\]\[4\]
+ _03130_ vssd1 vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout415_A _05726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1157_A net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07246_ datapath.rf.registers\[28\]\[26\] net750 net694 datapath.rf.registers\[8\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__a22o_1
XANTENNA__07471__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07177_ datapath.rf.registers\[22\]\[27\] net821 net815 datapath.rf.registers\[21\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02013_ sky130_fd_sc_hd__a22o_1
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07759__B1 _01772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout784_A net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout310 _06246_ vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__clkbuf_4
XFILLER_132_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout321 _03684_ vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__buf_1
Xfanout332 _03619_ vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout343 _03677_ vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__clkbuf_2
Xfanout354 net355 vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__buf_2
Xfanout365 _03629_ vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08184__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout376 net378 vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__buf_2
XANTENNA__09920__A1 _01786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout387 net389 vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__buf_4
X_09818_ _01889_ _01935_ net445 vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__mux2_1
XFILLER_87_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout398 net401 vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06734__A1 _01441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07931__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09749_ _04178_ _04207_ _04583_ vssd1 vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__nor3_1
XFILLER_27_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout837_X net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12760_ net2211 net182 net403 vssd1 vssd1 vccd1 vccd1 _00982_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09684__B1 _03604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ net28 net1033 net1023 net1400 vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__o22a_1
XFILLER_15_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12691_ datapath.mulitply_result\[30\] datapath.multiplication_module.multiplicand_i\[30\]
+ vssd1 vssd1 vccd1 vccd1 _06523_ sky130_fd_sc_hd__or2_1
XANTENNA__13043__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14430_ clknet_leaf_150_clk _01135_ net1059 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11642_ _05783_ _05823_ _05819_ vssd1 vssd1 vccd1 vccd1 _05866_ sky130_fd_sc_hd__o21ai_1
XFILLER_42_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14361_ clknet_leaf_9_clk _01066_ net1072 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12882__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11573_ net1008 _05762_ _05796_ net1006 vssd1 vssd1 vccd1 vccd1 _05797_ sky130_fd_sc_hd__o22a_1
Xinput18 DAT_I[24] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11794__A1 _01500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13312_ clknet_leaf_135_clk _00122_ net1104 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput29 DAT_I[5] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
X_10524_ screen.counter.ct\[1\] net1278 net1276 vssd1 vssd1 vccd1 vccd1 _05354_ sky130_fd_sc_hd__nor3_1
XANTENNA__07462__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14292_ clknet_leaf_93_clk _00997_ net1217 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11498__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13243_ clknet_leaf_39_clk _00053_ net1145 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10455_ mmio.wishbone.curr_state\[2\] mmio.wishbone.curr_state\[1\] vssd1 vssd1 vccd1
+ vccd1 _05289_ sky130_fd_sc_hd__nor2_1
XFILLER_136_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07214__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13174_ net2568 vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10386_ net377 _04504_ _05221_ net330 vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__o211a_1
XFILLER_112_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12125_ screen.counter.ct\[11\] net1275 net1274 _06161_ vssd1 vssd1 vccd1 vccd1 _06162_
+ sky130_fd_sc_hd__nand4_2
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12056_ screen.register.currentYbus\[20\] _05773_ _05778_ screen.register.currentYbus\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06097_ sky130_fd_sc_hd__a22o_1
XANTENNA__08175__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11007_ net304 net1650 net541 vssd1 vssd1 vccd1 vccd1 _00069_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_144_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07922__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12958_ net181 net2622 net395 vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12274__A2 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11909_ _02542_ net657 vssd1 vssd1 vccd1 vccd1 _05970_ sky130_fd_sc_hd__nand2_1
XFILLER_33_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12889_ net193 net2350 net398 vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__mux2_1
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14628_ clknet_leaf_18_clk _01333_ net1109 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14559_ clknet_leaf_13_clk _01264_ net1077 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12792__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07100_ datapath.rf.registers\[24\]\[29\] net767 net703 datapath.rf.registers\[9\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__a22o_1
XANTENNA__07989__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08080_ datapath.rf.registers\[30\]\[9\] net760 net752 datapath.rf.registers\[28\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02916_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_155_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07031_ datapath.rf.registers\[12\]\[30\] net955 net920 vssd1 vssd1 vccd1 vccd1 _01867_
+ sky130_fd_sc_hd__and3_1
XANTENNA__11201__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07205__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08982_ net337 _03816_ _03817_ vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__o21ai_2
XFILLER_103_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_143_Right_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07933_ datapath.rf.registers\[24\]\[12\] net769 net757 datapath.rf.registers\[12\]\[12\]
+ _02767_ vssd1 vssd1 vccd1 vccd1 _02769_ sky130_fd_sc_hd__a221o_1
XANTENNA__08166__B1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09902__A1 _01656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout198_A _05653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13128__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07864_ datapath.rf.registers\[10\]\[13\] net880 net827 datapath.rf.registers\[12\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__a22o_1
XFILLER_69_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09603_ _02857_ net440 _04317_ net362 vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__a211o_1
X_06815_ _01469_ net1002 net1018 net1027 datapath.ru.latched_instruction\[19\] vssd1
+ vssd1 vccd1 vccd1 _01651_ sky130_fd_sc_hd__a32o_1
XFILLER_95_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12967__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07795_ datapath.rf.registers\[19\]\[15\] net731 net680 datapath.rf.registers\[6\]\[15\]
+ _02630_ vssd1 vssd1 vccd1 vccd1 _02631_ sky130_fd_sc_hd__a221oi_1
XANTENNA__10060__B net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09534_ _02705_ _02751_ net441 vssd1 vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__mux2_1
X_06746_ _01461_ net1005 net1021 net1027 datapath.ru.latched_instruction\[3\] vssd1
+ vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__a32o_2
XANTENNA__12265__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11443__Y _05733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09465_ _03423_ _03554_ vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__xor2_1
X_06677_ datapath.ru.latched_instruction\[14\] _01513_ _01515_ vssd1 vssd1 vccd1 vccd1
+ _01516_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout532_A net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12268__A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08416_ datapath.rf.registers\[3\]\[2\] net803 net798 datapath.rf.registers\[29\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__a22o_1
XANTENNA__12017__A2 _05786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09396_ net328 _03988_ _04231_ net380 vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__a211o_1
XANTENNA__07692__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08347_ datapath.rf.registers\[5\]\[3\] net948 net936 vssd1 vssd1 vccd1 vccd1 _03183_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout418_X net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11900__A _02680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07444__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08278_ _03112_ _03113_ vssd1 vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_78_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07229_ datapath.rf.registers\[26\]\[26\] net836 net801 datapath.rf.registers\[3\]\[26\]
+ _02064_ vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__a221o_1
XFILLER_152_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11111__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10240_ _04841_ _05075_ vssd1 vssd1 vccd1 vccd1 _05076_ sky130_fd_sc_hd__nor2_1
XFILLER_145_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout787_X net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10171_ net228 _05001_ _05002_ _05006_ net1255 vssd1 vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__o221a_1
XANTENNA__10950__S net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1105 net1110 vssd1 vssd1 vccd1 vccd1 net1105 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_110_Right_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07825__A _02660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1116 net1119 vssd1 vssd1 vccd1 vccd1 net1116 sky130_fd_sc_hd__clkbuf_4
Xfanout1127 net1130 vssd1 vssd1 vccd1 vccd1 net1127 sky130_fd_sc_hd__clkbuf_4
Xfanout140 net142 vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__buf_2
Xfanout1138 net1139 vssd1 vssd1 vccd1 vccd1 net1138 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout954_X net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1149 net1151 vssd1 vssd1 vccd1 vccd1 net1149 sky130_fd_sc_hd__clkbuf_4
Xfanout151 _05886_ vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__buf_2
XANTENNA__08157__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout162 _05933_ vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__buf_2
XFILLER_59_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13038__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13930_ clknet_leaf_110_clk _00708_ net1201 vssd1 vssd1 vccd1 vccd1 screen.register.currentYbus\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout173 _05684_ vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_109_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout184 _05677_ vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__buf_1
XFILLER_86_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout195 _05659_ vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13861_ clknet_leaf_70_clk _00665_ net1244 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12877__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07263__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12812_ net1966 net249 net490 vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13792_ clknet_leaf_75_clk _00601_ net1242 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_70_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12743_ net1888 net264 net403 vssd1 vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__mux2_1
XFILLER_31_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12674_ datapath.mulitply_result\[27\] datapath.multiplication_module.multiplicand_i\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06509_ sky130_fd_sc_hd__nor2_1
XANTENNA__07683__A2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08943__X _03779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14413_ clknet_leaf_124_clk _01118_ net1207 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11625_ _05848_ vssd1 vssd1 vccd1 vccd1 _05849_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_42_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_85_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14344_ clknet_leaf_65_clk _01049_ net1238 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_155_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11556_ _05292_ _05754_ vssd1 vssd1 vccd1 vccd1 _05780_ sky130_fd_sc_hd__or2_2
XANTENNA__07435__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06904__A net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08391__A _03226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10507_ net1280 net1275 net1271 _05336_ vssd1 vssd1 vccd1 vccd1 _05337_ sky130_fd_sc_hd__a31o_1
X_14275_ clknet_leaf_119_clk _00980_ net1191 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11487_ net274 net2419 net512 vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__mux2_1
XFILLER_155_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11021__S net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13226_ clknet_leaf_58_clk _00036_ net1167 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10438_ datapath.PC\[3\] _01702_ vssd1 vssd1 vccd1 vccd1 _05274_ sky130_fd_sc_hd__nand2_1
XFILLER_152_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13157_ net1943 net183 net382 vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__mux2_1
X_10369_ net891 _04395_ vssd1 vssd1 vccd1 vccd1 _05205_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_143_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12108_ screen.counter.currentCt\[5\] screen.counter.currentCt\[4\] screen.counter.currentCt\[7\]
+ screen.counter.currentCt\[6\] vssd1 vssd1 vccd1 vccd1 _06145_ sky130_fd_sc_hd__or4_1
X_13088_ net2173 net194 net386 vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__mux2_1
XFILLER_112_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_23_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07454__B net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12039_ screen.register.currentXbus\[11\] _05768_ _05769_ screen.register.currentXbus\[19\]
+ _06080_ vssd1 vssd1 vccd1 vccd1 _06081_ sky130_fd_sc_hd__a221o_1
XFILLER_78_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12787__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_1_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_1_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08837__Y _03673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06600_ _01412_ _01438_ vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_0_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07580_ _02405_ _02406_ _02415_ vssd1 vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__or3b_1
XANTENNA__06638__X _01477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_38_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09014__X _03850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09250_ _03452_ _04085_ vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07674__A2 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08201_ datapath.rf.registers\[5\]\[6\] net945 net931 vssd1 vssd1 vccd1 vccd1 _03037_
+ sky130_fd_sc_hd__and3_1
XFILLER_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09181_ _03810_ _03813_ net448 vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__mux2_1
XANTENNA__11758__B2 _02487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08132_ datapath.rf.registers\[9\]\[8\] net705 net670 datapath.rf.registers\[21\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02968_ sky130_fd_sc_hd__a22o_1
XANTENNA__07426__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08063_ datapath.rf.registers\[2\]\[9\] net889 _02883_ _02884_ _02894_ vssd1 vssd1
+ vccd1 vccd1 _02899_ sky130_fd_sc_hd__a2111o_1
XFILLER_128_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07014_ datapath.rf.registers\[11\]\[31\] net711 net707 datapath.rf.registers\[10\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__a22o_1
XFILLER_108_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08387__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1022_A _01435_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10194__B1 net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08965_ _02856_ _02912_ net447 vssd1 vssd1 vccd1 vccd1 _03801_ sky130_fd_sc_hd__mux2_1
XFILLER_88_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout482_A _06554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08139__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07364__B net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07916_ datapath.rf.registers\[8\]\[12\] net695 net665 datapath.rf.registers\[15\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__a22o_1
XANTENNA__09887__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08896_ net469 _03480_ _03727_ _03731_ vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__a31o_1
XFILLER_57_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07847_ _02661_ _02681_ vssd1 vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout747_A net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07778_ datapath.rf.registers\[11\]\[15\] net711 net665 datapath.rf.registers\[15\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02614_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_88_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09517_ _02804_ _02856_ net452 vssd1 vssd1 vccd1 vccd1 _04353_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06729_ net1005 net1021 vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout535_X net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09448_ net356 _04106_ _04283_ net346 vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__a211o_1
XFILLER_24_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout702_X net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09379_ net552 net548 _02660_ vssd1 vssd1 vccd1 vccd1 _04215_ sky130_fd_sc_hd__a21o_1
XANTENNA__10945__S net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08923__B net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11749__B2 _02934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11410_ net209 net2328 net517 vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__mux2_1
XANTENNA__07417__A2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12390_ net1528 net133 _06342_ vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__a21o_1
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10421__A1 _03321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11341_ _05690_ _05692_ vssd1 vssd1 vccd1 vccd1 _05727_ sky130_fd_sc_hd__or2_1
XANTENNA__08090__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14060_ clknet_leaf_121_clk _00827_ net1199 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11272_ net170 net2288 net418 vssd1 vssd1 vccd1 vccd1 _00321_ sky130_fd_sc_hd__mux2_1
XANTENNA__08378__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13011_ net1930 net243 net391 vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__mux2_1
XANTENNA__09575__C1 _03614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10223_ _04893_ _04898_ vssd1 vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_18_Left_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10185__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10154_ _03745_ _04989_ net1040 vssd1 vssd1 vccd1 vccd1 _04990_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07274__B net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold7 keypad.debounce.debounce\[10\] vssd1 vssd1 vccd1 vccd1 net1355 sky130_fd_sc_hd__dlygate4sd3_1
X_10085_ net1265 datapath.PC\[23\] net1264 _03746_ datapath.PC\[25\] vssd1 vssd1 vccd1
+ vccd1 _04921_ sky130_fd_sc_hd__o41a_1
X_13913_ clknet_leaf_43_clk net1365 net1150 vssd1 vssd1 vccd1 vccd1 keypad.debounce.debounce\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_13844_ clknet_leaf_115_clk _00653_ net1189 vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__dfrtp_1
XFILLER_74_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_27_Left_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13775_ clknet_leaf_85_clk _00584_ net1258 vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__dfrtp_1
X_10987_ net1812 net218 net435 vssd1 vssd1 vccd1 vccd1 _00052_ sky130_fd_sc_hd__mux2_1
XANTENNA__08302__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11016__S net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12726_ columns.count\[8\] _06541_ columns.count\[9\] vssd1 vssd1 vccd1 vccd1 _06547_
+ sky130_fd_sc_hd__a21o_1
XFILLER_149_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_139_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12657_ _06486_ _06494_ vssd1 vssd1 vccd1 vccd1 _06495_ sky130_fd_sc_hd__or2_1
XANTENNA__08833__B _01614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07289__X _02125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11608_ _05782_ _05786_ _05826_ _05831_ vssd1 vssd1 vccd1 vccd1 _05832_ sky130_fd_sc_hd__or4_1
X_12588_ datapath.mulitply_result\[13\] datapath.multiplication_module.multiplicand_i\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06437_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_152_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14327_ clknet_leaf_130_clk _01032_ net1113 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_152_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11539_ screen.counter.ct\[2\] screen.counter.ct\[3\] vssd1 vssd1 vccd1 vccd1 _05763_
+ sky130_fd_sc_hd__nand2b_2
XANTENNA__07449__B _02284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08081__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold407 datapath.rf.registers\[14\]\[30\] vssd1 vssd1 vccd1 vccd1 net1755 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold418 datapath.rf.registers\[28\]\[11\] vssd1 vssd1 vccd1 vccd1 net1766 sky130_fd_sc_hd__dlygate4sd3_1
Xhold429 datapath.rf.registers\[12\]\[24\] vssd1 vssd1 vccd1 vccd1 net1777 sky130_fd_sc_hd__dlygate4sd3_1
X_14258_ clknet_leaf_30_clk _00963_ net1124 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_36_Left_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08369__B1 _03203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13209_ clknet_leaf_29_clk _00019_ net1131 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_14189_ clknet_leaf_91_clk datapath.multiplication_module.multiplicand_i_n\[0\] net1241
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_112_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout909 _01792_ vssd1 vssd1 vccd1 vccd1 net909 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07041__B1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1107 datapath.rf.registers\[16\]\[5\] vssd1 vssd1 vccd1 vccd1 net2455 sky130_fd_sc_hd__dlygate4sd3_1
X_08750_ _03502_ _03504_ _03585_ vssd1 vssd1 vccd1 vccd1 _03586_ sky130_fd_sc_hd__and3_1
Xhold1118 datapath.rf.registers\[24\]\[24\] vssd1 vssd1 vccd1 vccd1 net2466 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1129 datapath.rf.registers\[29\]\[0\] vssd1 vssd1 vccd1 vccd1 net2477 sky130_fd_sc_hd__dlygate4sd3_1
X_07701_ datapath.rf.registers\[17\]\[17\] net748 net724 datapath.rf.registers\[18\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__a22o_1
X_08681_ _03516_ vssd1 vssd1 vccd1 vccd1 _03517_ sky130_fd_sc_hd__inv_2
XANTENNA__11676__B1 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07632_ datapath.rf.registers\[3\]\[18\] net770 net691 datapath.rf.registers\[13\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__a22o_1
XFILLER_66_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07895__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07563_ datapath.rf.registers\[22\]\[19\] net952 net924 vssd1 vssd1 vccd1 vccd1 _02399_
+ sky130_fd_sc_hd__and3_1
X_09302_ net347 _04135_ net574 vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_24_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07647__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07494_ _02317_ _02318_ _02328_ _02329_ vssd1 vssd1 vccd1 vccd1 _02330_ sky130_fd_sc_hd__or4_1
XANTENNA__08583__X _03419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06855__B1 _01586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09233_ _02312_ _02365_ net453 vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__mux2_1
XFILLER_139_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13141__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09164_ net357 _03998_ _03999_ _03991_ vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__o31a_1
XANTENNA__08462__C _03294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08115_ datapath.rf.registers\[9\]\[8\] net886 net828 datapath.rf.registers\[12\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02951_ sky130_fd_sc_hd__a22o_1
XANTENNA__12980__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07359__B net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09095_ _03774_ _03930_ net354 vssd1 vssd1 vccd1 vccd1 _03931_ sky130_fd_sc_hd__mux2_1
XANTENNA__08072__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08046_ datapath.rf.registers\[15\]\[9\] net986 net915 vssd1 vssd1 vccd1 vccd1 _02882_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07280__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07078__C net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold930 datapath.rf.registers\[1\]\[28\] vssd1 vssd1 vccd1 vccd1 net2278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold941 datapath.rf.registers\[21\]\[26\] vssd1 vssd1 vccd1 vccd1 net2289 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold952 datapath.rf.registers\[1\]\[12\] vssd1 vssd1 vccd1 vccd1 net2300 sky130_fd_sc_hd__dlygate4sd3_1
Xhold963 datapath.rf.registers\[7\]\[27\] vssd1 vssd1 vccd1 vccd1 net2311 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold974 datapath.rf.registers\[18\]\[0\] vssd1 vssd1 vccd1 vccd1 net2322 sky130_fd_sc_hd__dlygate4sd3_1
Xhold985 datapath.rf.registers\[19\]\[7\] vssd1 vssd1 vccd1 vccd1 net2333 sky130_fd_sc_hd__dlygate4sd3_1
Xhold996 datapath.rf.registers\[0\]\[0\] vssd1 vssd1 vccd1 vccd1 net2344 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11609__B net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09997_ _04818_ _04832_ vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__xor2_1
XFILLER_131_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout864_A _01726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout485_X net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09309__C1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08948_ _02070_ _02126_ net445 vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__mux2_1
XANTENNA__14018__RESET_B net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08879_ _03707_ _03714_ net320 vssd1 vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__mux2_1
X_10910_ net1263 _05647_ vssd1 vssd1 vccd1 vccd1 _05654_ sky130_fd_sc_hd__and2_1
X_11890_ screen.register.currentYbus\[11\] net162 vssd1 vssd1 vccd1 vccd1 _05957_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__07886__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10841_ _05593_ _05594_ vssd1 vssd1 vccd1 vccd1 _05595_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout917_X net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13560_ clknet_leaf_4_clk _00370_ net1070 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[12\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10772_ net296 net2271 net545 vssd1 vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__mux2_1
XANTENNA__07638__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09493__D1 _03600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12511_ datapath.multiplication_module.multiplier_i\[0\] datapath.mulitply_result\[0\]
+ datapath.multiplication_module.multiplicand_i\[0\] net573 vssd1 vssd1 vccd1 vccd1
+ _06373_ sky130_fd_sc_hd__a31o_1
XANTENNA__09749__B _04207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13491_ clknet_leaf_33_clk _00301_ net1129 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13051__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12442_ net1424 net130 _06368_ vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__a21o_1
XFILLER_8_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12890__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12373_ _05242_ _05267_ net634 vssd1 vssd1 vccd1 vccd1 _06333_ sky130_fd_sc_hd__mux2_1
XANTENNA__07269__B net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08063__A2 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14112_ clknet_leaf_99_clk net1373 net1229 vssd1 vssd1 vccd1 vccd1 screen.register.xFill3
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11324_ net2082 net248 net415 vssd1 vssd1 vccd1 vccd1 _00369_ sky130_fd_sc_hd__mux2_1
XFILLER_141_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14043_ clknet_leaf_68_clk _00812_ net1245 vssd1 vssd1 vccd1 vccd1 datapath.PC\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11255_ net253 net2473 net419 vssd1 vssd1 vccd1 vccd1 _00304_ sky130_fd_sc_hd__mux2_1
XANTENNA__06901__B _01707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10206_ datapath.PC\[18\] _04600_ net469 vssd1 vssd1 vccd1 vccd1 _05042_ sky130_fd_sc_hd__mux2_1
X_11186_ net262 net2405 net423 vssd1 vssd1 vccd1 vccd1 _00238_ sky130_fd_sc_hd__mux2_1
XANTENNA__14441__RESET_B net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10137_ _04957_ _04971_ _04604_ vssd1 vssd1 vccd1 vccd1 _04973_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09315__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10068_ _01418_ _01593_ _01784_ _04900_ _04901_ vssd1 vssd1 vccd1 vccd1 _04904_ sky130_fd_sc_hd__o32a_1
XFILLER_85_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08523__B1 _03324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10330__B1 net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07877__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13827_ clknet_leaf_116_clk _00636_ net1187 vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__dfrtp_1
XFILLER_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13758_ clknet_leaf_76_clk _00567_ net1249 vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__dfrtp_1
XFILLER_44_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12709_ _05892_ _06530_ _06534_ net1378 vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__o22a_1
X_13689_ clknet_leaf_11_clk _00499_ net1081 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08563__B net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09787__C1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_44_Left_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold204 datapath.rf.registers\[7\]\[22\] vssd1 vssd1 vccd1 vccd1 net1552 sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 datapath.rf.registers\[27\]\[1\] vssd1 vssd1 vccd1 vccd1 net1563 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold226 datapath.rf.registers\[20\]\[26\] vssd1 vssd1 vccd1 vccd1 net1574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 datapath.rf.registers\[27\]\[0\] vssd1 vssd1 vccd1 vccd1 net1585 sky130_fd_sc_hd__dlygate4sd3_1
X_09920_ _01786_ _04754_ _04755_ datapath.PC\[11\] vssd1 vssd1 vccd1 vccd1 _04756_
+ sky130_fd_sc_hd__o31a_1
XANTENNA__12138__B2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold248 datapath.rf.registers\[3\]\[8\] vssd1 vssd1 vccd1 vccd1 net1596 sky130_fd_sc_hd__dlygate4sd3_1
Xhold259 datapath.rf.registers\[15\]\[20\] vssd1 vssd1 vccd1 vccd1 net1607 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_125_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07014__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout706 net709 vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__clkbuf_8
Xfanout717 _01815_ vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__clkbuf_4
X_09851_ _02442_ _02490_ vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__nand2_1
Xfanout728 _01812_ vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__buf_4
Xfanout739 net741 vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__clkbuf_4
X_08802_ _01603_ _03600_ vssd1 vssd1 vccd1 vccd1 _03638_ sky130_fd_sc_hd__or2_1
XFILLER_85_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09782_ net321 _04617_ vssd1 vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06994_ net968 _01820_ vssd1 vssd1 vccd1 vccd1 _01830_ sky130_fd_sc_hd__and2_1
XFILLER_105_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08733_ _03536_ _03537_ _03567_ _03534_ vssd1 vssd1 vccd1 vccd1 _03569_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_53_Left_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13136__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout278_A _05554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10949__A2_N _05686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08664_ _02284_ net563 vssd1 vssd1 vccd1 vccd1 _03500_ sky130_fd_sc_hd__and2b_1
XFILLER_38_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07615_ datapath.rf.registers\[8\]\[18\] net876 net801 datapath.rf.registers\[3\]\[18\]
+ _02450_ vssd1 vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_68_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08457__C net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12975__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07361__C net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08595_ _03032_ _03429_ _03033_ _02937_ _02984_ vssd1 vssd1 vccd1 vccd1 _03431_ sky130_fd_sc_hd__a2111o_1
XFILLER_121_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07546_ _02374_ _02375_ _02380_ _02381_ vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__or4_1
XFILLER_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07477_ datapath.rf.registers\[20\]\[21\] net718 net660 datapath.rf.registers\[5\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__a22o_1
XANTENNA__08293__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout612_A net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09216_ _03905_ _03907_ net340 vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__mux2_1
X_09147_ net375 _03982_ _03627_ vssd1 vssd1 vccd1 vccd1 _03983_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout400_X net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09242__A1 _02364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09078_ _03869_ _03870_ _03913_ vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout981_A net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08029_ datapath.rf.registers\[19\]\[10\] net732 _02863_ _02864_ net788 vssd1 vssd1
+ vccd1 vccd1 _02865_ sky130_fd_sc_hd__a2111o_1
Xhold760 datapath.rf.registers\[11\]\[25\] vssd1 vssd1 vccd1 vccd1 net2108 sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 datapath.rf.registers\[13\]\[23\] vssd1 vssd1 vccd1 vccd1 net2119 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07005__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold782 datapath.rf.registers\[10\]\[8\] vssd1 vssd1 vccd1 vccd1 net2130 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_112_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11040_ net288 net1774 net433 vssd1 vssd1 vccd1 vccd1 _00100_ sky130_fd_sc_hd__mux2_1
Xhold793 datapath.rf.registers\[22\]\[30\] vssd1 vssd1 vccd1 vccd1 net2141 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout867_X net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10811__X _05570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08488__X _03324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12991_ net181 net2536 net479 vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__mux2_1
XFILLER_92_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13046__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12301__B2 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11942_ _02001_ screen.counter.ack vssd1 vssd1 vccd1 vccd1 _05992_ sky130_fd_sc_hd__or2_1
XANTENNA__07859__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14661_ clknet_leaf_116_clk _01366_ net1188 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07271__C net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11873_ _03123_ net657 vssd1 vssd1 vccd1 vccd1 _05946_ sky130_fd_sc_hd__nand2_1
XANTENNA__12885__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13612_ clknet_leaf_18_clk _00422_ net1108 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10824_ datapath.mulitply_result\[13\] net598 net621 vssd1 vssd1 vccd1 vccd1 _05581_
+ sky130_fd_sc_hd__a21o_1
X_14592_ clknet_leaf_135_clk _01297_ net1102 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_13543_ clknet_leaf_142_clk _00353_ net1087 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_41_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10755_ datapath.mulitply_result\[3\] net600 _05520_ _05521_ net621 vssd1 vssd1 vccd1
+ vccd1 _05522_ sky130_fd_sc_hd__a221o_1
XANTENNA__08284__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07492__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13474_ clknet_leaf_152_clk _00284_ net1054 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10686_ button\[3\] _01435_ vssd1 vssd1 vccd1 vccd1 _05503_ sky130_fd_sc_hd__and2_1
XFILLER_9_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12425_ _05982_ net156 vssd1 vssd1 vccd1 vccd1 _06360_ sky130_fd_sc_hd__nor2_1
XFILLER_138_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09233__A1 _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07244__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09784__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12356_ net893 _04829_ vssd1 vssd1 vccd1 vccd1 _06321_ sky130_fd_sc_hd__nand2_1
XFILLER_153_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06912__A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11307_ _05692_ _05724_ vssd1 vssd1 vccd1 vccd1 _05725_ sky130_fd_sc_hd__or2_1
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12287_ net222 _04850_ vssd1 vssd1 vccd1 vccd1 _06271_ sky130_fd_sc_hd__nand2_1
XANTENNA__06765__A1_N datapath.ru.latched_instruction\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14026_ clknet_leaf_80_clk _00795_ net1254 vssd1 vssd1 vccd1 vccd1 datapath.PC\[16\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_113_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09536__A2 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11238_ net173 net2302 net528 vssd1 vssd1 vccd1 vccd1 _00288_ sky130_fd_sc_hd__mux2_1
XFILLER_110_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11169_ net178 net2253 net533 vssd1 vssd1 vccd1 vccd1 _00222_ sky130_fd_sc_hd__mux2_1
XANTENNA__08839__A _01637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08558__B net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12795__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07180__C1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07400_ _02230_ _02232_ _02233_ _02235_ vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__or4_1
XANTENNA__12056__B1 _05778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08380_ _03209_ _03211_ _03213_ _03215_ vssd1 vssd1 vccd1 vccd1 _03216_ sky130_fd_sc_hd__or4_2
X_07331_ datapath.rf.registers\[17\]\[24\] net849 net846 datapath.rf.registers\[1\]\[24\]
+ _02166_ vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__a221o_1
XFILLER_32_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08275__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_0_clk_X clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11204__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07483__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07262_ datapath.rf.registers\[27\]\[25\] net978 net938 vssd1 vssd1 vccd1 vccd1 _02098_
+ sky130_fd_sc_hd__and3_1
X_09001_ net374 _03836_ _03833_ net328 vssd1 vssd1 vccd1 vccd1 _03837_ sky130_fd_sc_hd__a211o_1
X_07193_ datapath.rf.registers\[25\]\[27\] net727 net719 datapath.rf.registers\[20\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02029_ sky130_fd_sc_hd__a22o_1
XANTENNA__08027__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07235__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08983__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09903_ datapath.PC\[16\] _04738_ vssd1 vssd1 vccd1 vccd1 _04739_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_4_9_0_clk_X clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout503 net505 vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__buf_2
Xfanout514 _05731_ vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__clkbuf_8
Xfanout525 _05723_ vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__clkbuf_4
XFILLER_101_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout395_A _06555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout536 net537 vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__buf_6
Xfanout547 _03656_ vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__buf_2
X_09834_ _03497_ _04669_ _03866_ _01910_ vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__nand4b_1
XANTENNA_fanout1102_A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout558 _03383_ vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__clkbuf_4
Xfanout569 _05368_ vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07653__A _02467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09765_ _04586_ _04600_ vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__nor2_1
X_06977_ net910 net907 vssd1 vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__and2_1
XFILLER_27_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08716_ _03549_ _03550_ _03545_ vssd1 vssd1 vccd1 vccd1 _03552_ sky130_fd_sc_hd__a21o_1
XFILLER_39_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09696_ net324 _03909_ vssd1 vssd1 vccd1 vccd1 _04532_ sky130_fd_sc_hd__or2_1
XFILLER_27_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08647_ _01935_ _01955_ vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout1092_X net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout827_A net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11903__A _02633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08578_ datapath.rf.registers\[11\]\[0\] net969 _01816_ vssd1 vssd1 vccd1 vccd1 _03414_
+ sky130_fd_sc_hd__and3_1
XFILLER_25_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07529_ datapath.rf.registers\[0\]\[20\] net870 _02363_ vssd1 vssd1 vccd1 vccd1 _02365_
+ sky130_fd_sc_hd__o21ai_4
XANTENNA__09463__A1 _03604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10519__A _05335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout615_X net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11114__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10073__A2 net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10540_ datapath.multiplication_module.mul_prev net615 vssd1 vssd1 vccd1 vccd1 _05368_
+ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_33_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08771__X _03607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10238__B _05073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10471_ net1278 net1279 net1277 _05300_ vssd1 vssd1 vccd1 vccd1 _05301_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_98_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12210_ screen.counter.currentCt\[7\] screen.counter.currentCt\[6\] _06214_ vssd1
+ vssd1 vccd1 vccd1 _06217_ sky130_fd_sc_hd__and3_1
XANTENNA__07226__B1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13190_ net1538 vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08974__A0 _03263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout984_X net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12141_ screen.counter.ct\[2\] _06175_ _06174_ vssd1 vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__o21a_1
XFILLER_150_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_756 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12072_ screen.register.currentXbus\[5\] net1000 _06018_ screen.register.currentYbus\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06112_ sky130_fd_sc_hd__a22o_1
Xhold590 datapath.rf.registers\[18\]\[4\] vssd1 vssd1 vccd1 vccd1 net1938 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07266__C net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11023_ net237 net2494 net540 vssd1 vssd1 vccd1 vccd1 _00085_ sky130_fd_sc_hd__mux2_1
XFILLER_150_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08659__A _02169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12974_ net262 net1816 net481 vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__mux2_1
Xhold1290 screen.counter.currentCt\[1\] vssd1 vssd1 vccd1 vccd1 net2638 sky130_fd_sc_hd__dlygate4sd3_1
X_11925_ net134 _05980_ _05979_ vssd1 vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_142_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14644_ clknet_leaf_20_clk _01349_ net1118 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11856_ _05074_ _05204_ _05284_ _05932_ vssd1 vssd1 vccd1 vccd1 _05934_ sky130_fd_sc_hd__or4_4
XANTENNA__08394__A _03204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10807_ datapath.PC\[11\] _05559_ vssd1 vssd1 vccd1 vccd1 _05566_ sky130_fd_sc_hd__nor2_1
X_14575_ clknet_leaf_36_clk _01280_ net1135 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11787_ datapath.ru.n_memwrite MemWrite net622 datapath.ru.n_memread vssd1 vssd1
+ vccd1 vccd1 _05899_ sky130_fd_sc_hd__a22o_1
XANTENNA__08257__A2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10429__A _03770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11024__S net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10738_ net1516 net568 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[24\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_31_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07465__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13526_ clknet_leaf_140_clk _00336_ net1096 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10863__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08009__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13457_ clknet_leaf_38_clk _00267_ net1141 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10669_ _05472_ _05486_ _05487_ _05447_ _01430_ vssd1 vssd1 vccd1 vccd1 _05488_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_124_Right_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12408_ net1415 net132 _06351_ vssd1 vssd1 vccd1 vccd1 _00828_ sky130_fd_sc_hd__a21o_1
XANTENNA__07217__B1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09459__A2_N net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13388_ clknet_leaf_15_clk _00198_ net1103 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 SEL_O[1] sky130_fd_sc_hd__buf_2
XFILLER_142_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08965__A0 _02856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput117 net117 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__buf_2
X_12339_ datapath.PC\[23\] _06308_ net306 vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__mux2_1
XFILLER_141_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_149_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14009_ clknet_leaf_75_clk _00000_ net1247 vssd1 vssd1 vccd1 vccd1 mmio.wishbone.curr_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_06900_ datapath.rf.registers\[11\]\[31\] net883 net849 datapath.rf.registers\[17\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__a22o_1
X_07880_ datapath.rf.registers\[22\]\[13\] net735 net695 datapath.rf.registers\[8\]\[13\]
+ _02715_ vssd1 vssd1 vccd1 vccd1 _02716_ sky130_fd_sc_hd__a221o_1
XANTENNA__13756__RESET_B net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06831_ datapath.ru.latched_instruction\[28\] net1045 net1014 net993 vssd1 vssd1
+ vccd1 vccd1 _01667_ sky130_fd_sc_hd__and4b_1
XANTENNA__10611__B _01435_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08288__B _01784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09550_ net363 _04063_ _04226_ net371 vssd1 vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__a211oi_1
XFILLER_110_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06762_ datapath.ru.latched_instruction\[27\] net1031 net994 _01597_ _01596_ vssd1
+ vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__a221oi_2
XFILLER_64_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08501_ datapath.rf.registers\[11\]\[1\] net970 _01816_ vssd1 vssd1 vccd1 vccd1 _03337_
+ sky130_fd_sc_hd__and3_1
X_09481_ net557 net576 net546 _02913_ vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_65_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06693_ net1289 net1283 mmio.memload_or_instruction\[25\] vssd1 vssd1 vccd1 vccd1
+ _01532_ sky130_fd_sc_hd__nor3b_1
XFILLER_24_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_19_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08496__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08432_ datapath.rf.registers\[11\]\[2\] net971 _01816_ vssd1 vssd1 vccd1 vccd1 _03268_
+ sky130_fd_sc_hd__and3_1
X_08363_ datapath.rf.registers\[24\]\[3\] net859 _03179_ _03193_ _03198_ vssd1 vssd1
+ vccd1 vccd1 _03199_ sky130_fd_sc_hd__a2111o_1
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout143_A net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07314_ datapath.rf.registers\[5\]\[24\] net946 net933 vssd1 vssd1 vccd1 vccd1 _02150_
+ sky130_fd_sc_hd__and3_1
X_08294_ datapath.rf.registers\[25\]\[4\] net841 net829 datapath.rf.registers\[14\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03130_ sky130_fd_sc_hd__a22o_1
XFILLER_20_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12472__A1_N net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07245_ _02079_ _02080_ vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__or2_1
XFILLER_149_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout310_A _06246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout408_A _05733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1052_A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07176_ _02009_ _02011_ vssd1 vssd1 vccd1 vccd1 _02012_ sky130_fd_sc_hd__or2_1
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10763__B1 _05527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07935__X _02771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout300 net301 vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__clkbuf_2
Xfanout311 _03620_ vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__buf_2
XANTENNA_fanout398_X net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout777_A _01796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout322 net323 vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__buf_2
Xfanout333 _05904_ vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__clkbuf_4
Xfanout344 _03676_ vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__buf_2
Xfanout355 _03649_ vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__clkbuf_2
Xfanout366 net369 vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__buf_2
XFILLER_87_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout377 _03621_ vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__buf_2
X_09817_ net348 _04220_ net575 vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__o21a_1
XFILLER_100_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout388 net389 vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__buf_6
Xfanout399 net401 vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__buf_4
XANTENNA_fanout565_X net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout944_A _01715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06734__A2 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11109__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09748_ _04207_ _04583_ vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__nor2_1
XANTENNA__09133__B1 _03770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout732_X net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09679_ net633 _04513_ _04514_ _03824_ vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_38_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08485__Y _03321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ net27 net1035 net1025 net1489 vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_124_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12690_ datapath.mulitply_result\[30\] datapath.multiplication_module.multiplicand_i\[30\]
+ vssd1 vssd1 vccd1 vccd1 _06522_ sky130_fd_sc_hd__nand2_1
XANTENNA__07695__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11641_ _05861_ _05864_ vssd1 vssd1 vccd1 vccd1 _05865_ sky130_fd_sc_hd__nand2_1
XANTENNA__09436__A1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07447__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14360_ clknet_leaf_7_clk _01065_ net1068 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[1\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11572_ _05293_ _05754_ _05753_ vssd1 vssd1 vccd1 vccd1 _05796_ sky130_fd_sc_hd__a21o_1
XANTENNA__11779__S _05894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13311_ clknet_leaf_12_clk _00121_ net1082 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput19 DAT_I[25] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
X_10523_ net1272 _05352_ vssd1 vssd1 vccd1 vccd1 _05353_ sky130_fd_sc_hd__nor2_1
X_14291_ clknet_leaf_64_clk _00996_ net1236 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[11\]
+ sky130_fd_sc_hd__dfrtp_2
X_13242_ clknet_leaf_2_clk _00052_ net1062 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10454_ net2547 _01419_ mmio.wishbone.curr_state\[0\] _05287_ vssd1 vssd1 vccd1 vccd1
+ _00001_ sky130_fd_sc_hd__a22o_1
XFILLER_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08947__A0 _01981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13173_ datapath.rf.registers\[0\]\[10\] vssd1 vssd1 vccd1 vccd1 _00995_ sky130_fd_sc_hd__clkbuf_1
X_10385_ net371 _04405_ _05220_ net329 vssd1 vssd1 vccd1 vccd1 _05221_ sky130_fd_sc_hd__a211o_1
XFILLER_151_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12124_ net1276 net1277 _05907_ _06154_ vssd1 vssd1 vccd1 vccd1 _06161_ sky130_fd_sc_hd__and4_1
XANTENNA__09773__A _01706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12055_ screen.register.currentXbus\[12\] net999 net997 screen.register.currentXbus\[20\]
+ vssd1 vssd1 vccd1 vccd1 _06096_ sky130_fd_sc_hd__a22o_1
XFILLER_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11006_ net287 net1734 net540 vssd1 vssd1 vccd1 vccd1 _00068_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_144_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11019__S net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08478__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12957_ net179 net2109 net396 vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__mux2_1
XANTENNA__09675__A1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06908__Y _01744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11908_ net2561 net162 vssd1 vssd1 vccd1 vccd1 _05969_ sky130_fd_sc_hd__nand2_1
XANTENNA__07686__B1 _02521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12888_ net198 net2521 net400 vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__mux2_1
X_14627_ clknet_leaf_139_clk _01332_ net1194 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11839_ _05914_ _05915_ _05917_ vssd1 vssd1 vccd1 vccd1 _05918_ sky130_fd_sc_hd__or3_1
XFILLER_20_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07438__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14558_ clknet_leaf_1_clk _01263_ net1062 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06924__X _01760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07989__A1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10442__C1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13509_ clknet_leaf_118_clk _00319_ net1189 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_14489_ clknet_leaf_31_clk _01194_ net1123 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_155_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07030_ datapath.rf.registers\[8\]\[30\] net955 _01712_ vssd1 vssd1 vccd1 vccd1 _01866_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_58_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08981_ net319 _03807_ vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__or2_1
XFILLER_142_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07932_ datapath.rf.registers\[31\]\[12\] net689 net681 datapath.rf.registers\[6\]\[12\]
+ _02761_ vssd1 vssd1 vccd1 vccd1 _02768_ sky130_fd_sc_hd__a221o_1
XFILLER_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07863_ datapath.rf.registers\[25\]\[13\] net843 net791 datapath.rf.registers\[18\]\[13\]
+ _02698_ vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__a221o_1
XFILLER_29_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06814_ _01469_ net1003 net1019 net1026 datapath.ru.latched_instruction\[19\] vssd1
+ vssd1 vccd1 vccd1 _01650_ sky130_fd_sc_hd__a32oi_2
X_09602_ _01609_ _04437_ _03770_ vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__o21a_1
XFILLER_56_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07794_ datapath.rf.registers\[26\]\[15\] net779 net727 datapath.rf.registers\[25\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02630_ sky130_fd_sc_hd__a22o_1
X_09533_ net643 _04366_ _04368_ vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__or3_1
X_06745_ _01582_ _01583_ vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__nand2_1
XFILLER_37_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08469__A2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout260_A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13144__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09464_ _04275_ _04299_ vssd1 vssd1 vccd1 vccd1 _04300_ sky130_fd_sc_hd__or2_1
X_06676_ net1287 net1282 datapath.ru.latched_instruction\[15\] mmio.memload_or_instruction\[15\]
+ vssd1 vssd1 vccd1 vccd1 _01515_ sky130_fd_sc_hd__or4b_1
XANTENNA__07141__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08415_ net875 _03248_ _03249_ _03250_ vssd1 vssd1 vccd1 vccd1 _03251_ sky130_fd_sc_hd__or4_1
XANTENNA__12983__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09395_ net328 _04230_ vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__nor2_1
XFILLER_11_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09418__B2 _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout525_A _05723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07429__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08346_ datapath.rf.registers\[22\]\[3\] net953 net926 vssd1 vssd1 vccd1 vccd1 _03182_
+ sky130_fd_sc_hd__and3_1
XANTENNA__11900__B net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08277_ datapath.rf.registers\[16\]\[5\] net739 net723 datapath.rf.registers\[18\]\[5\]
+ _03110_ vssd1 vssd1 vccd1 vccd1 _03113_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout313_X net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13458__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12284__A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07228_ datapath.rf.registers\[4\]\[26\] net864 net841 datapath.rf.registers\[25\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_95_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout894_A net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08929__A0 _01934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07159_ datapath.rf.registers\[1\]\[28\] net765 net717 datapath.rf.registers\[4\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1222_X net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10170_ net1043 _05003_ _05004_ _05005_ vssd1 vssd1 vccd1 vccd1 _05006_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout682_X net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1106 net1110 vssd1 vssd1 vccd1 vccd1 net1106 sky130_fd_sc_hd__clkbuf_4
XFILLER_121_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1117 net1119 vssd1 vssd1 vccd1 vccd1 net1117 sky130_fd_sc_hd__clkbuf_4
XFILLER_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout130 net132 vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__buf_2
Xfanout1128 net1130 vssd1 vssd1 vccd1 vccd1 net1128 sky130_fd_sc_hd__clkbuf_4
Xfanout141 net142 vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__buf_1
Xfanout1139 net1153 vssd1 vssd1 vccd1 vccd1 net1139 sky130_fd_sc_hd__clkbuf_2
Xfanout152 net155 vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__buf_2
Xfanout163 _05933_ vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__clkbuf_2
XFILLER_93_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout174 _05684_ vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_109_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout185 net188 vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout947_X net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout196 _05653_ vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__clkbuf_2
X_13860_ clknet_leaf_53_clk _00664_ net1180 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_28_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12811_ net1801 net251 net490 vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13791_ clknet_leaf_74_clk _00600_ net1247 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13054__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07560__B net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12742_ net2610 net269 net404 vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__mux2_1
XFILLER_42_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07132__A2 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_916 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12673_ datapath.mulitply_result\[27\] datapath.multiplication_module.multiplicand_i\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06508_ sky130_fd_sc_hd__and2_1
XFILLER_43_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12893__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11513__D _05335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11624_ _05358_ _05846_ vssd1 vssd1 vccd1 vccd1 _05848_ sky130_fd_sc_hd__or2_1
XFILLER_8_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14412_ clknet_leaf_17_clk _01117_ net1106 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09768__A _04023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08672__A _02419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14343_ clknet_leaf_137_clk _01048_ net1097 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11555_ _05292_ net1006 _05763_ vssd1 vssd1 vccd1 vccd1 _05779_ sky130_fd_sc_hd__nor3_1
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08093__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06904__B net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11302__S net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10506_ _05335_ vssd1 vssd1 vccd1 vccd1 _05336_ sky130_fd_sc_hd__inv_2
X_14274_ clknet_leaf_152_clk _00979_ net1056 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_21_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07840__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11486_ net279 net2291 net513 vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__mux2_1
Xwire586 _02749_ vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13225_ clknet_leaf_62_clk _00035_ net1165 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10437_ _04396_ _05272_ vssd1 vssd1 vccd1 vccd1 _05273_ sky130_fd_sc_hd__and2_1
XFILLER_124_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07199__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13156_ net1698 net178 net384 vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__mux2_1
X_10368_ _05085_ net180 net189 vssd1 vssd1 vccd1 vccd1 _05204_ sky130_fd_sc_hd__nand3_1
XANTENNA__06920__A net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12107_ _06144_ net1440 _06017_ vssd1 vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__mux2_1
XFILLER_151_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13087_ net2516 net197 net388 vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__mux2_1
XFILLER_97_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10299_ _05132_ _05134_ net224 vssd1 vssd1 vccd1 vccd1 _05135_ sky130_fd_sc_hd__mux2_1
X_12038_ screen.register.currentYbus\[11\] _06019_ _06078_ _06079_ vssd1 vssd1 vccd1
+ vccd1 _06080_ sky130_fd_sc_hd__a211o_1
XFILLER_66_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07454__C net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07371__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13989_ clknet_leaf_112_clk _00766_ net1219 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08200_ datapath.rf.registers\[29\]\[6\] net974 net917 vssd1 vssd1 vccd1 vccd1 _03036_
+ sky130_fd_sc_hd__and3_1
X_09180_ _03805_ _03809_ net448 vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__mux2_1
X_08131_ datapath.rf.registers\[3\]\[8\] net772 net765 datapath.rf.registers\[1\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02967_ sky130_fd_sc_hd__a22o_1
XANTENNA__08084__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11212__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08062_ datapath.rf.registers\[1\]\[9\] net847 net806 datapath.rf.registers\[28\]\[9\]
+ _02886_ vssd1 vssd1 vccd1 vccd1 _02898_ sky130_fd_sc_hd__a221o_1
XANTENNA__07831__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07629__C net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07013_ datapath.rf.registers\[12\]\[31\] net754 net664 datapath.rf.registers\[15\]\[31\]
+ _01848_ vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_73_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13139__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08964_ _02750_ _02804_ net447 vssd1 vssd1 vccd1 vccd1 _03800_ sky130_fd_sc_hd__mux2_1
XFILLER_69_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07915_ datapath.rf.registers\[0\]\[12\] net870 _02741_ net585 vssd1 vssd1 vccd1
+ vccd1 _02751_ sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12978__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07364__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08895_ datapath.PC\[31\] net468 net1038 vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout475_A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07846_ _02661_ _02681_ vssd1 vssd1 vccd1 vccd1 _02682_ sky130_fd_sc_hd__nor2_1
XANTENNA__07898__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07777_ _02612_ vssd1 vssd1 vccd1 vccd1 _02613_ sky130_fd_sc_hd__inv_2
XFILLER_37_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09516_ net457 _04349_ _04350_ vssd1 vssd1 vccd1 vccd1 _04352_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_104_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06728_ net1005 net1021 vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__and2_1
XANTENNA__07114__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09447_ net349 _04282_ _04277_ net359 vssd1 vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__o211a_1
X_06659_ net1287 net1282 mmio.memload_or_instruction\[29\] vssd1 vssd1 vccd1 vccd1
+ _01498_ sky130_fd_sc_hd__or3b_1
XANTENNA_fanout430_X net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout528_X net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09378_ _02612_ net554 net550 vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__or3_1
XFILLER_40_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11749__A2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08329_ datapath.rf.registers\[22\]\[4\] net735 net718 datapath.rf.registers\[20\]\[4\]
+ _03164_ vssd1 vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__a221o_1
XFILLER_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11122__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09875__X _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11340_ net1821 net168 net415 vssd1 vssd1 vccd1 vccd1 _00385_ sky130_fd_sc_hd__mux2_1
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout897_X net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11271_ net175 net1652 net420 vssd1 vssd1 vccd1 vccd1 _00320_ sky130_fd_sc_hd__mux2_1
XFILLER_106_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13010_ net1622 net247 net390 vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__mux2_1
X_10222_ net637 _05055_ _05057_ net226 vssd1 vssd1 vccd1 vccd1 _05058_ sky130_fd_sc_hd__a211o_1
XFILLER_152_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10185__A1 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13049__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10153_ datapath.PC\[20\] _03744_ vssd1 vssd1 vccd1 vccd1 _04989_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_7_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input36_A gpio_in[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10084_ datapath.PC\[25\] net1295 vssd1 vssd1 vccd1 vccd1 _04920_ sky130_fd_sc_hd__and2_1
XFILLER_48_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07274__C net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12888__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold8 keypad.debounce.debounce\[13\] vssd1 vssd1 vccd1 vccd1 net1356 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13912_ clknet_leaf_43_clk net1356 net1150 vssd1 vssd1 vccd1 vccd1 keypad.debounce.debounce\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08667__A _02312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13843_ clknet_leaf_76_clk _00652_ net1247 vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__dfrtp_1
XFILLER_62_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13774_ clknet_leaf_83_clk _00583_ net1260 vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__dfrtp_1
XFILLER_74_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10986_ net1785 net239 net436 vssd1 vssd1 vccd1 vccd1 _00051_ sky130_fd_sc_hd__mux2_1
XFILLER_90_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07105__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12725_ _01431_ _06538_ vssd1 vssd1 vccd1 vccd1 _06546_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_26_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12656_ _06481_ _06485_ _06487_ vssd1 vssd1 vccd1 vccd1 _06494_ sky130_fd_sc_hd__a21oi_1
X_11607_ _05302_ _05760_ _05784_ vssd1 vssd1 vccd1 vccd1 _05831_ sky130_fd_sc_hd__o21bai_1
XANTENNA__08066__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12587_ datapath.mulitply_result\[13\] datapath.multiplication_module.multiplicand_i\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06436_ sky130_fd_sc_hd__nand2_1
XFILLER_128_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11032__S net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14326_ clknet_leaf_137_clk _01031_ net1098 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07813__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11538_ _05749_ _05753_ vssd1 vssd1 vccd1 vccd1 _05762_ sky130_fd_sc_hd__or2_1
Xhold408 datapath.rf.registers\[9\]\[18\] vssd1 vssd1 vccd1 vccd1 net1756 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold419 datapath.rf.registers\[25\]\[4\] vssd1 vssd1 vccd1 vccd1 net1767 sky130_fd_sc_hd__dlygate4sd3_1
X_11469_ net2505 net197 net408 vssd1 vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__mux2_1
X_14257_ clknet_leaf_39_clk _00962_ net1142 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09945__B _03384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08369__A1 datapath.rf.registers\[0\]\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09566__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13208_ clknet_leaf_4_clk _00018_ net1069 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_14188_ clknet_leaf_69_clk net599 net1245 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.mul_prev
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_55_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13139_ net2427 net267 net384 vssd1 vssd1 vccd1 vccd1 _01380_ sky130_fd_sc_hd__mux2_1
XFILLER_112_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07592__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1108 datapath.rf.registers\[12\]\[3\] vssd1 vssd1 vccd1 vccd1 net2456 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12798__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1119 datapath.rf.registers\[11\]\[3\] vssd1 vssd1 vccd1 vccd1 net2467 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07700_ datapath.rf.registers\[30\]\[17\] net760 net677 datapath.rf.registers\[29\]\[17\]
+ _02535_ vssd1 vssd1 vccd1 vccd1 _02536_ sky130_fd_sc_hd__a221o_1
X_08680_ _02567_ _02588_ vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__nand2_1
XANTENNA__07344__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07631_ _02466_ vssd1 vssd1 vccd1 vccd1 _02467_ sky130_fd_sc_hd__inv_2
X_07562_ datapath.rf.registers\[6\]\[19\] net952 net934 vssd1 vssd1 vccd1 vccd1 _02398_
+ sky130_fd_sc_hd__and3_1
X_09301_ _03641_ _04136_ _04128_ vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__o21a_1
X_07493_ datapath.rf.registers\[12\]\[21\] net754 net738 datapath.rf.registers\[16\]\[21\]
+ _02327_ vssd1 vssd1 vccd1 vccd1 _02329_ sky130_fd_sc_hd__a221o_1
XFILLER_22_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09232_ net330 _04061_ _04067_ net311 vssd1 vssd1 vccd1 vccd1 _04068_ sky130_fd_sc_hd__a31oi_1
XANTENNA__09201__A net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09163_ net461 _03773_ _03992_ net351 vssd1 vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__o211a_1
XFILLER_30_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08114_ datapath.rf.registers\[25\]\[8\] net843 _02945_ _02949_ net875 vssd1 vssd1
+ vccd1 vccd1 _02950_ sky130_fd_sc_hd__a2111oi_1
X_09094_ _03928_ _03929_ net461 vssd1 vssd1 vccd1 vccd1 _03930_ sky130_fd_sc_hd__mux2_1
XANTENNA__07359__C net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08045_ _02856_ _02879_ vssd1 vssd1 vccd1 vccd1 _02881_ sky130_fd_sc_hd__or2_1
XFILLER_134_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold920 datapath.rf.registers\[2\]\[10\] vssd1 vssd1 vccd1 vccd1 net2268 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1132_A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold931 datapath.rf.registers\[13\]\[3\] vssd1 vssd1 vccd1 vccd1 net2279 sky130_fd_sc_hd__dlygate4sd3_1
Xhold942 datapath.rf.registers\[0\]\[7\] vssd1 vssd1 vccd1 vccd1 net2290 sky130_fd_sc_hd__dlygate4sd3_1
Xhold953 datapath.rf.registers\[6\]\[20\] vssd1 vssd1 vccd1 vccd1 net2301 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10167__A1 _04178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold964 datapath.rf.registers\[16\]\[15\] vssd1 vssd1 vccd1 vccd1 net2312 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold975 datapath.rf.registers\[25\]\[9\] vssd1 vssd1 vccd1 vccd1 net2323 sky130_fd_sc_hd__dlygate4sd3_1
Xhold986 datapath.rf.registers\[31\]\[29\] vssd1 vssd1 vccd1 vccd1 net2334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold997 datapath.rf.registers\[18\]\[31\] vssd1 vssd1 vccd1 vccd1 net2345 sky130_fd_sc_hd__dlygate4sd3_1
X_09996_ _04723_ _04816_ vssd1 vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__or2_1
XFILLER_135_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11609__C net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10513__C _05314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09871__A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08947_ _01981_ _02026_ net444 vssd1 vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout478_X net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout857_A net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_84_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11906__A _02587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12501__S net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08878_ _03710_ _03713_ net343 vssd1 vssd1 vccd1 vccd1 _03714_ sky130_fd_sc_hd__mux2_1
XANTENNA__08487__A _01663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07335__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07829_ datapath.rf.registers\[14\]\[14\] net775 net719 datapath.rf.registers\[20\]\[14\]
+ _02663_ vssd1 vssd1 vccd1 vccd1 _02665_ sky130_fd_sc_hd__a221o_1
XFILLER_84_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11117__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10840_ datapath.PC\[15\] _05583_ datapath.PC\[16\] vssd1 vssd1 vccd1 vccd1 _05594_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_72_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_99_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12092__A1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08296__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10771_ _01441_ net655 _05534_ _05535_ vssd1 vssd1 vccd1 vccd1 _05536_ sky130_fd_sc_hd__o22a_1
XANTENNA__12092__B2 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_145_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_145_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout812_X net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_142_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12510_ datapath.multiplication_module.multiplier_i\[0\] datapath.multiplication_module.multiplicand_i\[0\]
+ datapath.mulitply_result\[0\] vssd1 vssd1 vccd1 vccd1 _06372_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06846__A1 _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13490_ clknet_leaf_33_clk _00300_ net1123 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12441_ _05998_ net156 vssd1 vssd1 vccd1 vccd1 _06368_ sky130_fd_sc_hd__nor2_1
XFILLER_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_22_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12372_ _06332_ datapath.PC\[0\] net190 vssd1 vssd1 vccd1 vccd1 _00811_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07269__C net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14111_ clknet_leaf_110_clk _00877_ net1202 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11323_ net1641 net253 net415 vssd1 vssd1 vccd1 vccd1 _00368_ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_0_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_0_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09765__B _04600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11254_ net256 net2356 net419 vssd1 vssd1 vccd1 vccd1 _00303_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_37_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14042_ clknet_leaf_67_clk _00811_ net1239 vssd1 vssd1 vccd1 vccd1 datapath.PC\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10205_ datapath.PC\[23\] net1260 _05033_ _05040_ vssd1 vssd1 vccd1 vccd1 _05041_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__06901__C net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11185_ net267 datapath.rf.registers\[10\]\[11\] net424 vssd1 vssd1 vccd1 vccd1 _00237_
+ sky130_fd_sc_hd__mux2_1
XFILLER_122_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10136_ net894 _04023_ vssd1 vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__or2_1
X_10067_ _04898_ _04902_ _04893_ vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_50_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07326__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08523__A1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkload1_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11027__S net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13826_ clknet_leaf_113_clk _00635_ net1195 vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__dfrtp_1
XFILLER_62_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08287__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13757_ clknet_leaf_76_clk _00566_ net1248 vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_136_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_136_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10866__S net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12647__A datapath.mulitply_result\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10969_ datapath.mulitply_result\[2\] net598 net621 vssd1 vssd1 vccd1 vccd1 _05705_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_16_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12708_ _06534_ _06535_ vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__and2b_1
XFILLER_149_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13688_ clknet_leaf_7_clk _00498_ net1070 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08563__C _01831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12639_ _06477_ _06478_ _06476_ vssd1 vssd1 vccd1 vccd1 _06480_ sky130_fd_sc_hd__o21ai_1
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12386__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06932__X _01768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire180 _05202_ vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__buf_1
X_14309_ clknet_leaf_121_clk _01014_ net1199 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold205 datapath.multiplication_module.multiplicand_i\[13\] vssd1 vssd1 vccd1 vccd1
+ net1553 sky130_fd_sc_hd__dlygate4sd3_1
Xhold216 datapath.rf.registers\[5\]\[3\] vssd1 vssd1 vccd1 vccd1 net1564 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09539__A0 _03205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold227 datapath.rf.registers\[23\]\[2\] vssd1 vssd1 vccd1 vccd1 net1575 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold238 datapath.rf.registers\[5\]\[21\] vssd1 vssd1 vccd1 vccd1 net1586 sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 datapath.rf.registers\[2\]\[21\] vssd1 vssd1 vccd1 vccd1 net1597 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07476__A _02311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08211__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout707 net709 vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__clkbuf_4
X_09850_ _02545_ _03449_ _03513_ _04085_ vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__a211o_1
Xfanout718 net721 vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__buf_4
XFILLER_59_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout729 _01812_ vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__buf_2
X_08801_ _03636_ vssd1 vssd1 vccd1 vccd1 _03637_ sky130_fd_sc_hd__inv_2
XFILLER_98_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09781_ _04004_ _04616_ _03676_ vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__mux2_1
XFILLER_86_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06993_ net963 _01823_ vssd1 vssd1 vccd1 vccd1 _01829_ sky130_fd_sc_hd__and2_1
XFILLER_100_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Left_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08732_ _03536_ _03537_ _03567_ vssd1 vssd1 vccd1 vccd1 _03568_ sky130_fd_sc_hd__and3_1
X_08663_ _02217_ _02240_ vssd1 vssd1 vccd1 vccd1 _03499_ sky130_fd_sc_hd__or2_2
XANTENNA_fanout173_A _05684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07614_ datapath.rf.registers\[11\]\[18\] net882 net821 datapath.rf.registers\[22\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_68_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10872__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08594_ _03032_ _03429_ _03033_ vssd1 vssd1 vccd1 vccd1 _03430_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_101_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07545_ datapath.rf.registers\[14\]\[20\] net774 net679 datapath.rf.registers\[6\]\[20\]
+ _02371_ vssd1 vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__a221o_1
XFILLER_81_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_138_Right_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_127_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_127_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08817__A2 _03417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13152__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1082_A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_5_0_clk_X clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout438_A net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07476_ _02311_ vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_81_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09215_ _03503_ net627 net624 _03504_ net644 vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__a221oi_1
XANTENNA__12991__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout226_X net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout605_A net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09146_ net365 _03763_ _03630_ vssd1 vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09778__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06842__X _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10388__A1 _01610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08770__A _01859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09077_ _03892_ _03902_ _03912_ _03871_ net605 vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_116_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12292__A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08450__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11400__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08028_ datapath.rf.registers\[22\]\[10\] net736 net696 datapath.rf.registers\[8\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02864_ sky130_fd_sc_hd__a22o_1
Xhold750 datapath.rf.registers\[12\]\[6\] vssd1 vssd1 vccd1 vccd1 net2098 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout974_A net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold761 datapath.rf.registers\[3\]\[28\] vssd1 vssd1 vccd1 vccd1 net2109 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout595_X net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold772 datapath.rf.registers\[11\]\[10\] vssd1 vssd1 vccd1 vccd1 net2120 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_112_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold783 datapath.rf.registers\[17\]\[12\] vssd1 vssd1 vccd1 vccd1 net2131 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold794 datapath.rf.registers\[3\]\[18\] vssd1 vssd1 vccd1 vccd1 net2142 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09979_ datapath.PC\[21\] net596 vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout762_X net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12990_ net178 net2577 net480 vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11941_ net2569 net160 vssd1 vssd1 vccd1 vccd1 _05991_ sky130_fd_sc_hd__nand2_1
XFILLER_44_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08010__A net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07552__C net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14660_ clknet_leaf_22_clk _01365_ net1156 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11872_ screen.register.currentYbus\[5\] net161 vssd1 vssd1 vccd1 vccd1 _05945_ sky130_fd_sc_hd__nand2_1
X_13611_ clknet_leaf_55_clk _00421_ net1179 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10823_ _04272_ _05579_ net900 vssd1 vssd1 vccd1 vccd1 _05580_ sky130_fd_sc_hd__mux2_1
XANTENNA__08269__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_118_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_118_clk
+ sky130_fd_sc_hd__clkbuf_8
X_14591_ clknet_leaf_12_clk _01296_ net1082 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_105_Right_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06736__Y _01575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08664__B net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13062__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13542_ clknet_leaf_28_clk _00352_ net1133 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10754_ net897 _05276_ vssd1 vssd1 vccd1 vccd1 _05521_ sky130_fd_sc_hd__or2_1
XANTENNA__09481__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10685_ keypad.alpha _05459_ _05466_ vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__and3_1
X_13473_ clknet_leaf_25_clk _00283_ net1159 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_12424_ net1389 net130 _06359_ vssd1 vssd1 vccd1 vccd1 _00836_ sky130_fd_sc_hd__a21o_1
XANTENNA__08680__A _02567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08441__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12355_ net893 _03827_ vssd1 vssd1 vccd1 vccd1 _06320_ sky130_fd_sc_hd__or2_1
XANTENNA__06912__B net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11310__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07795__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11306_ _01648_ _03264_ vssd1 vssd1 vccd1 vccd1 _05724_ sky130_fd_sc_hd__or2_1
X_12286_ _06268_ _06270_ datapath.PC\[8\] net308 vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_142_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14025_ clknet_leaf_81_clk _00794_ net1255 vssd1 vssd1 vccd1 vccd1 datapath.PC\[15\]
+ sky130_fd_sc_hd__dfrtp_4
X_11237_ net182 net1843 net527 vssd1 vssd1 vccd1 vccd1 _00287_ sky130_fd_sc_hd__mux2_1
XFILLER_106_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_52_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11168_ net186 net2579 net531 vssd1 vssd1 vccd1 vccd1 _00221_ sky130_fd_sc_hd__mux2_1
X_10119_ datapath.PC\[21\] _03745_ vssd1 vssd1 vccd1 vccd1 _04955_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_147_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11099_ net194 net2014 net535 vssd1 vssd1 vccd1 vccd1 _00156_ sky130_fd_sc_hd__mux2_1
XFILLER_36_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13809_ clknet_leaf_73_clk _00618_ net1250 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[30\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_109_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_109_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09457__C1 _03614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12377__A _04909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08574__B net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07330_ datapath.rf.registers\[26\]\[24\] net837 net795 datapath.rf.registers\[31\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_63_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07261_ datapath.rf.registers\[10\]\[25\] net987 net937 vssd1 vssd1 vccd1 vccd1 _02097_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_14_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09000_ _03834_ _03835_ net367 vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__mux2_1
XFILLER_136_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07192_ datapath.rf.registers\[22\]\[27\] net735 net669 datapath.rf.registers\[21\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02028_ sky130_fd_sc_hd__a22o_1
XFILLER_144_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11220__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07786__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09902_ _01656_ _03670_ net604 vssd1 vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__a21o_1
Xfanout504 net505 vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__buf_2
Xfanout515 _05731_ vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__buf_4
XANTENNA__07538__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout526 _05721_ vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12531__A2 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout537 _05714_ vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__clkbuf_4
X_09833_ _04668_ _03828_ _02094_ _02092_ vssd1 vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__and4b_1
Xfanout548 _03656_ vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__buf_2
Xfanout559 _03320_ vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13147__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout388_A net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06884__A_N _01630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09764_ net630 _04587_ _04598_ _04599_ vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__a2bb2o_2
X_06976_ net965 net908 _01800_ vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__and3_2
XFILLER_132_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08715_ _03549_ _03550_ vssd1 vssd1 vccd1 vccd1 _03551_ sky130_fd_sc_hd__nand2_1
XANTENNA__12986__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09695_ _03538_ _03718_ _04530_ _01622_ vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__o211a_1
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08646_ _01910_ _01911_ vssd1 vssd1 vccd1 vccd1 _03482_ sky130_fd_sc_hd__nand2_1
XFILLER_27_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11903__B screen.counter.ack vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12287__A net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout722_A net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08577_ datapath.rf.registers\[5\]\[0\] net969 _01831_ vssd1 vssd1 vccd1 vccd1 _03413_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12598__A2 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07528_ datapath.rf.registers\[0\]\[20\] net870 _02363_ vssd1 vssd1 vccd1 vccd1 _02364_
+ sky130_fd_sc_hd__o21a_2
XFILLER_22_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07459_ datapath.rf.registers\[11\]\[21\] net882 net836 datapath.rf.registers\[26\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout510_X net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1252_X net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10470_ screen.counter.ct\[9\] _05297_ _05298_ _05299_ vssd1 vssd1 vccd1 vccd1 _05300_
+ sky130_fd_sc_hd__or4_1
XANTENNA__09215__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09129_ _03963_ _03964_ net350 vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__a21o_1
XFILLER_151_702 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11130__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12140_ _05292_ net567 vssd1 vssd1 vccd1 vccd1 _06175_ sky130_fd_sc_hd__nor2_1
XANTENNA__08974__A1 _03320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12071_ _05782_ _06108_ _06110_ vssd1 vssd1 vccd1 vccd1 _06111_ sky130_fd_sc_hd__or3_1
XFILLER_151_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold580 datapath.rf.registers\[23\]\[7\] vssd1 vssd1 vccd1 vccd1 net1928 sky130_fd_sc_hd__dlygate4sd3_1
Xhold591 datapath.rf.registers\[5\]\[30\] vssd1 vssd1 vccd1 vccd1 net1939 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08187__C1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11022_ net219 net1584 net538 vssd1 vssd1 vccd1 vccd1 _00084_ sky130_fd_sc_hd__mux2_1
XFILLER_150_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13057__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08659__B _02190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07563__B net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12896__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12973_ net267 net1983 net480 vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__mux2_1
XANTENNA__12286__B2 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1280 screen.register.currentYbus\[20\] vssd1 vssd1 vccd1 vccd1 net2628 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1291 datapath.rf.registers\[3\]\[25\] vssd1 vssd1 vccd1 vccd1 net2639 sky130_fd_sc_hd__dlygate4sd3_1
X_11924_ _02283_ net656 vssd1 vssd1 vccd1 vccd1 _05980_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_142_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07162__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07701__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14643_ clknet_leaf_36_clk _01348_ net1129 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_72_Left_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11855_ _04909_ _05073_ _05285_ _05932_ net659 vssd1 vssd1 vccd1 vccd1 _05933_ sky130_fd_sc_hd__o41a_2
XANTENNA__11305__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08394__B _03228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06907__B _01720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10806_ datapath.PC\[11\] _05559_ vssd1 vssd1 vccd1 vccd1 _05565_ sky130_fd_sc_hd__and2_1
XFILLER_14_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14574_ clknet_leaf_0_clk _01279_ net1055 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11786_ net616 datapath.ack_mul vssd1 vssd1 vccd1 vccd1 _05898_ sky130_fd_sc_hd__or2_1
XANTENNA__06626__C datapath.ru.latched_instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13525_ clknet_leaf_19_clk _00335_ net1116 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10737_ net1549 net568 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[23\]
+ sky130_fd_sc_hd__and2_1
XFILLER_9_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13456_ clknet_leaf_24_clk _00266_ net1160 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10668_ net1013 _05471_ _05464_ vssd1 vssd1 vccd1 vccd1 _05487_ sky130_fd_sc_hd__o21bai_1
XANTENNA__06923__A net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12407_ _05964_ net157 vssd1 vssd1 vccd1 vccd1 _06351_ sky130_fd_sc_hd__nor2_1
X_10599_ screen.register.currentYbus\[13\] screen.register.currentYbus\[12\] screen.register.currentYbus\[15\]
+ screen.register.currentYbus\[14\] vssd1 vssd1 vccd1 vccd1 _05420_ sky130_fd_sc_hd__or4_1
X_13387_ clknet_leaf_56_clk _00197_ net1161 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11040__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 SEL_O[2] sky130_fd_sc_hd__buf_2
XANTENNA__07768__A2 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08965__A1 _02912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput118 net118 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__buf_2
X_12338_ net894 _03978_ _06306_ _06307_ vssd1 vssd1 vccd1 vccd1 _06308_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_81_Left_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09953__B _03150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12269_ _05002_ net307 _06257_ _06253_ _05526_ vssd1 vssd1 vccd1 vccd1 _06258_ sky130_fd_sc_hd__a32o_1
XFILLER_96_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14008_ clknet_leaf_109_clk net1352 net1220 vssd1 vssd1 vccd1 vccd1 screen.screenEdge.enable2
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07754__A net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09390__A1 _02418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06830_ _01505_ net1004 net1020 net1028 datapath.ru.latched_instruction\[21\] vssd1
+ vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__a32o_4
X_06761_ datapath.ru.latched_instruction\[27\] net1030 net994 _01597_ vssd1 vssd1
+ vccd1 vccd1 _01598_ sky130_fd_sc_hd__a22oi_4
XFILLER_49_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09142__A1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08500_ datapath.rf.registers\[10\]\[1\] net709 _03333_ _03334_ _03335_ vssd1 vssd1
+ vccd1 vccd1 _03336_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09142__B2 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06692_ datapath.ru.latched_instruction\[6\] _01485_ _01528_ _01529_ _01530_ vssd1
+ vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__a2111o_1
X_09480_ net370 _04290_ _04288_ net327 vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_19_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_90_Left_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07153__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08431_ datapath.rf.registers\[31\]\[2\] net966 _01825_ vssd1 vssd1 vccd1 vccd1 _03267_
+ sky130_fd_sc_hd__and3_1
XANTENNA__06900__B1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11215__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08362_ datapath.rf.registers\[28\]\[3\] net806 _03178_ _03181_ _03190_ vssd1 vssd1
+ vccd1 vccd1 _03198_ sky130_fd_sc_hd__a2111o_1
X_07313_ datapath.rf.registers\[21\]\[24\] net946 net923 vssd1 vssd1 vccd1 vccd1 _02149_
+ sky130_fd_sc_hd__and3_1
XFILLER_149_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08293_ datapath.rf.registers\[22\]\[4\] net821 net817 datapath.rf.registers\[7\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__a22o_1
XFILLER_20_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout136_A _05934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07244_ datapath.rf.registers\[26\]\[26\] net778 net758 datapath.rf.registers\[30\]\[26\]
+ _02071_ vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__a221o_1
XFILLER_137_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07175_ datapath.rf.registers\[9\]\[27\] net886 net808 datapath.rf.registers\[27\]\[27\]
+ _02010_ vssd1 vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__a221o_1
XFILLER_117_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07759__A2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10763__A1 _01450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_93_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1212_A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout301 _05529_ vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout312 _03620_ vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout323 _03674_ vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__clkbuf_2
Xfanout334 _05904_ vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout672_A net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout345 net348 vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__buf_2
Xfanout356 net357 vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08184__A2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout367 net369 vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__clkbuf_4
X_09816_ net312 _04650_ _04651_ _03641_ vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__o22a_1
Xfanout378 _03621_ vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout389 _06560_ vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__buf_4
XANTENNA__07392__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07931__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09747_ _04239_ _04272_ _04582_ vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_129_Left_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06959_ _01636_ net990 vssd1 vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__nor2_2
XANTENNA_fanout558_X net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout937_A _01720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10279__B1 net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09133__A1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09678_ _03430_ _03565_ vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__xnor2_1
XFILLER_15_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08629_ _02147_ _03464_ vssd1 vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_124_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout725_X net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11125__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11640_ _05788_ _05863_ vssd1 vssd1 vccd1 vccd1 _05864_ sky130_fd_sc_hd__and2b_1
XFILLER_52_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11571_ net1008 _05765_ vssd1 vssd1 vccd1 vccd1 _05795_ sky130_fd_sc_hd__or2_2
XANTENNA__10964__S net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10817__X _05575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13310_ clknet_leaf_150_clk _00120_ net1059 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11794__A3 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10522_ _01423_ net1273 screen.counter.ct\[18\] screen.counter.ct\[21\] vssd1 vssd1
+ vccd1 vccd1 _05352_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_138_Left_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14290_ clknet_leaf_91_clk _00995_ net1232 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_109_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13241_ clknet_leaf_31_clk _00051_ net1122 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10453_ _04909_ _05073_ _05204_ _05282_ vssd1 vssd1 vccd1 vccd1 _05288_ sky130_fd_sc_hd__or4_4
XANTENNA__07558__B net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10384_ net369 _04375_ _05219_ net372 vssd1 vssd1 vccd1 vccd1 _05220_ sky130_fd_sc_hd__o211a_1
X_13172_ net2527 vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12123_ net1277 _05907_ _06154_ vssd1 vssd1 vccd1 vccd1 _06160_ sky130_fd_sc_hd__nand3_1
XFILLER_123_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12054_ screen.register.currentYbus\[28\] _05786_ net995 screen.register.currentXbus\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06095_ sky130_fd_sc_hd__a22o_1
XANTENNA__07574__A net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08175__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11005_ net258 net1563 net541 vssd1 vssd1 vccd1 vccd1 _00067_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_144_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07383__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout890 net896 vssd1 vssd1 vccd1 vccd1 net890 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07922__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_13_0_clk_X clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12956_ net187 net1841 net395 vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__mux2_1
XFILLER_34_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07135__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11907_ net136 _05968_ _05967_ vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07686__A1 datapath.rf.registers\[0\]\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12887_ net201 net2263 net399 vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__mux2_1
XANTENNA__11035__S net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14626_ clknet_leaf_152_clk _01331_ net1054 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11838_ screen.counter.ct\[17\] _01425_ _05806_ _05916_ vssd1 vssd1 vccd1 vccd1 _05917_
+ sky130_fd_sc_hd__or4_1
XFILLER_61_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14557_ clknet_leaf_146_clk _01262_ net1091 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10874__S net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11769_ net1499 net143 net138 _01954_ vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_60_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_40_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_clk sky130_fd_sc_hd__clkbuf_8
X_13508_ clknet_leaf_22_clk _00318_ net1156 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07989__A2 _02824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14488_ clknet_leaf_7_clk _01193_ net1068 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_155_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13439_ clknet_leaf_11_clk _00249_ net1082 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08980_ net344 _03811_ _03812_ _03815_ vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_58_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07931_ datapath.rf.registers\[10\]\[12\] net707 net661 datapath.rf.registers\[5\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02767_ sky130_fd_sc_hd__a22o_1
XANTENNA__08166__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07862_ datapath.rf.registers\[11\]\[13\] net882 net854 datapath.rf.registers\[19\]\[13\]
+ _02684_ vssd1 vssd1 vccd1 vccd1 _02698_ sky130_fd_sc_hd__a221o_1
XFILLER_96_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09601_ net325 _04043_ _04435_ _04436_ vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__o22ai_4
XFILLER_96_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06813_ _01490_ _01568_ net1029 datapath.ru.latched_instruction\[10\] vssd1 vssd1
+ vccd1 vccd1 _01649_ sky130_fd_sc_hd__a2bb2o_1
X_07793_ datapath.rf.registers\[9\]\[15\] net703 _02626_ _02628_ net787 vssd1 vssd1
+ vccd1 vccd1 _02629_ sky130_fd_sc_hd__a2111oi_1
X_09532_ net906 _03550_ net626 _03545_ _04367_ vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__a221o_1
X_06744_ _01502_ net1005 net1021 net1031 datapath.ru.latched_instruction\[1\] vssd1
+ vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__a32o_1
XFILLER_37_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07126__B1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06828__A _01663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06675_ datapath.ru.latched_instruction\[14\] _01513_ vssd1 vssd1 vccd1 vccd1 _01514_
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_35_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09463_ _03604_ _04276_ _04297_ _04298_ vssd1 vssd1 vccd1 vccd1 _04299_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout253_A _05588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08414_ datapath.rf.registers\[16\]\[2\] net863 _03242_ _03246_ _03247_ vssd1 vssd1
+ vccd1 vccd1 _03250_ sky130_fd_sc_hd__a2111o_1
X_09394_ _04227_ _04229_ _03625_ vssd1 vssd1 vccd1 vccd1 _04230_ sky130_fd_sc_hd__mux2_1
XANTENNA__10069__B net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08087__D1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08345_ datapath.rf.registers\[27\]\[3\] net979 net938 vssd1 vssd1 vccd1 vccd1 _03181_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout420_A _05722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_31_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1162_A net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout518_A net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13160__S net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10433__B1 net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08276_ datapath.rf.registers\[3\]\[5\] net771 net763 datapath.rf.registers\[1\]\[5\]
+ _03111_ vssd1 vssd1 vccd1 vccd1 _03112_ sky130_fd_sc_hd__a221o_1
XFILLER_137_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07227_ datapath.rf.registers\[5\]\[26\] net819 _02061_ _02062_ net872 vssd1 vssd1
+ vccd1 vccd1 _02063_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_95_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout306_X net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08929__A1 _01980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07158_ datapath.rf.registers\[25\]\[28\] net729 _01993_ net789 vssd1 vssd1 vccd1
+ vccd1 _01994_ sky130_fd_sc_hd__a211o_1
XFILLER_133_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout887_A net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11909__A _02542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07062__C1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07089_ datapath.rf.registers\[12\]\[29\] net827 net813 datapath.rf.registers\[23\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__a22o_1
XANTENNA__12504__S net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1107 net1110 vssd1 vssd1 vccd1 vccd1 net1107 sky130_fd_sc_hd__clkbuf_2
Xfanout1118 net1119 vssd1 vssd1 vccd1 vccd1 net1118 sky130_fd_sc_hd__clkbuf_2
Xfanout131 net132 vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__buf_2
XANTENNA_fanout675_X net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_98_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_98_clk sky130_fd_sc_hd__clkbuf_8
Xfanout1129 net1130 vssd1 vssd1 vccd1 vccd1 net1129 sky130_fd_sc_hd__clkbuf_4
Xfanout142 _05891_ vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08157__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout153 net155 vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__buf_1
XFILLER_75_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout164 net165 vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08777__X _03613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout175 _05684_ vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__buf_1
XANTENNA__08002__B net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout186 net187 vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_126_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout197 net198 vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__clkbuf_2
XFILLER_74_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout842_X net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12810_ net1587 net256 net491 vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__mux2_1
X_13790_ clknet_leaf_74_clk _00599_ net1242 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09114__A _03947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08865__A0 _02613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12741_ net2353 net272 net404 vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__mux2_1
XANTENNA__07560__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12672_ _06502_ _06506_ vssd1 vssd1 vccd1 vccd1 _06507_ sky130_fd_sc_hd__and2_1
XFILLER_31_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14411_ clknet_leaf_55_clk _01116_ net1173 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_146_Left_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11623_ _05846_ vssd1 vssd1 vccd1 vccd1 _05847_ sky130_fd_sc_hd__inv_2
XANTENNA__09768__B _04057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_22_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__13070__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14342_ clknet_leaf_29_clk _01047_ net1131 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11554_ net1006 _05777_ vssd1 vssd1 vccd1 vccd1 _05778_ sky130_fd_sc_hd__nor2_4
XFILLER_144_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10505_ _05315_ _05326_ _05334_ vssd1 vssd1 vccd1 vccd1 _05335_ sky130_fd_sc_hd__nor3_4
XTAP_TAPCELL_ROW_137_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14273_ clknet_leaf_45_clk _00978_ net1172 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_21_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11485_ net284 net2333 net512 vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__mux2_1
XFILLER_137_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire587 net588 vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__clkbuf_1
XFILLER_12_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13224_ clknet_leaf_60_clk _00034_ net1169 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10436_ _04338_ _04395_ vssd1 vssd1 vccd1 vccd1 _05272_ sky130_fd_sc_hd__or2_1
XFILLER_136_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10727__A1 _02704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13155_ net2281 net185 net382 vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__mux2_1
XFILLER_98_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10367_ _05126_ _05136_ _05157_ vssd1 vssd1 vccd1 vccd1 _05203_ sky130_fd_sc_hd__nor3_1
XANTENNA__06920__B net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12106_ _06089_ _06140_ _06143_ vssd1 vssd1 vccd1 vccd1 _06144_ sky130_fd_sc_hd__o21ai_1
XFILLER_124_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_155_Left_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13086_ net1747 net199 net386 vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__mux2_1
X_10298_ _04843_ _05133_ vssd1 vssd1 vccd1 vccd1 _05134_ sky130_fd_sc_hd__nand2_1
X_12037_ screen.register.currentXbus\[3\] net1000 _05837_ screen.register.currentYbus\[19\]
+ vssd1 vssd1 vccd1 vccd1 _06079_ sky130_fd_sc_hd__a22o_1
XFILLER_77_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07356__B1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07108__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13988_ clknet_leaf_108_clk _00765_ net1219 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12101__B1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08566__C _01797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12939_ net272 net1697 net396 vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__mux2_1
X_14609_ clknet_leaf_41_clk _01314_ net1143 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_13_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_8
X_08130_ datapath.rf.registers\[16\]\[8\] net740 net720 datapath.rf.registers\[20\]\[8\]
+ _02965_ vssd1 vssd1 vccd1 vccd1 _02966_ sky130_fd_sc_hd__a221o_1
XANTENNA_wire590_A _02428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10966__A1 _01502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08061_ datapath.rf.registers\[9\]\[9\] net986 net944 vssd1 vssd1 vccd1 vccd1 _02897_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10109__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07012_ datapath.rf.registers\[3\]\[31\] net770 net714 datapath.rf.registers\[4\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01848_ sky130_fd_sc_hd__a22o_1
XANTENNA__10179__C1 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10718__A1 _03104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08387__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07595__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08963_ net338 _03798_ _03788_ _03673_ vssd1 vssd1 vccd1 vccd1 _03799_ sky130_fd_sc_hd__o211ai_1
XANTENNA__08139__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07914_ _02741_ net586 datapath.rf.registers\[0\]\[12\] net870 vssd1 vssd1 vccd1
+ vccd1 _02750_ sky130_fd_sc_hd__o2bb2a_2
X_08894_ datapath.i_ack datapath.pc_module.i_ack2 vssd1 vssd1 vccd1 vccd1 _03730_
+ sky130_fd_sc_hd__nand2b_1
XANTENNA__07347__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07845_ net612 _02680_ net564 vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__a21o_1
XANTENNA__11694__A2 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout468_A net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13155__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07776_ datapath.rf.registers\[0\]\[15\] net871 _02599_ _02611_ vssd1 vssd1 vccd1
+ vccd1 _02612_ sky130_fd_sc_hd__o22a_4
XFILLER_140_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09515_ _04349_ _04350_ vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_88_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06727_ _01407_ datapath.pc_module.i_ack2 datapath.ru.n_memwrite2 net1031 datapath.ru.zero_multi1
+ vssd1 vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__a311oi_2
XANTENNA__08847__A0 _03228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout635_A net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08311__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06708__D datapath.ru.latched_instruction\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09446_ net455 _04247_ _04281_ vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__a21o_1
X_06658_ mmio.memload_or_instruction\[29\] net1050 vssd1 vssd1 vccd1 vccd1 _01497_
+ sky130_fd_sc_hd__and2_2
XANTENNA__08773__A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout423_X net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09377_ _04069_ _04158_ net461 vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout802_A _01769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06589_ keypad.alpha vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__inv_2
XANTENNA__11403__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08328_ datapath.rf.registers\[19\]\[4\] net730 _03162_ _03163_ net787 vssd1 vssd1
+ vccd1 vccd1 _03164_ sky130_fd_sc_hd__a2111o_1
XFILLER_149_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14283__Q datapath.rf.registers\[0\]\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08259_ datapath.rf.registers\[5\]\[5\] net819 net811 datapath.rf.registers\[13\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03095_ sky130_fd_sc_hd__a22o_1
XFILLER_137_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11270_ net184 net2332 net419 vssd1 vssd1 vccd1 vccd1 _00319_ sky130_fd_sc_hd__mux2_1
Xteam_04_1340 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] team_04_1340/LO sky130_fd_sc_hd__conb_1
XANTENNA__09024__B1 _03721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10709__A1 _02680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout792_X net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08378__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10221_ net1044 _05056_ _05054_ net898 vssd1 vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__o211a_1
XANTENNA__07586__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09891__X _04727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10152_ datapath.PC\[20\] _04084_ net469 vssd1 vssd1 vccd1 vccd1 _04988_ sky130_fd_sc_hd__mux2_1
XFILLER_0_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07555__C net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10262__B _04272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10830__X _05586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10083_ _04916_ _04918_ datapath.PC\[30\] net1258 vssd1 vssd1 vccd1 vccd1 _04919_
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__07338__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold9 keypad.debounce.debounce\[8\] vssd1 vssd1 vccd1 vccd1 net1357 sky130_fd_sc_hd__dlygate4sd3_1
X_13911_ clknet_leaf_43_clk net1366 net1149 vssd1 vssd1 vccd1 vccd1 keypad.debounce.debounce\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input29_A DAT_I[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13065__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10893__B1 _05635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13842_ clknet_leaf_115_clk _00651_ net1195 vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__dfrtp_1
X_13773_ clknet_leaf_81_clk _00582_ net1255 vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__dfrtp_1
XFILLER_15_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10985_ net1618 net243 net435 vssd1 vssd1 vccd1 vccd1 _00050_ sky130_fd_sc_hd__mux2_1
XANTENNA__08302__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12724_ _05893_ _06544_ _06545_ _06530_ vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_26_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08683__A _02612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_139_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12655_ _06491_ _06492_ vssd1 vssd1 vccd1 vccd1 _06493_ sky130_fd_sc_hd__nand2_1
XANTENNA__11313__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11606_ _05829_ vssd1 vssd1 vccd1 vccd1 _05830_ sky130_fd_sc_hd__inv_2
XFILLER_11_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12586_ _06431_ _06433_ _06430_ vssd1 vssd1 vccd1 vccd1 _06435_ sky130_fd_sc_hd__a21boi_2
X_14325_ clknet_leaf_130_clk _01030_ net1111 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11537_ screen.counter.ct\[1\] screen.counter.ct\[0\] screen.counter.ct\[2\] vssd1
+ vssd1 vccd1 vccd1 _05761_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_152_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold409 datapath.rf.registers\[11\]\[7\] vssd1 vssd1 vccd1 vccd1 net1757 sky130_fd_sc_hd__dlygate4sd3_1
X_14256_ clknet_leaf_24_clk _00961_ net1160 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11468_ net1691 net201 net407 vssd1 vssd1 vccd1 vccd1 _00506_ sky130_fd_sc_hd__mux2_1
XFILLER_143_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13207_ clknet_leaf_131_clk _00017_ net1114 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09566__A1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10419_ net358 _04521_ _05254_ net345 vssd1 vssd1 vccd1 vccd1 _05255_ sky130_fd_sc_hd__a211o_1
X_14187_ clknet_leaf_75_clk net1385 net1246 vssd1 vssd1 vccd1 vccd1 datapath.pc_module.i_ack1
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10453__A _04909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11399_ net1760 net211 net410 vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__mux2_1
XFILLER_98_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07041__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13138_ net1737 net270 net384 vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__mux2_1
XANTENNA__09318__A1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13069_ net1659 net285 net388 vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__mux2_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1109 datapath.rf.registers\[3\]\[22\] vssd1 vssd1 vccd1 vccd1 net2457 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_39_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_119_Right_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08577__B net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10884__A0 _04023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07630_ _02458_ _02465_ datapath.rf.registers\[0\]\[18\] net867 vssd1 vssd1 vccd1
+ vccd1 _02466_ sky130_fd_sc_hd__o2bb2a_4
X_07561_ datapath.rf.registers\[9\]\[19\] net886 net791 datapath.rf.registers\[18\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__a22o_1
XFILLER_80_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09300_ _03642_ net347 _04135_ net649 vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__o31a_1
X_07492_ datapath.rf.registers\[1\]\[21\] net762 net671 datapath.rf.registers\[7\]\[21\]
+ _02322_ vssd1 vssd1 vccd1 vccd1 _02328_ sky130_fd_sc_hd__a221o_1
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09231_ net372 _04064_ _04065_ net329 vssd1 vssd1 vccd1 vccd1 _04067_ sky130_fd_sc_hd__a211o_1
XANTENNA__11223__S net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09162_ net461 _03929_ _03997_ net354 vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__o211a_1
X_08113_ _02939_ _02946_ _02947_ _02948_ vssd1 vssd1 vccd1 vccd1 _02949_ sky130_fd_sc_hd__or4_1
XFILLER_108_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10915__X _05659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09093_ _02126_ _02170_ net453 vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__mux2_1
XANTENNA__07937__A _02750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08044_ _02856_ _02879_ vssd1 vssd1 vccd1 vccd1 _02880_ sky130_fd_sc_hd__and2_1
XANTENNA__07280__A2 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold910 datapath.rf.registers\[14\]\[19\] vssd1 vssd1 vccd1 vccd1 net2258 sky130_fd_sc_hd__dlygate4sd3_1
Xhold921 datapath.rf.registers\[30\]\[18\] vssd1 vssd1 vccd1 vccd1 net2269 sky130_fd_sc_hd__dlygate4sd3_1
Xhold932 datapath.rf.registers\[28\]\[15\] vssd1 vssd1 vccd1 vccd1 net2280 sky130_fd_sc_hd__dlygate4sd3_1
Xhold943 datapath.rf.registers\[19\]\[8\] vssd1 vssd1 vccd1 vccd1 net2291 sky130_fd_sc_hd__dlygate4sd3_1
Xhold954 datapath.rf.registers\[18\]\[30\] vssd1 vssd1 vccd1 vccd1 net2302 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07656__B net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold965 datapath.rf.registers\[22\]\[19\] vssd1 vssd1 vccd1 vccd1 net2313 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold976 datapath.rf.registers\[16\]\[31\] vssd1 vssd1 vccd1 vccd1 net2324 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12561__B1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold987 screen.counter.currentCt\[3\] vssd1 vssd1 vccd1 vccd1 net2335 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_1_0_clk_X clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold998 datapath.rf.registers\[23\]\[28\] vssd1 vssd1 vccd1 vccd1 net2346 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07032__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09995_ _04821_ _04830_ vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__nor2_1
XANTENNA__12989__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09309__A1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08946_ _03780_ _03781_ net450 vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11906__B net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08877_ _03711_ _03712_ net448 vssd1 vssd1 vccd1 vccd1 _03713_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout752_A _01804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08532__A2 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07828_ datapath.rf.registers\[8\]\[14\] net695 net665 datapath.rf.registers\[15\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__a22o_1
XFILLER_151_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07740__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07759_ datapath.rf.registers\[25\]\[15\] net841 _01772_ datapath.rf.registers\[15\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout540_X net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10770_ datapath.mulitply_result\[5\] net598 net620 vssd1 vssd1 vccd1 vccd1 _05535_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_23_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09429_ net904 _04240_ vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__nor2_1
XFILLER_52_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14027__RESET_B net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout805_X net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11133__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12440_ net1387 net130 _06367_ vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__a21o_1
XFILLER_21_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10972__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12371_ net891 net222 _04781_ _05239_ _06331_ vssd1 vssd1 vccd1 vccd1 _06332_ sky130_fd_sc_hd__a41o_1
XANTENNA__10825__X _05582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14110_ clknet_leaf_111_clk _00876_ net1202 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11322_ net1892 net255 net415 vssd1 vssd1 vccd1 vccd1 _00367_ sky130_fd_sc_hd__mux2_1
XANTENNA__07847__A _02661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14041_ clknet_leaf_88_clk _00810_ net1253 vssd1 vssd1 vccd1 vccd1 datapath.PC\[31\]
+ sky130_fd_sc_hd__dfrtp_4
X_11253_ net265 net2554 net421 vssd1 vssd1 vccd1 vccd1 _00302_ sky130_fd_sc_hd__mux2_1
XANTENNA__07566__B net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10204_ net230 _05037_ _05039_ net1295 vssd1 vssd1 vccd1 vccd1 _05040_ sky130_fd_sc_hd__a31o_1
X_11184_ net272 net2386 net424 vssd1 vssd1 vccd1 vccd1 _00236_ sky130_fd_sc_hd__mux2_1
XANTENNA__12899__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10135_ net894 _04023_ vssd1 vssd1 vccd1 vccd1 _04971_ sky130_fd_sc_hd__nor2_1
XFILLER_79_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08678__A _02523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10066_ _04900_ _04901_ vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__xor2_2
XFILLER_94_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08397__B net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08523__A2 _03357_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09720__B2 _03673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13825_ clknet_leaf_113_clk _00634_ net1195 vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__dfrtp_1
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13756_ clknet_leaf_76_clk _00565_ net1248 vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__dfrtp_1
X_10968_ net1269 _04395_ net897 vssd1 vssd1 vccd1 vccd1 _05704_ sky130_fd_sc_hd__mux2_1
XFILLER_71_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12707_ columns.count\[1\] columns.count\[0\] _06531_ columns.count\[2\] vssd1 vssd1
+ vccd1 vccd1 _06535_ sky130_fd_sc_hd__a31o_1
X_13687_ clknet_leaf_124_clk _00497_ net1208 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10899_ datapath.mulitply_result\[24\] net615 net652 vssd1 vssd1 vccd1 vccd1 _05645_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__11043__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12638_ _06476_ _06477_ _06478_ vssd1 vssd1 vccd1 vccd1 _06479_ sky130_fd_sc_hd__or3_1
XANTENNA__11043__A0 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09787__A1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12569_ datapath.mulitply_result\[10\] datapath.multiplication_module.multiplicand_i\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06421_ sky130_fd_sc_hd__or2_1
XFILLER_156_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14308_ clknet_leaf_20_clk _01013_ net1163 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold206 mmio.memload_or_instruction\[16\] vssd1 vssd1 vccd1 vccd1 net1554 sky130_fd_sc_hd__dlygate4sd3_1
Xhold217 datapath.rf.registers\[31\]\[0\] vssd1 vssd1 vccd1 vccd1 net1565 sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 datapath.rf.registers\[10\]\[5\] vssd1 vssd1 vccd1 vccd1 net1576 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09539__A1 _03263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14239_ clknet_leaf_124_clk datapath.multiplication_module.multiplier_i_n\[7\] net1214
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i\[7\] sky130_fd_sc_hd__dfrtp_1
Xhold239 datapath.rf.registers\[1\]\[13\] vssd1 vssd1 vccd1 vccd1 net1587 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12543__B1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07014__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout708 net709 vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__clkbuf_8
Xfanout719 net721 vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__buf_4
X_08800_ _01574_ _01607_ vssd1 vssd1 vccd1 vccd1 _03636_ sky130_fd_sc_hd__or2_2
X_09780_ _03785_ _03780_ net450 vssd1 vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06992_ net968 net910 _01809_ vssd1 vssd1 vccd1 vccd1 _01828_ sky130_fd_sc_hd__and3_2
XANTENNA__06773__B2 _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07970__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08731_ _02912_ _02936_ _03564_ _03565_ _03539_ vssd1 vssd1 vccd1 vccd1 _03567_ sky130_fd_sc_hd__a221o_1
XANTENNA__10306__C1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11218__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1290 mmio.key_en3 vssd1 vssd1 vccd1 vccd1 net1290 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10857__B1 _05608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10122__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08662_ _02217_ _02240_ vssd1 vssd1 vccd1 vccd1 _03498_ sky130_fd_sc_hd__and2_1
XANTENNA__07722__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10321__A2 net1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07613_ datapath.rf.registers\[30\]\[18\] net832 net818 datapath.rf.registers\[7\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__a22o_1
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_max_cap972_X net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08593_ _03081_ _03128_ _03426_ _03427_ _03080_ vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__a41o_1
XFILLER_81_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout166_A _05288_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07544_ datapath.rf.registers\[1\]\[20\] net762 net664 datapath.rf.registers\[15\]\[20\]
+ _02379_ vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__a221o_1
XFILLER_22_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14191__RESET_B net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07475_ _02300_ _02310_ datapath.rf.registers\[0\]\[21\] net866 vssd1 vssd1 vccd1
+ vccd1 _02311_ sky130_fd_sc_hd__o2bb2a_4
XFILLER_14_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1075_A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09214_ net337 _04047_ _04049_ net322 vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__a211o_1
XANTENNA__09227__A0 _02312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09778__A1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09145_ _03586_ _03980_ net578 vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_101_Left_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout500_A net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1242_A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09076_ net904 _03866_ _03909_ net318 _03911_ vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__o221a_1
X_08027_ datapath.rf.registers\[4\]\[10\] net716 net670 datapath.rf.registers\[21\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__a22o_1
XANTENNA__10093__A net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold740 datapath.rf.registers\[21\]\[30\] vssd1 vssd1 vccd1 vccd1 net2088 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold751 datapath.rf.registers\[16\]\[19\] vssd1 vssd1 vccd1 vccd1 net2099 sky130_fd_sc_hd__dlygate4sd3_1
Xhold762 datapath.rf.registers\[17\]\[19\] vssd1 vssd1 vccd1 vccd1 net2110 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07005__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold773 datapath.rf.registers\[2\]\[12\] vssd1 vssd1 vccd1 vccd1 net2121 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout490_X net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold784 datapath.rf.registers\[31\]\[25\] vssd1 vssd1 vccd1 vccd1 net2132 sky130_fd_sc_hd__dlygate4sd3_1
Xhold795 datapath.rf.registers\[29\]\[5\] vssd1 vssd1 vccd1 vccd1 net2143 sky130_fd_sc_hd__dlygate4sd3_1
X_09978_ _04729_ _04812_ _04730_ _04726_ vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__o211a_1
XANTENNA__07961__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08929_ _01934_ _01980_ net443 vssd1 vssd1 vccd1 vccd1 _03765_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_110_Left_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout755_X net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10540__B net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11128__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11940_ net136 _05990_ _05989_ vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_28_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11871_ net135 _05944_ _05943_ vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__o21ai_1
XFILLER_44_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10967__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11652__A _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13610_ clknet_leaf_59_clk _00420_ net1169 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[13\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10822_ _05578_ vssd1 vssd1 vccd1 vccd1 _05579_ sky130_fd_sc_hd__inv_2
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14590_ clknet_leaf_1_clk _01295_ net1062 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12255__A1_N datapath.multiplication_module.zero_multi vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10539__Y _05367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13541_ clknet_leaf_118_clk _00351_ net1192 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10753_ net897 _04338_ vssd1 vssd1 vccd1 vccd1 _05520_ sky130_fd_sc_hd__nand2_1
XANTENNA__11812__A2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13472_ clknet_leaf_135_clk _00282_ net1098 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_41_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10684_ keypad.alpha _05444_ vssd1 vssd1 vccd1 vccd1 _05501_ sky130_fd_sc_hd__nor2_1
XANTENNA__07492__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12423_ _05980_ net156 vssd1 vssd1 vccd1 vccd1 _06359_ sky130_fd_sc_hd__nor2_1
XFILLER_138_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12354_ datapath.PC\[27\] net309 _06319_ vssd1 vssd1 vccd1 vccd1 _00806_ sky130_fd_sc_hd__a21o_1
XANTENNA__07244__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10715__B net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11305_ net168 net2515 net523 vssd1 vssd1 vccd1 vccd1 _00353_ sky130_fd_sc_hd__mux2_1
XFILLER_4_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12285_ _05550_ _06254_ _06269_ net190 vssd1 vssd1 vccd1 vccd1 _06270_ sky130_fd_sc_hd__o22a_1
XFILLER_107_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12525__B1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14024_ clknet_leaf_77_clk _00793_ net1255 vssd1 vssd1 vccd1 vccd1 datapath.PC\[14\]
+ sky130_fd_sc_hd__dfrtp_4
X_11236_ net178 net1824 net528 vssd1 vssd1 vccd1 vccd1 _00286_ sky130_fd_sc_hd__mux2_1
XANTENNA__07583__Y _02419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11167_ net195 net2223 net530 vssd1 vssd1 vccd1 vccd1 _00220_ sky130_fd_sc_hd__mux2_1
X_10118_ datapath.PC\[19\] net1256 _04950_ _04953_ vssd1 vssd1 vccd1 vccd1 _04954_
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_147_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11098_ net198 net2506 net536 vssd1 vssd1 vccd1 vccd1 _00155_ sky130_fd_sc_hd__mux2_1
XANTENNA__11038__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10049_ _04882_ _04884_ vssd1 vssd1 vccd1 vccd1 _04885_ sky130_fd_sc_hd__nand2_1
XFILLER_91_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13808_ clknet_leaf_73_clk _00617_ net1243 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12056__A2 _05773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12377__B _05073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09032__A net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13739_ clknet_leaf_50_clk _00549_ net1176 vssd1 vssd1 vccd1 vccd1 mmio.key_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_91_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09209__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07260_ datapath.rf.registers\[19\]\[25\] net978 net928 vssd1 vssd1 vccd1 vccd1 _02096_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07483__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07191_ datapath.rf.registers\[17\]\[27\] net747 net723 datapath.rf.registers\[18\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__a22o_1
XFILLER_118_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_83_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11501__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07235__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13513__RESET_B net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09901_ _04727_ _04734_ datapath.PC\[17\] vssd1 vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_98_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout505 _06374_ vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__buf_2
XFILLER_113_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout516 _05731_ vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__clkbuf_8
Xfanout527 _05721_ vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__clkbuf_4
XFILLER_99_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09832_ _03487_ _04628_ vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__or2_1
XANTENNA__12332__S net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout538 net541 vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__clkbuf_8
XFILLER_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_141_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout549 _03655_ vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09763_ net609 _04587_ _04588_ net578 net605 vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__a221oi_1
XFILLER_101_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06975_ _01797_ net907 vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__and2_2
XANTENNA_clkbuf_leaf_21_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08714_ _03263_ _03295_ vssd1 vssd1 vccd1 vccd1 _03550_ sky130_fd_sc_hd__xnor2_2
XFILLER_55_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09694_ _03537_ net625 _04518_ net906 vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__a22oi_1
XFILLER_26_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08645_ _01888_ _01909_ vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__and2_1
XFILLER_27_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08765__B _01603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08576_ datapath.rf.registers\[23\]\[0\] net966 _01820_ vssd1 vssd1 vccd1 vccd1 _03412_
+ sky130_fd_sc_hd__and3_1
XFILLER_42_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_36_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07527_ _02353_ _02358_ _02362_ vssd1 vssd1 vccd1 vccd1 _02363_ sky130_fd_sc_hd__or3_4
XFILLER_23_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout715_A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07458_ datapath.rf.registers\[14\]\[21\] net981 net919 vssd1 vssd1 vccd1 vccd1 _02294_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_33_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08781__A net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10375__X _05211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12507__S net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07389_ datapath.rf.registers\[2\]\[23\] net742 net738 datapath.rf.registers\[16\]\[23\]
+ _02224_ vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__a221o_1
XANTENNA__11411__S net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09128_ _03884_ _03885_ net462 vssd1 vssd1 vccd1 vccd1 _03964_ sky130_fd_sc_hd__a21o_1
XANTENNA__07226__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09059_ _03691_ _03701_ net449 vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__mux2_1
XANTENNA__08005__B net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12070_ screen.register.currentYbus\[21\] _05773_ net997 screen.register.currentXbus\[21\]
+ _06109_ vssd1 vssd1 vccd1 vccd1 _06110_ sky130_fd_sc_hd__a221o_1
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout872_X net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold570 datapath.rf.registers\[27\]\[13\] vssd1 vssd1 vccd1 vccd1 net1918 sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 datapath.rf.registers\[19\]\[26\] vssd1 vssd1 vccd1 vccd1 net1929 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold592 datapath.rf.registers\[27\]\[23\] vssd1 vssd1 vccd1 vccd1 net1940 sky130_fd_sc_hd__dlygate4sd3_1
X_11021_ net241 net1619 net540 vssd1 vssd1 vccd1 vccd1 _00083_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_109_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07563__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_129_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12972_ net271 net2238 net480 vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__mux2_1
Xhold1270 datapath.rf.registers\[3\]\[11\] vssd1 vssd1 vccd1 vccd1 net2618 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input11_A DAT_I[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11923_ net2596 net160 vssd1 vssd1 vccd1 vccd1 _05979_ sky130_fd_sc_hd__nand2_1
Xhold1281 datapath.rf.registers\[9\]\[19\] vssd1 vssd1 vccd1 vccd1 net2629 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1292 datapath.rf.registers\[20\]\[3\] vssd1 vssd1 vccd1 vccd1 net2640 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06747__Y _01586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13073__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14642_ clknet_leaf_32_clk _01347_ net1123 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11854_ _05281_ _05283_ _05282_ vssd1 vssd1 vccd1 vccd1 _05932_ sky130_fd_sc_hd__o21ai_1
X_10805_ net272 net2091 net543 vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__mux2_1
X_14573_ clknet_leaf_126_clk _01278_ net1205 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11785_ keypad.apps.app_c\[0\] net2432 _05896_ vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__mux2_1
XFILLER_25_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08111__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13524_ clknet_leaf_20_clk _00334_ net1118 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10736_ net1612 net568 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[22\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_45_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07465__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08691__A _02751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13455_ clknet_leaf_26_clk _00265_ net1137 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10667_ _05443_ _05468_ _05444_ vssd1 vssd1 vccd1 vccd1 _05486_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06923__B net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11321__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12406_ net1401 net130 _06350_ vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__a21o_1
XANTENNA__07217__A2 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09611__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13386_ clknet_leaf_54_clk _00196_ net1180 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10598_ screen.register.currentYbus\[9\] screen.register.currentYbus\[8\] screen.register.currentYbus\[11\]
+ screen.register.currentYbus\[10\] vssd1 vssd1 vccd1 vccd1 _05419_ sky130_fd_sc_hd__or4_1
XANTENNA__10221__A1 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 SEL_O[3] sky130_fd_sc_hd__buf_2
X_12337_ net226 _05638_ net895 vssd1 vssd1 vccd1 vccd1 _06307_ sky130_fd_sc_hd__o21ai_1
Xoutput119 net119 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__buf_2
XFILLER_99_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12268_ net634 _04840_ vssd1 vssd1 vccd1 vccd1 _06257_ sky130_fd_sc_hd__or2_1
XANTENNA__08178__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14007_ clknet_leaf_109_clk screen.screenEdge.enableIn net1220 vssd1 vssd1 vccd1
+ vccd1 screen.screenEdge.enable1 sky130_fd_sc_hd__dfrtp_1
X_11219_ net267 net2583 net528 vssd1 vssd1 vccd1 vccd1 _00269_ sky130_fd_sc_hd__mux2_1
XFILLER_110_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12199_ screen.counter.currentCt\[3\] _06209_ vssd1 vssd1 vccd1 vccd1 _06210_ sky130_fd_sc_hd__and2_1
Xoutput90 net90 vssd1 vssd1 vccd1 vccd1 DAT_O[25] sky130_fd_sc_hd__buf_2
XANTENNA__07925__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09390__A2 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06760_ mmio.memload_or_instruction\[27\] net1050 net1017 vssd1 vssd1 vccd1 vccd1
+ _01597_ sky130_fd_sc_hd__and3_2
XFILLER_49_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12277__A2 _06254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06691_ _01459_ _01460_ datapath.ru.latched_instruction\[3\] vssd1 vssd1 vccd1 vccd1
+ _01530_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_65_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08430_ datapath.rf.registers\[0\]\[2\] net783 vssd1 vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__nor2_1
X_08361_ _03191_ _03194_ _03195_ _03196_ vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__or4_1
X_07312_ datapath.rf.registers\[6\]\[24\] net824 net813 datapath.rf.registers\[23\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__a22o_1
X_08292_ net464 _03125_ vssd1 vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__nand2_1
X_07243_ datapath.rf.registers\[19\]\[26\] net730 net687 datapath.rf.registers\[31\]\[26\]
+ _02078_ vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_30_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06833__B net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11231__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout129_A _06369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07174_ datapath.rf.registers\[30\]\[27\] net833 net817 datapath.rf.registers\[7\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__a22o_1
XFILLER_11_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09602__B1 _03770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1038_A net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10763__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08169__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13158__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout302 net305 vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__clkbuf_2
Xfanout313 _05905_ vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07664__B net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout324 _03674_ vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__buf_2
XFILLER_143_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout335 net336 vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1205_A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07916__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout346 net348 vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__buf_2
XANTENNA_input3_A DAT_I[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09815_ _03642_ net347 _04220_ net649 vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__o31a_1
Xfanout357 net358 vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__buf_2
Xfanout368 net369 vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12997__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout379 net381 vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__buf_2
XANTENNA_fanout665_A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09746_ _04564_ _04580_ vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__or2_1
XFILLER_100_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06958_ net963 net910 net908 vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__and3_2
XFILLER_86_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10279__A1 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09677_ _03604_ _04497_ _04511_ _04512_ net616 vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout832_A net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06889_ _01630_ _01638_ net988 vssd1 vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_38_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_915 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08495__B net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11406__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08628_ _02170_ _02190_ vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_124_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07695__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08559_ datapath.rf.registers\[12\]\[0\] net969 net913 _01795_ vssd1 vssd1 vccd1
+ vccd1 _03395_ sky130_fd_sc_hd__and4_1
XFILLER_30_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout718_X net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11930__A _02189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11570_ net1008 _05760_ vssd1 vssd1 vccd1 vccd1 _05794_ sky130_fd_sc_hd__or2_2
XFILLER_11_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10521_ _05329_ _05350_ vssd1 vssd1 vccd1 vccd1 _05351_ sky130_fd_sc_hd__nor2_1
XFILLER_11_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11141__S net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13240_ clknet_leaf_6_clk _00050_ net1067 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[7\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10452_ _05074_ _05285_ _05286_ vssd1 vssd1 vccd1 vccd1 _05287_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07558__C net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10980__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13171_ net2058 vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__clkbuf_1
X_10383_ _03383_ net443 _05218_ vssd1 vssd1 vccd1 vccd1 _05219_ sky130_fd_sc_hd__a21o_1
X_12122_ net1270 screen.counter.ct\[18\] _06158_ vssd1 vssd1 vccd1 vccd1 _06159_ sky130_fd_sc_hd__and3_1
XANTENNA__07080__B1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13068__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12053_ _05343_ _05824_ _06021_ _06093_ vssd1 vssd1 vccd1 vccd1 _06094_ sky130_fd_sc_hd__a211o_1
XFILLER_77_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07907__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11004_ net209 net1585 net540 vssd1 vssd1 vccd1 vccd1 _00066_ sky130_fd_sc_hd__mux2_1
XFILLER_120_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_144_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout880 net881 vssd1 vssd1 vccd1 vccd1 net880 sky130_fd_sc_hd__clkbuf_4
XFILLER_19_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout891 net896 vssd1 vssd1 vccd1 vccd1 net891 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06758__X _01595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08686__A _02660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12259__A2 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12955_ net194 net2396 net394 vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__mux2_1
XFILLER_80_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08332__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06918__B net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11316__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11906_ _02587_ net657 vssd1 vssd1 vccd1 vccd1 _05968_ sky130_fd_sc_hd__nand2_1
XFILLER_45_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10220__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12886_ net205 net2452 net398 vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__mux2_1
XFILLER_45_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14625_ clknet_leaf_45_clk _01330_ net1148 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11837_ screen.counter.ct\[6\] screen.counter.ct\[14\] screen.counter.ct\[15\] net1278
+ vssd1 vssd1 vccd1 vccd1 _05916_ sky130_fd_sc_hd__or4bb_1
XANTENNA__07438__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14556_ clknet_leaf_8_clk _01261_ net1071 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11768_ net1501 net145 net140 _02002_ vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_60_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10442__A1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13507_ clknet_leaf_120_clk _00317_ net1193 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10719_ net1556 net572 vssd1 vssd1 vccd1 vccd1 _05512_ sky130_fd_sc_hd__nor2_1
X_14487_ clknet_leaf_129_clk _01192_ net1209 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11699_ _05072_ _05885_ net149 net1423 vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__11051__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13438_ clknet_leaf_148_clk _00248_ net1061 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_155_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13369_ clknet_leaf_10_clk _00179_ net1080 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07930_ _02764_ _02765_ vssd1 vssd1 vccd1 vccd1 _02766_ sky130_fd_sc_hd__or2_1
XFILLER_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07861_ datapath.rf.registers\[4\]\[13\] net865 _02694_ _02695_ _02696_ vssd1 vssd1
+ vccd1 vccd1 _02697_ sky130_fd_sc_hd__a2111o_1
X_09600_ net358 _04244_ _04250_ net345 vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__a31o_1
XANTENNA__08571__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06812_ datapath.ru.latched_instruction\[10\] net1029 _01568_ _01490_ vssd1 vssd1
+ vccd1 vccd1 _01648_ sky130_fd_sc_hd__o2bb2a_1
X_07792_ datapath.rf.registers\[24\]\[15\] net767 net706 datapath.rf.registers\[10\]\[15\]
+ _02627_ vssd1 vssd1 vccd1 vccd1 _02628_ sky130_fd_sc_hd__a221o_1
XANTENNA__08596__A _02913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09531_ _03263_ _03296_ net623 vssd1 vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__a21oi_1
XFILLER_83_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06743_ net1002 net1018 _01581_ net1026 datapath.ru.latched_instruction\[0\] vssd1
+ vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__a32o_1
XFILLER_25_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11226__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08323__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09462_ net607 _04274_ net555 vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__o21a_1
X_06674_ net1288 net1283 mmio.memload_or_instruction\[14\] vssd1 vssd1 vccd1 vccd1
+ _01513_ sky130_fd_sc_hd__or3b_4
XTAP_TAPCELL_ROW_35_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08413_ datapath.rf.registers\[30\]\[2\] net834 _03233_ _03243_ _03245_ vssd1 vssd1
+ vccd1 vccd1 _03249_ sky130_fd_sc_hd__a2111o_1
X_09393_ _04152_ _04228_ net369 vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout246_A _05599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08344_ datapath.rf.registers\[9\]\[3\] net986 net943 vssd1 vssd1 vccd1 vccd1 _03180_
+ sky130_fd_sc_hd__and3_1
XFILLER_149_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07429__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09823__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10433__A1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08275_ datapath.rf.registers\[11\]\[5\] net711 net661 datapath.rf.registers\[5\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03111_ sky130_fd_sc_hd__a22o_1
XANTENNA__07659__B net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout413_A _05730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1155_A net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07226_ datapath.rf.registers\[6\]\[26\] net824 net815 datapath.rf.registers\[21\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__a22o_1
XFILLER_153_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07157_ datapath.rf.registers\[22\]\[28\] net736 _01832_ datapath.rf.registers\[21\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01993_ sky130_fd_sc_hd__a22o_1
XANTENNA__10197__B1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11909__B net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07088_ datapath.rf.registers\[4\]\[29\] net864 net821 datapath.rf.registers\[22\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout782_A net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1108 net1109 vssd1 vssd1 vccd1 vccd1 net1108 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1110_X net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1119 net1120 vssd1 vssd1 vccd1 vccd1 net1119 sky130_fd_sc_hd__clkbuf_2
XFILLER_102_931 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout132 net133 vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__clkbuf_2
Xfanout143 net147 vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__buf_2
Xfanout154 net155 vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__buf_2
Xfanout165 _05288_ vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout668_X net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout176 _05670_ vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08002__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout187 net188 vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_126_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout198 _05653_ vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__clkbuf_2
XFILLER_28_720 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09729_ _03439_ _03529_ vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout835_X net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11136__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12740_ net2084 net275 net404 vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__mux2_1
XFILLER_16_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08865__A1 _02661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12671_ net499 _06505_ _06506_ net503 net2612 vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__a32o_1
XANTENNA__10975__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14410_ clknet_leaf_58_clk _01115_ net1167 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[2\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11622_ _05736_ net1010 vssd1 vssd1 vccd1 vccd1 _05846_ sky130_fd_sc_hd__or2_2
XFILLER_30_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14341_ clknet_leaf_139_clk _01046_ net1099 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11553_ _05750_ _05763_ vssd1 vssd1 vccd1 vccd1 _05777_ sky130_fd_sc_hd__or2_2
XANTENNA__08093__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10504_ _05316_ screen.controlBus\[7\] screen.controlBus\[6\] vssd1 vssd1 vccd1 vccd1
+ _05334_ sky130_fd_sc_hd__or3b_1
XFILLER_156_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14272_ clknet_leaf_138_clk _00977_ net1097 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07840__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11484_ net291 net1599 net510 vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_137_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13223_ clknet_leaf_143_clk _00033_ net1086 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire588 _02703_ vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__clkbuf_1
X_10435_ _05211_ _05240_ _05270_ vssd1 vssd1 vccd1 vccd1 _05271_ sky130_fd_sc_hd__nor3_1
XFILLER_137_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07053__B1 _01887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13154_ net1949 net194 net383 vssd1 vssd1 vccd1 vccd1 _01395_ sky130_fd_sc_hd__mux2_1
X_10366_ _05095_ _05200_ _05201_ vssd1 vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__nor3_1
XFILLER_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12105_ _06134_ _06142_ net1011 vssd1 vssd1 vccd1 vccd1 _06143_ sky130_fd_sc_hd__o21ai_1
X_13085_ net1571 net203 net386 vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__mux2_1
X_10297_ _04841_ _04842_ vssd1 vssd1 vccd1 vccd1 _05133_ sky130_fd_sc_hd__or2_1
XFILLER_151_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12036_ screen.register.currentXbus\[27\] _05772_ _06076_ _06077_ vssd1 vssd1 vccd1
+ vccd1 _06078_ sky130_fd_sc_hd__a211o_1
XFILLER_38_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06929__A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13987_ clknet_leaf_108_clk _00764_ net1219 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08305__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11046__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12938_ net276 net2581 net396 vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__mux2_1
XFILLER_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12869_ net292 net2349 net398 vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__mux2_1
X_14608_ clknet_leaf_23_clk _01313_ net1155 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12385__B net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10415__A1 _03321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09281__A1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14539_ clknet_leaf_55_clk _01244_ net1173 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08084__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10966__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07292__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08060_ datapath.rf.registers\[4\]\[9\] net959 net934 vssd1 vssd1 vccd1 vccd1 _02896_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07831__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07011_ datapath.rf.registers\[1\]\[31\] net762 _01846_ net786 vssd1 vssd1 vccd1
+ vccd1 _01847_ sky130_fd_sc_hd__a211o_1
XANTENNA__07044__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08792__A0 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08962_ _03793_ _03797_ net341 vssd1 vssd1 vccd1 vccd1 _03798_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_90_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07913_ _02735_ _02743_ _02746_ _02748_ vssd1 vssd1 vccd1 vccd1 _02749_ sky130_fd_sc_hd__nor4_1
X_08893_ datapath.i_ack datapath.pc_module.i_ack2 vssd1 vssd1 vccd1 vccd1 _03729_
+ sky130_fd_sc_hd__and2b_1
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08544__B1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout196_A _05653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09741__C1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07844_ datapath.rf.registers\[0\]\[14\] net784 _02676_ _02679_ vssd1 vssd1 vccd1
+ vccd1 _02680_ sky130_fd_sc_hd__o22a_4
XANTENNA__07942__B net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10351__B1 net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07898__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07775_ datapath.rf.registers\[6\]\[15\] net824 _02602_ _02606_ _02610_ vssd1 vssd1
+ vccd1 vccd1 _02611_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07661__C net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09514_ net552 net548 _02750_ vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__a21o_1
XFILLER_83_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06726_ _01406_ datapath.multiplication_module.mul_prev datapath.ru.n_memread datapath.ru.n_memwrite
+ vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_88_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08847__A1 _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09502__X _04338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09445_ _04278_ _04279_ net454 vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06858__B1 _01614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06657_ mmio.memload_or_instruction\[31\] net1050 datapath.ru.latched_instruction\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01496_ sky130_fd_sc_hd__a21bo_1
XFILLER_13_918 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10795__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout530_A net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout628_A net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08773__B net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09221__Y _04057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09376_ net609 _04208_ vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__nand2_1
X_06588_ datapath.mulitply_result\[30\] vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__inv_2
X_08327_ datapath.rf.registers\[4\]\[4\] net715 net706 datapath.rf.registers\[10\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__a22o_1
XFILLER_137_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout416_X net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08258_ datapath.rf.registers\[19\]\[5\] net853 net795 datapath.rf.registers\[31\]\[5\]
+ _03083_ vssd1 vssd1 vccd1 vccd1 _03094_ sky130_fd_sc_hd__a221o_1
XANTENNA__07822__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07209_ datapath.rf.registers\[0\]\[27\] net784 net591 _02044_ vssd1 vssd1 vccd1
+ vccd1 _02045_ sky130_fd_sc_hd__a2bb2o_2
Xteam_04_1330 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] team_04_1330/LO sky130_fd_sc_hd__conb_1
X_08189_ datapath.rf.registers\[28\]\[7\] net752 net704 datapath.rf.registers\[9\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03025_ sky130_fd_sc_hd__a22o_1
Xteam_04_1341 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] team_04_1341/LO sky130_fd_sc_hd__conb_1
X_10220_ datapath.PC\[29\] _04645_ net469 vssd1 vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__mux2_1
XFILLER_3_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout785_X net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08783__A0 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10151_ _04983_ _04986_ net1263 net1259 vssd1 vssd1 vccd1 vccd1 _04987_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_58_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10082_ net229 _04917_ net1258 vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout952_X net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08535__B1 _01768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13910_ clknet_leaf_42_clk net1370 net1149 vssd1 vssd1 vccd1 vccd1 keypad.debounce.debounce\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07889__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06749__A _01585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10893__A1 datapath.mulitply_result\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09125__A _02169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_807 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13841_ clknet_leaf_113_clk _00650_ net1195 vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10893__B2 _05639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12189__C net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13772_ clknet_leaf_83_clk _00581_ net1260 vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12095__B1 _05786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10984_ net2128 net247 net434 vssd1 vssd1 vccd1 vccd1 _00049_ sky130_fd_sc_hd__mux2_1
X_12723_ columns.count\[8\] _06541_ vssd1 vssd1 vccd1 vccd1 _06545_ sky130_fd_sc_hd__nand2_1
XFILLER_15_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13081__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12654_ datapath.mulitply_result\[24\] datapath.multiplication_module.multiplicand_i\[24\]
+ vssd1 vssd1 vccd1 vccd1 _06492_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_139_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11605_ _05799_ _05826_ _05828_ vssd1 vssd1 vccd1 vccd1 _05829_ sky130_fd_sc_hd__nor3_1
XANTENNA__08066__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12585_ net2195 net504 net500 _06434_ vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__a22o_1
X_11536_ _05293_ _05750_ vssd1 vssd1 vccd1 vccd1 _05760_ sky130_fd_sc_hd__or2_2
X_14324_ clknet_leaf_128_clk _01029_ net1117 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07813__A2 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14255_ clknet_leaf_27_clk _00960_ net1134 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11467_ net1732 net205 net406 vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__mux2_1
XFILLER_125_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13206_ clknet_leaf_142_clk _00016_ net1093 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_99_73 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10418_ net353 _04434_ _05253_ net359 vssd1 vssd1 vccd1 vccd1 _05254_ sky130_fd_sc_hd__o211a_1
X_14186_ clknet_leaf_55_clk _00941_ net1179 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_125_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11398_ net1634 net214 net410 vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__mux2_1
XANTENNA__10453__B _05073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08774__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13137_ net2078 net276 net384 vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__mux2_1
X_10349_ _04835_ _04851_ vssd1 vssd1 vccd1 vccd1 _05185_ sky130_fd_sc_hd__nand2_1
XFILLER_140_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13068_ net2558 net290 net386 vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__mux2_1
XANTENNA__12322__B2 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12019_ screen.register.currentYbus\[2\] _05778_ net997 screen.register.currentXbus\[18\]
+ vssd1 vssd1 vccd1 vccd1 _06062_ sky130_fd_sc_hd__a22o_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08577__C _01831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12086__B1 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07560_ datapath.rf.registers\[23\]\[19\] net942 net924 vssd1 vssd1 vccd1 vccd1 _02396_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08829__A1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06946__X _01782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07491_ datapath.rf.registers\[3\]\[21\] net770 net706 datapath.rf.registers\[10\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__a22o_1
XFILLER_62_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11504__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09230_ net372 _04064_ _04065_ vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_14_Left_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09161_ net459 _03994_ _03995_ vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__nand3_1
XANTENNA__09254__A1 _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08112_ datapath.rf.registers\[2\]\[8\] net889 net838 datapath.rf.registers\[26\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02948_ sky130_fd_sc_hd__a22o_1
X_09092_ _03926_ _03927_ vssd1 vssd1 vccd1 vccd1 _03928_ sky130_fd_sc_hd__nand2_1
XFILLER_119_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08043_ net611 _02876_ _02878_ vssd1 vssd1 vccd1 vccd1 _02879_ sky130_fd_sc_hd__o21ai_1
XFILLER_147_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold900 datapath.rf.registers\[28\]\[24\] vssd1 vssd1 vccd1 vccd1 net2248 sky130_fd_sc_hd__dlygate4sd3_1
Xhold911 datapath.rf.registers\[16\]\[7\] vssd1 vssd1 vccd1 vccd1 net2259 sky130_fd_sc_hd__dlygate4sd3_1
Xhold922 datapath.rf.registers\[4\]\[26\] vssd1 vssd1 vccd1 vccd1 net2270 sky130_fd_sc_hd__dlygate4sd3_1
Xhold933 datapath.rf.registers\[6\]\[27\] vssd1 vssd1 vccd1 vccd1 net2281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold944 datapath.rf.registers\[2\]\[5\] vssd1 vssd1 vccd1 vccd1 net2292 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07656__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold955 datapath.rf.registers\[24\]\[10\] vssd1 vssd1 vccd1 vccd1 net2303 sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 datapath.rf.registers\[21\]\[12\] vssd1 vssd1 vccd1 vccd1 net2314 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12561__A1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold977 datapath.rf.registers\[30\]\[31\] vssd1 vssd1 vccd1 vccd1 net2325 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Left_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09994_ _04820_ _04722_ vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout1020_A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold988 datapath.rf.registers\[9\]\[26\] vssd1 vssd1 vccd1 vccd1 net2336 sky130_fd_sc_hd__dlygate4sd3_1
Xhold999 datapath.rf.registers\[21\]\[5\] vssd1 vssd1 vccd1 vccd1 net2347 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08945_ _02264_ _02311_ net445 vssd1 vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout480_A _06556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout578_A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08876_ net559 net558 net446 vssd1 vssd1 vccd1 vccd1 _03712_ sky130_fd_sc_hd__mux2_1
XANTENNA__10324__B1 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07827_ datapath.rf.registers\[11\]\[14\] net711 net707 datapath.rf.registers\[10\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02663_ sky130_fd_sc_hd__a22o_1
XFILLER_57_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07758_ datapath.rf.registers\[29\]\[15\] net975 net917 vssd1 vssd1 vccd1 vccd1 _02594_
+ sky130_fd_sc_hd__and3_1
X_06709_ datapath.ru.latched_instruction\[8\] datapath.ru.latched_instruction\[9\]
+ datapath.ru.latched_instruction\[10\] datapath.ru.latched_instruction\[11\] vssd1
+ vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__or4_1
XFILLER_71_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08296__A2 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09493__A1 _01603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07689_ datapath.rf.registers\[22\]\[17\] net736 net670 datapath.rf.registers\[21\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02525_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout533_X net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11414__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09428_ net574 _04254_ _04255_ _04263_ vssd1 vssd1 vccd1 vccd1 _04264_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_23_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09359_ net557 net577 net546 _02612_ vssd1 vssd1 vccd1 vccd1 _04195_ sky130_fd_sc_hd__o211ai_1
XANTENNA_fanout700_X net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09245__A1 _01620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12370_ net634 _05237_ vssd1 vssd1 vccd1 vccd1 _06331_ sky130_fd_sc_hd__and2_1
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11321_ net2206 net264 net415 vssd1 vssd1 vccd1 vccd1 _00366_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07008__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14040_ clknet_leaf_87_clk _00809_ net1253 vssd1 vssd1 vccd1 vccd1 datapath.PC\[30\]
+ sky130_fd_sc_hd__dfrtp_4
X_11252_ net268 net1647 net420 vssd1 vssd1 vccd1 vccd1 _00301_ sky130_fd_sc_hd__mux2_1
XFILLER_4_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07566__C net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10203_ _04605_ _05038_ vssd1 vssd1 vccd1 vccd1 _05039_ sky130_fd_sc_hd__or2_1
XFILLER_106_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11183_ net276 net2175 net424 vssd1 vssd1 vccd1 vccd1 _00235_ sky130_fd_sc_hd__mux2_1
XFILLER_121_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10134_ _03729_ _04969_ _04968_ net640 vssd1 vssd1 vccd1 vccd1 _04970_ sky130_fd_sc_hd__a211o_1
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13076__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10065_ _04894_ _04895_ _04896_ vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_50_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08397__C net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12068__B1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13824_ clknet_leaf_112_clk _00633_ net1197 vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__dfrtp_1
XANTENNA__06766__X _01603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09142__X _03978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13755_ clknet_leaf_76_clk _00564_ net1248 vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09484__A1 _02961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10967_ net1541 net259 net436 vssd1 vssd1 vccd1 vccd1 _00035_ sky130_fd_sc_hd__mux2_1
XFILLER_43_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11324__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12706_ columns.count\[1\] columns.count\[0\] columns.count\[2\] _06531_ vssd1 vssd1
+ vccd1 vccd1 _06534_ sky130_fd_sc_hd__and4_1
XANTENNA__07495__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10898_ net903 _03950_ _05643_ vssd1 vssd1 vccd1 vccd1 _05644_ sky130_fd_sc_hd__o21ai_4
X_13686_ clknet_leaf_141_clk _00496_ net1095 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_12637_ datapath.mulitply_result\[21\] datapath.multiplication_module.multiplicand_i\[21\]
+ vssd1 vssd1 vccd1 vccd1 _06478_ sky130_fd_sc_hd__nor2_1
XFILLER_8_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07247__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12568_ datapath.mulitply_result\[10\] datapath.multiplication_module.multiplicand_i\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06420_ sky130_fd_sc_hd__nand2_1
XFILLER_8_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_152_Right_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11519_ _05346_ _05739_ _05740_ vssd1 vssd1 vccd1 vccd1 _05744_ sky130_fd_sc_hd__and3_1
X_14307_ clknet_leaf_121_clk _01012_ net1200 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07757__B net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12499_ net214 net2448 net506 vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__mux2_1
XFILLER_8_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold207 datapath.rf.registers\[29\]\[1\] vssd1 vssd1 vccd1 vccd1 net1555 sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 datapath.rf.registers\[20\]\[24\] vssd1 vssd1 vccd1 vccd1 net1566 sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 datapath.rf.registers\[28\]\[0\] vssd1 vssd1 vccd1 vccd1 net1577 sky130_fd_sc_hd__dlygate4sd3_1
X_14238_ clknet_leaf_123_clk datapath.multiplication_module.multiplier_i_n\[6\] net1214
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i\[6\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12543__A1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14169_ clknet_leaf_54_clk _00924_ net1180 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08211__A2 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout709 _01818_ vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08221__X _03057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06991_ net966 _01816_ vssd1 vssd1 vccd1 vccd1 _01827_ sky130_fd_sc_hd__and2_1
XFILLER_86_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08730_ _03564_ _03565_ _03539_ vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09172__A0 _03796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1280 screen.counter.ct\[4\] vssd1 vssd1 vccd1 vccd1 net1280 sky130_fd_sc_hd__buf_2
Xfanout1291 net72 vssd1 vssd1 vccd1 vccd1 net1291 sky130_fd_sc_hd__clkbuf_2
X_08661_ _02191_ _03464_ vssd1 vssd1 vccd1 vccd1 _03497_ sky130_fd_sc_hd__or2_2
XFILLER_39_689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07612_ datapath.rf.registers\[27\]\[18\] net974 net939 vssd1 vssd1 vccd1 vccd1 _02448_
+ sky130_fd_sc_hd__and3_1
X_08592_ _03128_ _03426_ _03427_ vssd1 vssd1 vccd1 vccd1 _03428_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_85_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07543_ datapath.rf.registers\[4\]\[20\] net714 net660 datapath.rf.registers\[5\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _02379_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_101_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11234__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout159_A _06335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07486__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07474_ _02302_ _02306_ _02307_ _02309_ vssd1 vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__nor4_1
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09213_ net337 _04048_ vssd1 vssd1 vccd1 vccd1 _04049_ sky130_fd_sc_hd__nor2_1
XANTENNA__09227__A1 _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10926__X _05668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07238__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1068_A net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09144_ _03504_ _03585_ _03502_ vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__a21oi_1
XFILLER_30_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08986__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07667__B net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09075_ _03910_ vssd1 vssd1 vccd1 vccd1 _03911_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_116_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08450__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08026_ datapath.rf.registers\[17\]\[10\] net748 net724 datapath.rf.registers\[18\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__a22o_1
Xhold730 datapath.rf.registers\[6\]\[9\] vssd1 vssd1 vccd1 vccd1 net2078 sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 datapath.rf.registers\[21\]\[1\] vssd1 vssd1 vccd1 vccd1 net2089 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout695_A net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold752 datapath.rf.registers\[17\]\[8\] vssd1 vssd1 vccd1 vccd1 net2100 sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 datapath.rf.registers\[10\]\[20\] vssd1 vssd1 vccd1 vccd1 net2111 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09882__B net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold774 datapath.rf.registers\[22\]\[8\] vssd1 vssd1 vccd1 vccd1 net2122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold785 datapath.rf.registers\[8\]\[7\] vssd1 vssd1 vccd1 vccd1 net2133 sky130_fd_sc_hd__dlygate4sd3_1
Xhold796 datapath.rf.registers\[26\]\[31\] vssd1 vssd1 vccd1 vccd1 net2144 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07410__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09977_ _04729_ _04812_ _04730_ vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout483_X net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout862_A net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08498__B net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08928_ net364 _03763_ vssd1 vssd1 vccd1 vccd1 _03764_ sky130_fd_sc_hd__nand2_1
XFILLER_85_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout650_X net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08859_ _03694_ _03685_ net451 vssd1 vssd1 vccd1 vccd1 _03695_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout748_X net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11933__A _02145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11870_ _03170_ net656 vssd1 vssd1 vccd1 vccd1 _05944_ sky130_fd_sc_hd__nand2_1
XFILLER_72_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10821_ _05576_ _05577_ vssd1 vssd1 vccd1 vccd1 _05578_ sky130_fd_sc_hd__or2_1
XANTENNA__11652__B _05874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08269__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout915_X net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11144__S net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07477__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13540_ clknet_leaf_19_clk _00350_ net1109 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10752_ _05515_ _05518_ vssd1 vssd1 vccd1 vccd1 _05519_ sky130_fd_sc_hd__or2_1
X_13471_ clknet_leaf_17_clk _00281_ net1106 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10683_ keypad.alpha _05496_ _05499_ _05500_ vssd1 vssd1 vccd1 vccd1 keypad.decode.button_n\[2\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10983__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09218__A1 _01620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07229__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12422_ net1386 net130 _06358_ vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__a21o_1
XFILLER_138_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12353_ net893 _03865_ _06317_ _06318_ net306 vssd1 vssd1 vccd1 vccd1 _06319_ sky130_fd_sc_hd__o221a_1
XFILLER_126_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08441__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10784__B1 _05545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11304_ net174 net1581 net524 vssd1 vssd1 vccd1 vccd1 _00352_ sky130_fd_sc_hd__mux2_1
X_12284_ net634 _04847_ vssd1 vssd1 vccd1 vccd1 _06269_ sky130_fd_sc_hd__nor2_1
X_14023_ clknet_leaf_76_clk _00792_ net1249 vssd1 vssd1 vccd1 vccd1 datapath.PC\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_4_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11235_ net187 net1744 net527 vssd1 vssd1 vccd1 vccd1 _00285_ sky130_fd_sc_hd__mux2_1
XANTENNA__08689__A _02705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11166_ net197 net2603 net532 vssd1 vssd1 vccd1 vccd1 _00219_ sky130_fd_sc_hd__mux2_1
XANTENNA__11319__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10117_ net225 _04952_ net1294 vssd1 vssd1 vccd1 vccd1 _04953_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_147_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12289__B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11097_ net199 net1759 net534 vssd1 vssd1 vccd1 vccd1 _00154_ sky130_fd_sc_hd__mux2_1
XANTENNA__08201__B net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10048_ _04822_ _04883_ vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__xnor2_1
XFILLER_64_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold90 net113 vssd1 vssd1 vccd1 vccd1 net1438 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07180__A2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13807_ clknet_leaf_73_clk _00616_ net1243 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_63_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11999_ _05741_ _05793_ _06042_ _05320_ _06024_ vssd1 vssd1 vccd1 vccd1 _06043_ sky130_fd_sc_hd__a221o_1
XANTENNA__11054__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08114__D1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09032__B _03867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07468__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13738_ clknet_leaf_103_clk _00548_ net1225 vssd1 vssd1 vccd1 vccd1 screen.screenLogic.currentWrx
+ sky130_fd_sc_hd__dfstp_1
XFILLER_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09209__A1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13669_ clknet_leaf_114_clk _00479_ net1190 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06943__Y _01779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07190_ _02025_ vssd1 vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__inv_2
XFILLER_118_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12393__B net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12961__X _06556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_756 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09900_ _04735_ vssd1 vssd1 vccd1 vccd1 _04736_ sky130_fd_sc_hd__inv_2
Xfanout506 net509 vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_111_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09831_ _03477_ _03478_ _04666_ vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__a21oi_1
Xfanout517 _05731_ vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__clkbuf_4
Xfanout528 _05721_ vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__clkbuf_8
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout539 net541 vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__buf_4
XFILLER_113_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload13_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06746__A2 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11229__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06974_ net963 net910 _01809_ vssd1 vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__and3_1
X_09762_ _01619_ _03513_ _04597_ vssd1 vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__a21bo_1
XANTENNA__09145__B1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08713_ _03547_ _03548_ _03546_ vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__a21o_1
X_09693_ net574 _04523_ _04524_ _04528_ vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__a22o_1
XFILLER_82_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07950__B net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08644_ _01706_ _03479_ vssd1 vssd1 vccd1 vccd1 _03480_ sky130_fd_sc_hd__or2_1
XFILLER_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08765__C _01604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08575_ datapath.rf.registers\[6\]\[0\] net682 _03408_ _03409_ _03410_ vssd1 vssd1
+ vccd1 vccd1 _03411_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10369__A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1185_A net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07459__B1 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07526_ _02359_ _02360_ _02361_ vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__or3_1
XFILLER_23_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07457_ datapath.rf.registers\[8\]\[21\] net876 net849 datapath.rf.registers\[17\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__a22o_1
XFILLER_50_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout610_A _01782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout708_A net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06682__B2 datapath.ru.latched_instruction\[29\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07388_ datapath.rf.registers\[14\]\[23\] net774 net687 datapath.rf.registers\[31\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__a22o_1
X_09127_ _03961_ _03962_ net454 vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_98_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08423__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09058_ _03688_ _03690_ net449 vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout698_X net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08009_ datapath.rf.registers\[13\]\[10\] net812 _02833_ _02839_ _02842_ vssd1 vssd1
+ vccd1 vccd1 _02845_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08005__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold560 datapath.rf.registers\[17\]\[28\] vssd1 vssd1 vccd1 vccd1 net1908 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold571 datapath.rf.registers\[4\]\[28\] vssd1 vssd1 vccd1 vccd1 net1919 sky130_fd_sc_hd__dlygate4sd3_1
X_11020_ net245 net2327 net538 vssd1 vssd1 vccd1 vccd1 _00082_ sky130_fd_sc_hd__mux2_1
Xhold582 datapath.rf.registers\[4\]\[16\] vssd1 vssd1 vccd1 vccd1 net1930 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold593 datapath.rf.registers\[15\]\[23\] vssd1 vssd1 vccd1 vccd1 net1941 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout865_X net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11730__A2 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_129_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12971_ net275 net2214 net480 vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__mux2_1
XANTENNA__10978__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1260 datapath.rf.registers\[18\]\[15\] vssd1 vssd1 vccd1 vccd1 net2608 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1271 datapath.rf.registers\[14\]\[9\] vssd1 vssd1 vccd1 vccd1 net2619 sky130_fd_sc_hd__dlygate4sd3_1
X_11922_ net134 _05978_ _05977_ vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__o21ai_1
Xhold1282 screen.register.currentYbus\[27\] vssd1 vssd1 vccd1 vccd1 net2630 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07698__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1293 datapath.rf.registers\[3\]\[31\] vssd1 vssd1 vccd1 vccd1 net2641 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07162__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14641_ clknet_leaf_34_clk _01346_ net1127 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11853_ _05281_ _05283_ vssd1 vssd1 vccd1 vccd1 _05931_ sky130_fd_sc_hd__nor2_1
XFILLER_60_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10804_ _01490_ net620 _05562_ _05563_ vssd1 vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__o2bb2a_2
X_11784_ _05897_ _05896_ net2655 vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__mux2_1
X_14572_ clknet_leaf_16_clk _01277_ net1104 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08972__A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13523_ clknet_leaf_34_clk _00333_ net1128 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10735_ net1709 net568 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[21\]
+ sky130_fd_sc_hd__and2_1
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06673__A1 datapath.ru.latched_instruction\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__06673__B2 datapath.ru.latched_instruction\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10666_ _05471_ _05484_ vssd1 vssd1 vccd1 vccd1 _05485_ sky130_fd_sc_hd__nor2_1
XFILLER_139_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13454_ clknet_leaf_5_clk _00264_ net1068 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07870__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12405_ _05962_ net156 vssd1 vssd1 vccd1 vccd1 _06350_ sky130_fd_sc_hd__nor2_1
X_13385_ clknet_leaf_91_clk _00195_ net1232 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10597_ screen.register.currentYbus\[1\] screen.register.currentYbus\[0\] screen.register.currentYbus\[3\]
+ screen.register.currentYbus\[2\] vssd1 vssd1 vccd1 vccd1 _05418_ sky130_fd_sc_hd__or4_1
XANTENNA__09611__A1 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08414__A2 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 STB_O sky130_fd_sc_hd__buf_2
X_12336_ net230 _04880_ vssd1 vssd1 vccd1 vccd1 _06306_ sky130_fd_sc_hd__nor2_1
XFILLER_56_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12267_ net891 _04428_ vssd1 vssd1 vccd1 vccd1 _06256_ sky130_fd_sc_hd__or2_1
XFILLER_141_247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14006_ clknet_leaf_107_clk net1363 net1220 vssd1 vssd1 vccd1 vccd1 screen.screenEdge.enable3
+ sky130_fd_sc_hd__dfrtp_1
X_11218_ net272 net2469 net528 vssd1 vssd1 vccd1 vccd1 _00268_ sky130_fd_sc_hd__mux2_1
XANTENNA__09375__B1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12198_ _06168_ _06208_ _06209_ vssd1 vssd1 vccd1 vccd1 _00760_ sky130_fd_sc_hd__nor3_1
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 DAT_O[16] sky130_fd_sc_hd__buf_2
Xoutput91 net91 vssd1 vssd1 vccd1 vccd1 DAT_O[26] sky130_fd_sc_hd__buf_2
XANTENNA__11049__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11149_ net280 net2186 net532 vssd1 vssd1 vccd1 vccd1 _00202_ sky130_fd_sc_hd__mux2_1
XFILLER_110_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07689__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06690_ mmio.memload_or_instruction\[5\] net1051 _01440_ _01411_ vssd1 vssd1 vccd1
+ vccd1 _01529_ sky130_fd_sc_hd__a211oi_1
XFILLER_36_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07153__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06900__A2 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08360_ datapath.rf.registers\[23\]\[3\] net814 _03175_ _03177_ _03188_ vssd1 vssd1
+ vccd1 vccd1 _03196_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08882__A _01610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07311_ _02125_ _02146_ vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__and2_1
X_08291_ net464 _03125_ vssd1 vssd1 vccd1 vccd1 _03127_ sky130_fd_sc_hd__nor2_1
X_07242_ datapath.rf.registers\[11\]\[26\] net710 net675 datapath.rf.registers\[29\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_30_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07173_ datapath.rf.registers\[10\]\[27\] net880 net836 datapath.rf.registers\[26\]\[27\]
+ _02008_ vssd1 vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__a221o_1
XANTENNA__09602__A1 _01609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08106__B net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07613__B1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07945__B net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout303 net305 vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__clkbuf_2
Xfanout314 _05905_ vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__clkbuf_2
Xfanout325 net326 vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07664__C net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11712__A2 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout336 _05904_ vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__clkbuf_2
XFILLER_143_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09814_ net380 _04225_ vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__nor2_1
Xfanout347 net348 vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__buf_2
Xfanout358 _03647_ vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__buf_2
Xfanout369 _03628_ vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__buf_2
XANTENNA__07392__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09745_ _04564_ _04580_ vssd1 vssd1 vccd1 vccd1 _04581_ sky130_fd_sc_hd__nor2_1
XFILLER_28_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10798__S net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout560_A _03057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06957_ _01637_ net990 vssd1 vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout658_A net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09676_ net324 _03943_ _04508_ vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__o21ai_1
X_06888_ _01707_ net955 vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__nand2_4
XANTENNA__12298__B _04580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07144__A2 _01724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_6_Left_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08627_ _02125_ _02146_ vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__or2_1
XFILLER_15_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout825_A _01753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08558_ datapath.rf.registers\[28\]\[0\] net965 net913 _01795_ vssd1 vssd1 vccd1
+ vccd1 _03394_ sky130_fd_sc_hd__and4_1
XANTENNA__11930__B net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07509_ datapath.rf.registers\[3\]\[20\] net982 net927 vssd1 vssd1 vccd1 vccd1 _02345_
+ sky130_fd_sc_hd__and3_1
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08489_ datapath.rf.registers\[29\]\[1\] net963 _01823_ vssd1 vssd1 vccd1 vccd1 _03325_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout613_X net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11422__S net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10520_ _05335_ _05343_ vssd1 vssd1 vccd1 vccd1 _05350_ sky130_fd_sc_hd__or2_1
XANTENNA__07852__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10451_ datapath.i_ack mmio.WEN2 _01576_ _01589_ vssd1 vssd1 vccd1 vccd1 _05286_
+ sky130_fd_sc_hd__nor4_1
XFILLER_136_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07604__B1 _01787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13170_ net2290 vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__clkbuf_1
X_10382_ _03320_ net440 net363 vssd1 vssd1 vccd1 vccd1 _05218_ sky130_fd_sc_hd__a21o_1
XFILLER_109_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12121_ net1271 net1272 screen.counter.ct\[16\] _06157_ vssd1 vssd1 vccd1 vccd1 _06158_
+ sky130_fd_sc_hd__and4_1
XFILLER_123_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09357__B1 _03661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12052_ _05335_ net998 _05847_ _06024_ _06073_ vssd1 vssd1 vccd1 vccd1 _06093_ sky130_fd_sc_hd__a2111o_1
Xhold390 datapath.rf.registers\[30\]\[3\] vssd1 vssd1 vccd1 vccd1 net1738 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11003_ _05517_ _05708_ vssd1 vssd1 vccd1 vccd1 _05709_ sky130_fd_sc_hd__nand2_1
XANTENNA__07383__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout870 net871 vssd1 vssd1 vccd1 vccd1 net870 sky130_fd_sc_hd__buf_4
XANTENNA__09109__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09415__X _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout881 _01721_ vssd1 vssd1 vccd1 vccd1 net881 sky130_fd_sc_hd__clkbuf_8
Xfanout892 net896 vssd1 vssd1 vccd1 vccd1 net892 sky130_fd_sc_hd__buf_2
XFILLER_19_924 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13084__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_82_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12954_ net197 net2639 net396 vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__mux2_1
Xhold1090 datapath.rf.registers\[17\]\[30\] vssd1 vssd1 vccd1 vccd1 net2438 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07135__A2 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06918__C net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11905_ screen.register.currentYbus\[16\] net162 vssd1 vssd1 vccd1 vccd1 _05967_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_47_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12885_ net210 net2316 net398 vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__mux2_1
XANTENNA__07540__C1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14624_ clknet_leaf_135_clk _01329_ net1104 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06774__X _01611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11836_ screen.counter.ct\[13\] screen.counter.ct\[12\] screen.counter.ct\[18\] screen.counter.ct\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05915_ sky130_fd_sc_hd__or4b_1
XFILLER_61_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_97_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14555_ clknet_leaf_37_clk _01260_ net1136 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_11767_ net1476 net145 net140 _02046_ vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__a22o_1
XANTENNA__11332__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_140_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13506_ clknet_leaf_151_clk _00316_ net1052 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10718_ _03104_ net572 _05511_ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[5\]
+ sky130_fd_sc_hd__a21oi_1
X_14486_ clknet_leaf_142_clk _01191_ net1093 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_11698_ _04944_ _05885_ net149 net1459 vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_155_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13437_ clknet_leaf_149_clk _00247_ net1092 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_20_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10649_ _05453_ _05464_ _05443_ _05444_ vssd1 vssd1 vccd1 vccd1 _05469_ sky130_fd_sc_hd__a2bb2o_1
X_13368_ clknet_leaf_4_clk _00178_ net1069 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06950__A net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12319_ net894 _04600_ vssd1 vssd1 vccd1 vccd1 _06294_ sky130_fd_sc_hd__nor2_1
XFILLER_5_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13299_ clknet_leaf_34_clk _00109_ net1128 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_58_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_35_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11855__X _05933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07860_ datapath.rf.registers\[1\]\[13\] net846 net817 datapath.rf.registers\[7\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02696_ sky130_fd_sc_hd__a22o_1
XANTENNA__08020__B1 _02855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07374__A2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06811_ net1004 net1020 _01645_ net1028 datapath.ru.latched_instruction\[23\] vssd1
+ vssd1 vccd1 vccd1 _01647_ sky130_fd_sc_hd__a32o_4
X_07791_ datapath.rf.registers\[28\]\[15\] net751 net661 datapath.rf.registers\[5\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__a22o_1
XFILLER_84_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11507__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06742_ datapath.ru.latched_instruction\[0\] _01500_ net1014 vssd1 vssd1 vccd1 vccd1
+ _01581_ sky130_fd_sc_hd__mux2_1
XANTENNA__11458__A1 _05588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09530_ net324 _04365_ vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__nor2_1
XANTENNA__07126__A2 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09461_ net904 _04273_ _04296_ vssd1 vssd1 vccd1 vccd1 _04297_ sky130_fd_sc_hd__o21ai_1
X_06673_ datapath.ru.latched_instruction\[30\] _01466_ _01511_ datapath.ru.latched_instruction\[15\]
+ vssd1 vssd1 vccd1 vccd1 _01512_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_35_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08412_ datapath.rf.registers\[19\]\[2\] net854 net792 datapath.rf.registers\[18\]\[2\]
+ _03244_ vssd1 vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__a221o_1
X_09392_ _02613_ _02661_ net443 vssd1 vssd1 vccd1 vccd1 _04228_ sky130_fd_sc_hd__mux2_1
XFILLER_40_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08343_ datapath.rf.registers\[30\]\[3\] net979 net919 vssd1 vssd1 vccd1 vccd1 _03179_
+ sky130_fd_sc_hd__and3_1
XFILLER_149_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout141_A net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09823__A1 _01888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_108_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11242__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07834__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08274_ datapath.rf.registers\[2\]\[5\] net743 net680 datapath.rf.registers\[6\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03110_ sky130_fd_sc_hd__a22o_1
XANTENNA__07659__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07225_ datapath.rf.registers\[28\]\[26\] net804 net790 datapath.rf.registers\[18\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02061_ sky130_fd_sc_hd__a22o_1
XFILLER_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10934__X _05675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1050_A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout406_A _05733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07156_ datapath.rf.registers\[16\]\[28\] net741 net724 datapath.rf.registers\[18\]\[28\]
+ _01989_ vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__a221o_1
XFILLER_145_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07087_ datapath.rf.registers\[6\]\[29\] net824 net817 datapath.rf.registers\[7\]\[29\]
+ _01914_ vssd1 vssd1 vccd1 vccd1 _01923_ sky130_fd_sc_hd__a221o_1
XFILLER_154_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout775_A _01796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1109 net1110 vssd1 vssd1 vccd1 vccd1 net1109 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout396_X net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout133 _06336_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08011__B1 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11697__A1 _04987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09890__B net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout144 net147 vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12801__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout155 _05884_ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__buf_2
Xfanout166 _05288_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__clkbuf_2
Xfanout177 _05670_ vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_126_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout188 _05664_ vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_126_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout199 net200 vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__clkbuf_2
XFILLER_87_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout942_A _01717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout563_X net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07989_ net614 _02824_ net564 vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11417__S net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09728_ _04275_ _04299_ _04561_ _04538_ vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__or4b_2
XTAP_TAPCELL_ROW_2_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14297__Q datapath.rf.registers\[0\]\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08314__B2 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout730_X net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09659_ _03824_ _04493_ _04494_ _04492_ net632 vssd1 vssd1 vccd1 vccd1 _04495_ sky130_fd_sc_hd__o32a_1
XFILLER_16_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout828_X net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06594__X _01435_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12670_ _06498_ _06504_ _06503_ _06502_ vssd1 vssd1 vccd1 vccd1 _06506_ sky130_fd_sc_hd__o211ai_1
XFILLER_151_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10409__C1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11621_ _05794_ _05843_ vssd1 vssd1 vccd1 vccd1 _05845_ sky130_fd_sc_hd__nand2_1
XANTENNA__08078__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11152__S net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14340_ clknet_leaf_17_clk _01045_ net1109 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11552_ net1006 _05775_ vssd1 vssd1 vccd1 vccd1 _05776_ sky130_fd_sc_hd__nor2_4
XFILLER_156_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10503_ screen.counter.ct\[2\] _05331_ vssd1 vssd1 vccd1 vccd1 _05333_ sky130_fd_sc_hd__nand2_1
XANTENNA__10991__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11483_ net294 net1833 net510 vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__mux2_1
X_14271_ clknet_leaf_4_clk _00976_ net1077 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09027__C1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13222_ clknet_leaf_29_clk _00032_ net1133 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10434_ datapath.PC\[1\] net1240 _05242_ _05269_ vssd1 vssd1 vccd1 vccd1 _05270_
+ sky130_fd_sc_hd__o22a_2
Xwire589 _02691_ vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__buf_1
XANTENNA__08314__X _03150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06770__A _01571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13079__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07053__A1 datapath.rf.registers\[0\]\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10365_ _05146_ _05167_ _05177_ vssd1 vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__or3_1
X_13153_ net1886 net198 net384 vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__mux2_1
XANTENNA__08250__B1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12104_ screen.register.currentXbus\[31\] net996 net995 screen.register.currentXbus\[7\]
+ _06141_ vssd1 vssd1 vccd1 vccd1 _06142_ sky130_fd_sc_hd__a221o_1
X_13084_ net2202 net210 net386 vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__mux2_1
XFILLER_151_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10296_ net892 _05127_ _05131_ vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__o21a_1
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12035_ screen.register.currentYbus\[27\] _05757_ _06018_ screen.register.currentYbus\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06077_ sky130_fd_sc_hd__a22o_1
XFILLER_104_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07356__A2 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_69_Left_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11327__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06929__B net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13986_ clknet_leaf_108_clk _00763_ net1219 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_93_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07108__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12937_ net281 net1596 net397 vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__mux2_1
XFILLER_34_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12868_ net297 net2292 net399 vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__mux2_1
X_14607_ clknet_leaf_25_clk _01312_ net1137 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11819_ _01532_ net1017 net316 net336 datapath.ru.latched_instruction\[25\] vssd1
+ vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__a32o_1
XANTENNA__11062__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12799_ net1753 net288 net493 vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__mux2_1
XANTENNA__07816__B1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14538_ clknet_leaf_61_clk _01243_ net1164 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_78_Left_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14469_ clknet_leaf_141_clk _01174_ net1187 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_146_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06951__Y _01787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07010_ datapath.rf.registers\[17\]\[31\] net746 net722 datapath.rf.registers\[18\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_77_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07595__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08961_ _03795_ _03796_ net450 vssd1 vssd1 vccd1 vccd1 _03797_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11679__A1 _05199_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07912_ datapath.rf.registers\[8\]\[12\] net876 net832 datapath.rf.registers\[30\]\[12\]
+ _02747_ vssd1 vssd1 vccd1 vccd1 _02748_ sky130_fd_sc_hd__a221o_1
XFILLER_97_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_87_Left_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08892_ _03480_ _03727_ vssd1 vssd1 vccd1 vccd1 _03728_ sky130_fd_sc_hd__and2_1
XANTENNA__07347__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09741__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07843_ _02665_ _02666_ _02673_ _02678_ vssd1 vssd1 vccd1 vccd1 _02679_ sky130_fd_sc_hd__or4_1
XFILLER_68_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10351__A1 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07942__C net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11237__S net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07774_ _02607_ _02608_ _02609_ vssd1 vssd1 vccd1 vccd1 _02610_ sky130_fd_sc_hd__or3_1
X_09513_ _02704_ net554 net550 vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__or3_1
X_06725_ _01540_ _01563_ datapath.ru.n_memread datapath.ru.n_memwrite vssd1 vssd1
+ vccd1 vccd1 _01564_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_88_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06858__A1 datapath.ru.latched_instruction\[29\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06656_ mmio.memload_or_instruction\[20\] datapath.ru.latched_instruction\[20\] net1049
+ vssd1 vssd1 vccd1 vccd1 _01495_ sky130_fd_sc_hd__and3_1
X_09444_ _04278_ _04279_ vssd1 vssd1 vccd1 vccd1 _04280_ sky130_fd_sc_hd__nand2_1
XFILLER_80_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07303__X _02139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06587_ screen.screenEdge.enable3 vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__inv_2
X_09375_ _03574_ _04210_ net580 vssd1 vssd1 vccd1 vccd1 _04211_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout523_A _05723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_96_Left_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07807__B1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08326_ datapath.rf.registers\[9\]\[4\] net703 net660 datapath.rf.registers\[5\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03162_ sky130_fd_sc_hd__a22o_1
XFILLER_137_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08257_ datapath.rf.registers\[8\]\[5\] net877 _03090_ _03091_ _03092_ vssd1 vssd1
+ vccd1 vccd1 _03093_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout311_X net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08480__B1 _01768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout409_X net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07208_ _02036_ _02037_ _02042_ _02043_ vssd1 vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__nor4_1
XFILLER_137_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xteam_04_1320 vssd1 vssd1 vccd1 vccd1 team_04_1320/HI gpio_out[24] sky130_fd_sc_hd__conb_1
X_08188_ datapath.rf.registers\[19\]\[7\] net732 net689 datapath.rf.registers\[31\]\[7\]
+ _03023_ vssd1 vssd1 vccd1 vccd1 _03024_ sky130_fd_sc_hd__a221o_1
Xteam_04_1331 vssd1 vssd1 vccd1 vccd1 gpio_oeb[5] team_04_1331/LO sky130_fd_sc_hd__conb_1
XFILLER_146_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xteam_04_1342 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] team_04_1342/LO sky130_fd_sc_hd__conb_1
XANTENNA_fanout892_A net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07139_ datapath.rf.registers\[4\]\[28\] net864 net818 datapath.rf.registers\[7\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01975_ sky130_fd_sc_hd__a22o_1
XANTENNA__08232__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07586__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10150_ net224 _04985_ net1293 vssd1 vssd1 vccd1 vccd1 _04986_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout680_X net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout778_X net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11936__A _02090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10081_ _04899_ _04902_ vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07338__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11655__B _05874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout945_X net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire1045 _01534_ vssd1 vssd1 vccd1 vccd1 net1045 sky130_fd_sc_hd__buf_2
XANTENNA__11147__S net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13840_ clknet_leaf_141_clk _00649_ net1095 vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10893__A2 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13771_ clknet_leaf_82_clk _00580_ net1256 vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_148_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_148_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08299__B1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10986__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10983_ net1694 net253 net434 vssd1 vssd1 vccd1 vccd1 _00048_ sky130_fd_sc_hd__mux2_1
XFILLER_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12722_ columns.count\[8\] _06541_ vssd1 vssd1 vccd1 vccd1 _06544_ sky130_fd_sc_hd__or2_1
XFILLER_15_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_133_Right_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12653_ datapath.mulitply_result\[24\] datapath.multiplication_module.multiplicand_i\[24\]
+ vssd1 vssd1 vccd1 vccd1 _06491_ sky130_fd_sc_hd__nand2_1
XFILLER_130_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_139_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11604_ net999 net997 net995 _05827_ vssd1 vssd1 vccd1 vccd1 _05828_ sky130_fd_sc_hd__or4b_1
XANTENNA__12398__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09799__B1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12584_ _06432_ _06433_ vssd1 vssd1 vccd1 vccd1 _06434_ sky130_fd_sc_hd__xnor2_1
XFILLER_11_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14323_ clknet_leaf_34_clk _01028_ net1127 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11535_ _05293_ _05750_ vssd1 vssd1 vccd1 vccd1 _05759_ sky130_fd_sc_hd__nor2_1
XANTENNA__08471__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14254_ clknet_leaf_2_clk _00959_ net1062 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_137_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11466_ net2408 net210 net406 vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__mux2_1
X_13205_ clknet_leaf_19_clk _00015_ net1116 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08223__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10417_ _05250_ _05251_ _05252_ net351 vssd1 vssd1 vccd1 vccd1 _05253_ sky130_fd_sc_hd__a211o_1
X_14185_ clknet_leaf_47_clk _00940_ net1175 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11397_ net1927 net233 net410 vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__mux2_1
XFILLER_99_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08204__B net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07577__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13136_ net1674 net278 net385 vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__mux2_1
XFILLER_151_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10348_ net634 _05183_ _05179_ net227 vssd1 vssd1 vccd1 vccd1 _05184_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_55_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10279_ net222 _05114_ net1292 vssd1 vssd1 vccd1 vccd1 _05115_ sky130_fd_sc_hd__a21o_1
X_13067_ net1749 net294 net387 vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__mux2_1
XANTENNA__07329__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12018_ screen.register.currentYbus\[10\] _05776_ net999 screen.register.currentXbus\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06061_ sky130_fd_sc_hd__a22o_1
XANTENNA__11057__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09035__B _03867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_139_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_139_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13969_ clknet_leaf_106_clk _00747_ net1223 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07490_ _02315_ _02323_ _02324_ _02325_ vssd1 vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__or4_1
XFILLER_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09160_ _03994_ _03995_ vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__nand2_1
X_08111_ datapath.rf.registers\[30\]\[8\] net834 net812 datapath.rf.registers\[13\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02947_ sky130_fd_sc_hd__a22o_1
X_09091_ net552 net548 _02069_ vssd1 vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__a21o_1
XANTENNA__07777__Y _02613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10484__X _05314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08042_ net614 _02877_ vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__or2_1
XFILLER_116_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold901 mmio.memload_or_instruction\[31\] vssd1 vssd1 vccd1 vccd1 net2249 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold912 screen.controlBus\[3\] vssd1 vssd1 vccd1 vccd1 net2260 sky130_fd_sc_hd__dlygate4sd3_1
Xhold923 datapath.rf.registers\[17\]\[5\] vssd1 vssd1 vccd1 vccd1 net2271 sky130_fd_sc_hd__dlygate4sd3_1
Xhold934 mmio.memload_or_instruction\[29\] vssd1 vssd1 vccd1 vccd1 net2282 sky130_fd_sc_hd__dlygate4sd3_1
Xhold945 datapath.rf.registers\[8\]\[24\] vssd1 vssd1 vccd1 vccd1 net2293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold956 datapath.rf.registers\[13\]\[27\] vssd1 vssd1 vccd1 vccd1 net2304 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold967 datapath.rf.registers\[2\]\[31\] vssd1 vssd1 vccd1 vccd1 net2315 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold978 mmio.key_data\[4\] vssd1 vssd1 vccd1 vccd1 net2326 sky130_fd_sc_hd__dlygate4sd3_1
Xhold989 datapath.rf.registers\[25\]\[29\] vssd1 vssd1 vccd1 vccd1 net2337 sky130_fd_sc_hd__dlygate4sd3_1
X_09993_ _04719_ _04828_ vssd1 vssd1 vccd1 vccd1 _04829_ sky130_fd_sc_hd__xor2_1
XFILLER_135_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08944_ _02169_ _02217_ net445 vssd1 vssd1 vccd1 vccd1 _03780_ sky130_fd_sc_hd__mux2_1
XANTENNA__07953__B net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08875_ _03205_ _03263_ net446 vssd1 vssd1 vccd1 vccd1 _03711_ sky130_fd_sc_hd__mux2_1
XFILLER_151_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07826_ datapath.rf.registers\[3\]\[14\] net771 net692 datapath.rf.registers\[13\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__a22o_1
XFILLER_57_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07740__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07757_ datapath.rf.registers\[11\]\[15\] net983 net939 vssd1 vssd1 vccd1 vccd1 _02593_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout261_X net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout738_A net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10088__B1 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06708_ datapath.ru.latched_instruction\[12\] datapath.ru.latched_instruction\[13\]
+ datapath.ru.latched_instruction\[14\] datapath.ru.latched_instruction\[15\] vssd1
+ vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__or4_1
XANTENNA__11824__B2 datapath.ru.latched_instruction\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_13_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07688_ datapath.rf.registers\[25\]\[17\] net728 net720 datapath.rf.registers\[20\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__a22o_1
XANTENNA__09493__A2 _04328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09427_ net331 _04256_ _04262_ _03613_ vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__o211a_1
X_06639_ net1288 net1283 datapath.ru.latched_instruction\[31\] mmio.memload_or_instruction\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_23_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout526_X net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07968__X _02804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09358_ net648 _04193_ net438 vssd1 vssd1 vccd1 vccd1 _04194_ sky130_fd_sc_hd__a21o_1
X_08309_ datapath.rf.registers\[20\]\[4\] net839 net819 datapath.rf.registers\[5\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__a22o_1
XANTENNA__07687__Y _02523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08453__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09289_ net365 _04124_ _04123_ vssd1 vssd1 vccd1 vccd1 _04125_ sky130_fd_sc_hd__o21a_1
XANTENNA__11430__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11320_ net1980 net268 net416 vssd1 vssd1 vccd1 vccd1 _00365_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11251_ net270 net2120 net420 vssd1 vssd1 vccd1 vccd1 _00300_ sky130_fd_sc_hd__mux2_1
XFILLER_134_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10202_ _03978_ _04604_ net895 vssd1 vssd1 vccd1 vccd1 _05038_ sky130_fd_sc_hd__a21o_1
XFILLER_140_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11182_ net280 net2130 net425 vssd1 vssd1 vccd1 vccd1 _00234_ sky130_fd_sc_hd__mux2_1
XFILLER_134_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14036__RESET_B net1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10133_ net1265 _03746_ vssd1 vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__xnor2_1
XFILLER_121_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12304__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input34_A en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10064_ datapath.PC\[30\] net596 vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__xnor2_2
XFILLER_85_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07192__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07731__A2 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13823_ clknet_leaf_112_clk _00632_ net1197 vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__dfrtp_1
XFILLER_47_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13092__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11815__A1 datapath.ru.latched_instruction\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13754_ clknet_leaf_88_clk _00563_ net1253 vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__dfrtp_1
XFILLER_141_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11815__B2 _01505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10966_ _01502_ net655 _05701_ _05702_ vssd1 vssd1 vccd1 vccd1 _05703_ sky130_fd_sc_hd__o22a_1
XANTENNA__09484__A2 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12705_ net1559 _06532_ vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__xnor2_1
XFILLER_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13685_ clknet_leaf_94_clk _00495_ net1211 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10897_ net898 _05642_ net616 vssd1 vssd1 vccd1 vccd1 _05643_ sky130_fd_sc_hd__o21a_1
XFILLER_148_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12636_ datapath.mulitply_result\[21\] datapath.multiplication_module.multiplicand_i\[21\]
+ vssd1 vssd1 vccd1 vccd1 _06477_ sky130_fd_sc_hd__and2_1
XFILLER_34_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12567_ net501 _06418_ _06419_ net505 net2075 vssd1 vssd1 vccd1 vccd1 _00919_ sky130_fd_sc_hd__a32o_1
XANTENNA__11340__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14306_ clknet_leaf_1_clk _01011_ net1056 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11518_ screen.counter.ct\[2\] _01425_ net1001 net1276 vssd1 vssd1 vccd1 vccd1 _05743_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__07757__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12498_ net232 net2436 net507 vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__mux2_1
Xhold208 datapath.multiplication_module.multiplicand_i\[5\] vssd1 vssd1 vccd1 vccd1
+ net1556 sky130_fd_sc_hd__dlygate4sd3_1
Xhold219 datapath.rf.registers\[4\]\[3\] vssd1 vssd1 vccd1 vccd1 net1567 sky130_fd_sc_hd__dlygate4sd3_1
X_14237_ clknet_leaf_122_clk datapath.multiplication_module.multiplier_i_n\[5\] net1214
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i\[5\] sky130_fd_sc_hd__dfrtp_1
X_11449_ datapath.rf.registers\[14\]\[5\] net296 net407 vssd1 vssd1 vccd1 vccd1 _00487_
+ sky130_fd_sc_hd__mux2_1
X_14168_ clknet_leaf_70_clk _00923_ net1244 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_125_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13119_ net200 net2248 net470 vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__mux2_1
XFILLER_86_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14099_ clknet_leaf_122_clk _00865_ net1201 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_06990_ net966 _01825_ vssd1 vssd1 vccd1 vccd1 _01826_ sky130_fd_sc_hd__and2_1
XANTENNA__07118__X _01954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07970__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1270 screen.counter.ct\[17\] vssd1 vssd1 vccd1 vccd1 net1270 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09172__A1 _03800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13759__RESET_B net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1281 net1285 vssd1 vssd1 vccd1 vccd1 net1281 sky130_fd_sc_hd__buf_2
X_08660_ _02169_ _02190_ vssd1 vssd1 vccd1 vccd1 _03496_ sky130_fd_sc_hd__or2_1
Xfanout1292 _01436_ vssd1 vssd1 vccd1 vccd1 net1292 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08885__A _01611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07722__A2 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07611_ datapath.rf.registers\[10\]\[18\] net879 net845 datapath.rf.registers\[1\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__a22o_1
XFILLER_26_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08591_ _03230_ _03423_ _03231_ _03127_ _03174_ vssd1 vssd1 vccd1 vccd1 _03427_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_85_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07542_ datapath.rf.registers\[9\]\[20\] net702 net671 datapath.rf.registers\[7\]\[20\]
+ _02377_ vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_101_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07473_ datapath.rf.registers\[25\]\[21\] net841 net804 datapath.rf.registers\[28\]\[21\]
+ _02308_ vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__a221o_1
XFILLER_62_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09212_ _03898_ _03904_ net342 vssd1 vssd1 vccd1 vccd1 _04048_ sky130_fd_sc_hd__mux2_1
XFILLER_50_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09143_ _03459_ _03502_ vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12346__S net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07948__B net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout221_A _05610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11250__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09074_ _03493_ net628 _03721_ _03494_ net645 vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__a221o_1
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07667__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08125__A _02960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06997__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11990__B1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08025_ datapath.rf.registers\[26\]\[10\] net780 net677 datapath.rf.registers\[29\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__a22o_1
XFILLER_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold720 datapath.rf.registers\[20\]\[2\] vssd1 vssd1 vccd1 vccd1 net2068 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1130_A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold731 datapath.rf.registers\[22\]\[16\] vssd1 vssd1 vccd1 vccd1 net2079 sky130_fd_sc_hd__dlygate4sd3_1
Xhold742 datapath.rf.registers\[12\]\[1\] vssd1 vssd1 vccd1 vccd1 net2090 sky130_fd_sc_hd__dlygate4sd3_1
Xhold753 datapath.rf.registers\[23\]\[21\] vssd1 vssd1 vccd1 vccd1 net2101 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold764 datapath.rf.registers\[30\]\[24\] vssd1 vssd1 vccd1 vccd1 net2112 sky130_fd_sc_hd__dlygate4sd3_1
Xhold775 screen.register.currentYbus\[0\] vssd1 vssd1 vccd1 vccd1 net2123 sky130_fd_sc_hd__dlygate4sd3_1
Xhold786 datapath.rf.registers\[0\]\[14\] vssd1 vssd1 vccd1 vccd1 net2134 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout688_A net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11742__B1 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08779__B net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold797 datapath.rf.registers\[3\]\[17\] vssd1 vssd1 vccd1 vccd1 net2145 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09976_ _04733_ _04735_ _04810_ _04732_ vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__a31o_1
XANTENNA__08498__C _01825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07961__A2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08927_ net566 _03761_ _03762_ vssd1 vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__a21oi_1
XFILLER_29_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout476_X net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08858_ net566 _01889_ net445 vssd1 vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__mux2_1
XANTENNA__07174__B1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07809_ datapath.rf.registers\[15\]\[14\] net800 net792 datapath.rf.registers\[18\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02645_ sky130_fd_sc_hd__a22o_1
XANTENNA__11933__B net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06921__B1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08789_ _03296_ net576 _03624_ vssd1 vssd1 vccd1 vccd1 _03625_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout643_X net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11425__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10820_ net1266 _05565_ datapath.PC\[13\] vssd1 vssd1 vccd1 vccd1 _05577_ sky130_fd_sc_hd__a21oi_1
XFILLER_26_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout810_X net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10751_ _01640_ _05516_ vssd1 vssd1 vccd1 vccd1 _05518_ sky130_fd_sc_hd__or2_2
XFILLER_71_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13470_ clknet_leaf_148_clk _00280_ net1061 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10682_ net1013 _05444_ _05464_ _05489_ _01430_ vssd1 vssd1 vccd1 vccd1 _05500_ sky130_fd_sc_hd__o41a_1
XFILLER_139_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12421_ _05978_ net156 vssd1 vssd1 vccd1 vccd1 _06358_ sky130_fd_sc_hd__nor2_1
XANTENNA__08426__B1 _03261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11160__S net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12352_ net229 _05661_ net638 vssd1 vssd1 vccd1 vccd1 _06318_ sky130_fd_sc_hd__a21o_1
XANTENNA__10784__A1 _01438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11303_ net184 net2337 net523 vssd1 vssd1 vccd1 vccd1 _00351_ sky130_fd_sc_hd__mux2_1
XANTENNA__10852__X _05605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12283_ net891 _04515_ vssd1 vssd1 vccd1 vccd1 _06268_ sky130_fd_sc_hd__nor2_1
X_14022_ clknet_leaf_77_clk _00791_ net1249 vssd1 vssd1 vccd1 vccd1 datapath.PC\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12525__A2 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11234_ net194 net1866 net526 vssd1 vssd1 vccd1 vccd1 _00284_ sky130_fd_sc_hd__mux2_1
XFILLER_4_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13087__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11165_ net201 net1837 net531 vssd1 vssd1 vccd1 vccd1 _00218_ sky130_fd_sc_hd__mux2_1
XFILLER_96_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10116_ _04873_ _04951_ vssd1 vssd1 vccd1 vccd1 _04952_ sky130_fd_sc_hd__nand2_1
XANTENNA__12289__A1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11096_ net203 net2124 net535 vssd1 vssd1 vccd1 vccd1 _00153_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_147_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08201__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10047_ datapath.PC\[24\] net594 _04821_ vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__a21o_1
XANTENNA__13852__RESET_B net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_42_Left_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold80 net84 vssd1 vssd1 vccd1 vccd1 net1428 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold91 net52 vssd1 vssd1 vccd1 vccd1 net1439 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_63_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11335__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06937__B net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13806_ clknet_leaf_73_clk _00615_ net1242 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11998_ _06041_ vssd1 vssd1 vccd1 vccd1 _06042_ sky130_fd_sc_hd__inv_2
XFILLER_90_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13737_ clknet_leaf_77_clk _00547_ net1246 vssd1 vssd1 vccd1 vccd1 datapath.i_ack
+ sky130_fd_sc_hd__dfrtp_1
X_10949_ _05687_ _05686_ net653 _01477_ vssd1 vssd1 vccd1 vccd1 _05688_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_32_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_70_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_31_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13668_ clknet_leaf_21_clk _00478_ net1163 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06953__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12619_ _06456_ _06458_ vssd1 vssd1 vccd1 vccd1 _06463_ sky130_fd_sc_hd__nor2_1
XANTENNA__08417__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13599_ clknet_leaf_13_clk _00409_ net1079 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10775__A1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09983__B net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09830_ _01610_ net904 vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__nor2_1
Xfanout507 net508 vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__clkbuf_8
Xfanout518 net519 vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_111_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout529 _05721_ vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__clkbuf_4
XFILLER_99_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06746__A3 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09761_ net317 _04365_ _04592_ _04595_ _04596_ vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__o2111a_1
X_06973_ _01636_ _01647_ vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__nor2_2
X_08712_ net559 _03358_ vssd1 vssd1 vccd1 vccd1 _03548_ sky130_fd_sc_hd__xnor2_2
X_09692_ net379 _03879_ _04527_ _03614_ vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__a211o_1
XFILLER_132_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07156__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_722 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08643_ _03477_ _03478_ vssd1 vssd1 vccd1 vccd1 _03479_ sky130_fd_sc_hd__and2_1
XANTENNA__07950__C net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout171_A _05688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11245__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout269_A _05570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08574_ datapath.rf.registers\[2\]\[0\] net914 net910 vssd1 vssd1 vccd1 vccd1 _03410_
+ sky130_fd_sc_hd__and3_1
XFILLER_81_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07024__A _01859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07525_ datapath.rf.registers\[8\]\[20\] net876 _02335_ _02336_ _02345_ vssd1 vssd1
+ vccd1 vccd1 _02361_ sky130_fd_sc_hd__a2111o_1
XFILLER_35_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1080_A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_61_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout436_A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1178_A net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07959__A net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07456_ datapath.rf.registers\[7\]\[21\] _01717_ net933 vssd1 vssd1 vccd1 vccd1 _02292_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_33_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout224_X net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07387_ _02219_ _02220_ _02221_ _02222_ vssd1 vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__or4_1
XFILLER_6_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09126_ net551 net547 _02217_ vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_98_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09057_ _03681_ _03687_ net449 vssd1 vssd1 vccd1 vccd1 _03893_ sky130_fd_sc_hd__mux2_1
XANTENNA__12804__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08008_ datapath.rf.registers\[1\]\[10\] net847 _02829_ _02832_ _02841_ vssd1 vssd1
+ vccd1 vccd1 _02844_ sky130_fd_sc_hd__a2111o_1
Xhold550 datapath.rf.registers\[23\]\[29\] vssd1 vssd1 vccd1 vccd1 net1898 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10518__A1 _05335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold561 datapath.rf.registers\[16\]\[2\] vssd1 vssd1 vccd1 vccd1 net1909 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold572 datapath.rf.registers\[27\]\[8\] vssd1 vssd1 vccd1 vccd1 net1920 sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 datapath.rf.registers\[11\]\[15\] vssd1 vssd1 vccd1 vccd1 net1931 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08187__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold594 datapath.rf.registers\[9\]\[8\] vssd1 vssd1 vccd1 vccd1 net1942 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07395__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout760_X net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09959_ datapath.PC\[8\] _02981_ vssd1 vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout858_X net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12970_ net280 net2052 net481 vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__mux2_1
XANTENNA__07147__B1 _01824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1250 screen.controlBus\[0\] vssd1 vssd1 vccd1 vccd1 net2598 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1261 datapath.rf.registers\[30\]\[2\] vssd1 vssd1 vccd1 vccd1 net2609 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11663__B _05874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11921_ _02331_ net656 vssd1 vssd1 vccd1 vccd1 _05978_ sky130_fd_sc_hd__nand2_1
Xhold1272 datapath.rf.registers\[26\]\[19\] vssd1 vssd1 vccd1 vccd1 net2620 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1283 datapath.rf.registers\[26\]\[1\] vssd1 vssd1 vccd1 vccd1 net2631 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11155__S net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1294 datapath.multiplication_module.multiplicand_i\[12\] vssd1 vssd1 vccd1 vccd1
+ net2642 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_61_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14640_ clknet_leaf_25_clk _01345_ net1158 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[28\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_142_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ screen.csx _05930_ _05926_ vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__mux2_1
XFILLER_73_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ datapath.mulitply_result\[10\] net598 net620 vssd1 vssd1 vccd1 vccd1 _05563_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__10994__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14571_ clknet_leaf_57_clk _01276_ net1160 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11783_ keypad.apps.app_c\[1\] _05896_ vssd1 vssd1 vccd1 vccd1 _05897_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_52_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08111__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13522_ clknet_leaf_30_clk _00332_ net1124 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10734_ net1561 net568 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[20\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__07855__D1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06673__A2 _01466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13453_ clknet_leaf_125_clk _00263_ net1205 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10665_ _05443_ _05465_ _05483_ vssd1 vssd1 vccd1 vccd1 _05484_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_11_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12404_ net1406 net130 _06349_ vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__a21o_1
X_13384_ clknet_leaf_64_clk _00194_ net1236 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[26\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10596_ screen.register.currentYbus\[5\] screen.register.currentYbus\[4\] screen.register.currentYbus\[7\]
+ screen.register.currentYbus\[6\] vssd1 vssd1 vccd1 vccd1 _05417_ sky130_fd_sc_hd__or4_1
XFILLER_5_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12335_ net1265 net310 _06305_ _04972_ vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__a22o_1
XANTENNA__07083__C1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12266_ datapath.PC\[3\] net308 _06250_ _06255_ vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__a22o_1
X_14005_ clknet_leaf_111_clk screen.counter.ack net1198 vssd1 vssd1 vccd1 vccd1 screen.counter.ack1
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08178__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11217_ net277 net1838 net528 vssd1 vssd1 vccd1 vccd1 _00267_ sky130_fd_sc_hd__mux2_1
XFILLER_96_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 ADR_O[8] sky130_fd_sc_hd__buf_2
X_12197_ screen.counter.currentCt\[1\] screen.counter.currentCt\[2\] _06205_ vssd1
+ vssd1 vccd1 vccd1 _06209_ sky130_fd_sc_hd__and3_1
XANTENNA__07386__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 DAT_O[17] sky130_fd_sc_hd__buf_2
XANTENNA__07925__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput92 net92 vssd1 vssd1 vccd1 vccd1 DAT_O[27] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_50_Left_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11148_ net283 net2176 net532 vssd1 vssd1 vccd1 vccd1 _00201_ sky130_fd_sc_hd__mux2_1
X_11079_ net291 net1989 net535 vssd1 vssd1 vccd1 vccd1 _00136_ sky130_fd_sc_hd__mux2_1
XFILLER_37_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07138__B1 _01760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11065__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_43_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_32_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07310_ net613 _02145_ net565 vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__a21oi_2
XFILLER_20_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08290_ _03125_ vssd1 vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__inv_2
XANTENNA__07310__B1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_9_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07241_ datapath.rf.registers\[14\]\[26\] net774 net726 datapath.rf.registers\[25\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02077_ sky130_fd_sc_hd__a22o_1
XANTENNA__07498__B net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07172_ datapath.rf.registers\[13\]\[27\] net811 net805 datapath.rf.registers\[28\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__a22o_1
XANTENNA__08106__C _01712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wire561_X net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07945__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10652__B _01435_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08169__A2 _01716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout304 net305 vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__clkbuf_2
Xfanout315 net316 vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__buf_2
XANTENNA__07377__B1 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout326 _03663_ vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__buf_2
XANTENNA__07019__A _01854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07916__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout337 net339 vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__buf_2
X_09813_ _03598_ _04648_ net579 vssd1 vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__o21ai_1
Xfanout348 _03662_ vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout359 net361 vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__buf_2
XANTENNA_fanout386_A net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09744_ net631 _04565_ _04567_ _04579_ vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__a22o_2
X_06956_ net991 net972 vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__nor2_1
XANTENNA__07129__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09675_ net906 _03565_ _04509_ _04510_ vssd1 vssd1 vccd1 vccd1 _04511_ sky130_fd_sc_hd__a211o_1
X_06887_ _01707_ net956 vssd1 vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__and2_4
XANTENNA_fanout1295_A _01436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08626_ _02241_ _03460_ _02242_ _02147_ _02191_ vssd1 vssd1 vccd1 vccd1 _03462_ sky130_fd_sc_hd__a2111o_1
XFILLER_70_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_124_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout720_A net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08557_ datapath.rf.registers\[16\]\[0\] net913 _01805_ vssd1 vssd1 vccd1 vccd1 _03393_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout818_A _01758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout439_X net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_34_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_51_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07508_ datapath.rf.registers\[23\]\[20\] net940 net922 vssd1 vssd1 vccd1 vccd1 _02344_
+ sky130_fd_sc_hd__and3_1
X_08488_ net614 _03322_ _03323_ vssd1 vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__or3_2
XANTENNA__07301__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07439_ datapath.rf.registers\[14\]\[22\] net774 net754 datapath.rf.registers\[12\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1250_X net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout606_X net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10450_ _05074_ _05285_ vssd1 vssd1 vccd1 vccd1 WEN sky130_fd_sc_hd__nor2_1
XFILLER_6_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06880__X _01716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09109_ net317 _03943_ net905 _03497_ vssd1 vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__11939__A _02045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07604__A1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10381_ _03547_ net626 _04172_ _03673_ _05216_ vssd1 vssd1 vccd1 vccd1 _05217_ sky130_fd_sc_hd__a221o_1
XFILLER_151_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12120_ screen.counter.ct\[11\] net1275 net1273 _06156_ vssd1 vssd1 vccd1 vccd1 _06157_
+ sky130_fd_sc_hd__and4_1
XANTENNA__09409__A _02660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_107_Left_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07080__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout975_X net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12051_ screen.register.currentXbus\[4\] net1000 _06018_ screen.register.currentYbus\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06092_ sky130_fd_sc_hd__a22o_1
Xhold380 datapath.rf.registers\[21\]\[20\] vssd1 vssd1 vccd1 vccd1 net1728 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold391 datapath.rf.registers\[30\]\[13\] vssd1 vssd1 vccd1 vccd1 net1739 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07368__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12361__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07907__A2 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11002_ _05689_ _05707_ vssd1 vssd1 vccd1 vccd1 _05708_ sky130_fd_sc_hd__nor2_1
XFILLER_78_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10989__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10372__C1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout860 net863 vssd1 vssd1 vccd1 vccd1 net860 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_144_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout871 _01724_ vssd1 vssd1 vccd1 vccd1 net871 sky130_fd_sc_hd__clkbuf_8
Xfanout882 net883 vssd1 vssd1 vccd1 vccd1 net882 sky130_fd_sc_hd__clkbuf_8
Xfanout893 net896 vssd1 vssd1 vccd1 vccd1 net893 sky130_fd_sc_hd__clkbuf_2
XFILLER_93_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08868__A0 _02805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12953_ net200 net2220 net395 vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__mux2_1
Xhold1080 datapath.rf.registers\[8\]\[15\] vssd1 vssd1 vccd1 vccd1 net2428 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1091 datapath.rf.registers\[19\]\[14\] vssd1 vssd1 vccd1 vccd1 net2439 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08332__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11904_ net134 _05966_ _05965_ vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_47_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_116_Left_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12884_ net216 net1597 net398 vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__mux2_1
XANTENNA__09154__A_N net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14623_ clknet_leaf_13_clk _01328_ net1077 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_11835_ net1277 screen.counter.ct\[11\] screen.counter.ct\[19\] net1276 vssd1 vssd1
+ vccd1 vccd1 _05914_ sky130_fd_sc_hd__or4b_1
XFILLER_26_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_25_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__10427__B1 _03667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14554_ clknet_leaf_2_clk _01259_ net1064 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_11766_ net1508 net143 net138 _02090_ vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__a22o_1
XANTENNA__08194__S net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13505_ clknet_leaf_46_clk _00315_ net1172 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10717_ net1851 net572 vssd1 vssd1 vccd1 vccd1 _05511_ sky130_fd_sc_hd__nor2_1
X_14485_ clknet_leaf_130_clk _01190_ net1111 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11697_ _04987_ net153 net148 net1418 vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__a22o_1
XFILLER_146_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13436_ clknet_leaf_7_clk _00246_ net1073 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10648_ _05437_ _05439_ _05440_ vssd1 vssd1 vccd1 vccd1 _05468_ sky130_fd_sc_hd__or3_1
XANTENNA__06790__X _01626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13367_ clknet_leaf_126_clk _00177_ net1205 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_125_Left_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10579_ _02217_ net563 _02311_ _02364_ vssd1 vssd1 vccd1 vccd1 _05402_ sky130_fd_sc_hd__or4_1
XANTENNA__10753__A net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06950__B net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12318_ datapath.PC\[17\] net307 _06293_ _05024_ vssd1 vssd1 vccd1 vccd1 _00796_
+ sky130_fd_sc_hd__o22a_1
XFILLER_5_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13298_ clknet_leaf_32_clk _00108_ net1123 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_75_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12249_ screen.counter.currentCt\[21\] screen.counter.currentCt\[20\] _06238_ vssd1
+ vssd1 vccd1 vccd1 _06242_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_75_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08020__A1 datapath.rf.registers\[0\]\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08571__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06810_ net1004 net1020 _01645_ net1028 datapath.ru.latched_instruction\[23\] vssd1
+ vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__a32oi_4
X_07790_ datapath.rf.registers\[22\]\[15\] net735 net668 datapath.rf.registers\[21\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02626_ sky130_fd_sc_hd__a22o_1
XANTENNA__12104__B1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_147_Right_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09054__A net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_134_Left_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06741_ _01579_ vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__inv_2
XANTENNA__08323__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09460_ net324 _03859_ _04294_ _04295_ net642 vssd1 vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__o2111a_1
X_06672_ net1287 net1282 mmio.memload_or_instruction\[15\] vssd1 vssd1 vccd1 vccd1
+ _01511_ sky130_fd_sc_hd__or3b_1
XFILLER_52_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07531__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08411_ datapath.rf.registers\[13\]\[2\] net988 net918 vssd1 vssd1 vccd1 vccd1 _03247_
+ sky130_fd_sc_hd__and3_1
X_09391_ net362 _04063_ _04226_ vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_16_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_51_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08342_ datapath.rf.registers\[15\]\[3\] net989 net916 vssd1 vssd1 vccd1 vccd1 _03178_
+ sky130_fd_sc_hd__and3_1
XFILLER_32_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08273_ datapath.rf.registers\[4\]\[5\] net715 net665 datapath.rf.registers\[15\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03109_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout134_A net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07224_ datapath.rf.registers\[22\]\[26\] net821 net818 datapath.rf.registers\[7\]\[26\]
+ _02059_ vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__a221o_1
XANTENNA__07021__B net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07155_ datapath.rf.registers\[19\]\[28\] net733 net690 datapath.rf.registers\[31\]\[28\]
+ _01990_ vssd1 vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__a221o_1
XANTENNA__13955__RESET_B net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout301_A _05529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1043_A net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12591__B1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07086_ datapath.rf.registers\[14\]\[29\] net831 net796 datapath.rf.registers\[29\]\[29\]
+ _01921_ vssd1 vssd1 vccd1 vccd1 _01922_ sky130_fd_sc_hd__a221o_1
XANTENNA__07062__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1210_A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout134 net135 vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__buf_2
Xfanout145 net147 vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__buf_2
XANTENNA_fanout670_A _01832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout156 net157 vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__buf_2
XFILLER_86_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout167 _05288_ vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__buf_1
XANTENNA_fanout768_A net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout389_X net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout178 _05670_ vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_126_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07988_ datapath.rf.registers\[0\]\[11\] net783 _02820_ _02823_ vssd1 vssd1 vccd1
+ vccd1 _02824_ sky130_fd_sc_hd__o22a_4
XTAP_TAPCELL_ROW_126_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_114_Right_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09727_ _04538_ _04562_ vssd1 vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__nand2_1
XFILLER_101_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06939_ net976 net915 vssd1 vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__and2_1
XFILLER_28_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout556_X net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout935_A net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09511__A1 _03263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09658_ _03429_ _03563_ vssd1 vssd1 vccd1 vccd1 _04494_ sky130_fd_sc_hd__nor2_1
X_08609_ _03440_ _03443_ vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout723_X net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09589_ _04424_ _04403_ net648 _04411_ vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__and4b_1
XANTENNA__11433__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11620_ _05836_ _05843_ vssd1 vssd1 vccd1 vccd1 _05844_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_42_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11551_ _05749_ _05774_ vssd1 vssd1 vccd1 vccd1 _05775_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_42_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10502_ _05324_ _05330_ vssd1 vssd1 vccd1 vccd1 _05332_ sky130_fd_sc_hd__or2_1
X_14270_ clknet_leaf_150_clk _00975_ net1059 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11482_ net299 net2366 net511 vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_137_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13221_ clknet_leaf_114_clk _00031_ net1189 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10433_ net227 _05268_ net1292 vssd1 vssd1 vccd1 vccd1 _05269_ sky130_fd_sc_hd__a21o_1
XANTENNA__06770__B _01579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07589__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13152_ net2367 net200 net382 vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__mux2_1
X_10364_ _05106_ _05116_ _05188_ _05199_ vssd1 vssd1 vccd1 vccd1 _05200_ sky130_fd_sc_hd__or4_1
XFILLER_3_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12103_ screen.register.currentYbus\[23\] _05773_ net999 screen.register.currentXbus\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06141_ sky130_fd_sc_hd__a22o_1
XFILLER_124_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13083_ net1586 net216 net386 vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__mux2_1
X_10295_ net1038 _05128_ _05130_ net639 vssd1 vssd1 vccd1 vccd1 _05131_ sky130_fd_sc_hd__a211o_1
XANTENNA__12334__B1 _06253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12034_ _05840_ _06058_ vssd1 vssd1 vccd1 vccd1 _06076_ sky130_fd_sc_hd__or2_1
XANTENNA__13095__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07761__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout690 _01826_ vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__clkbuf_4
X_13985_ clknet_leaf_108_clk _00762_ net1221 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08305__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12936_ net285 net1995 net396 vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__mux2_1
X_12867_ net300 net2645 net398 vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__mux2_1
XFILLER_34_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11343__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11818_ datapath.ru.latched_instruction\[24\] net334 net314 _01463_ vssd1 vssd1 vccd1
+ vccd1 _00684_ sky130_fd_sc_hd__a22o_1
X_14606_ clknet_leaf_5_clk _01311_ net1067 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12798_ net2105 net260 net493 vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__mux2_1
XFILLER_30_931 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14537_ clknet_leaf_62_clk _01242_ net1234 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11749_ net1445 net147 net142 _02934_ vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__a22o_1
XFILLER_41_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07292__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14468_ clknet_leaf_21_clk _01173_ net1163 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06961__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13419_ clknet_leaf_56_clk _00229_ net1173 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_14399_ clknet_leaf_12_clk _01104_ net1082 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12573__B1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07044__A2 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08960_ _02660_ _02704_ net447 vssd1 vssd1 vccd1 vccd1 _03796_ sky130_fd_sc_hd__mux2_1
XANTENNA__13273__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12902__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_5_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_90_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07911_ datapath.rf.registers\[12\]\[12\] net826 net803 datapath.rf.registers\[3\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__a22o_1
XANTENNA__08240__X _03076_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08891_ _03599_ net579 _03606_ _03726_ vssd1 vssd1 vccd1 vccd1 _03727_ sky130_fd_sc_hd__a31o_1
XANTENNA__08544__A2 _01753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07842_ datapath.rf.registers\[30\]\[14\] net759 net661 datapath.rf.registers\[5\]\[14\]
+ _02677_ vssd1 vssd1 vccd1 vccd1 _02678_ sky130_fd_sc_hd__a221o_1
XFILLER_69_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07752__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08400__B net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07773_ datapath.rf.registers\[8\]\[15\] net877 net793 datapath.rf.registers\[31\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02609_ sky130_fd_sc_hd__a22o_1
XFILLER_65_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09512_ net458 _04345_ _04347_ net351 vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__a211oi_1
X_06724_ _01410_ _01546_ _01550_ net1015 vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__a31o_1
XFILLER_140_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09443_ net552 net548 _02804_ vssd1 vssd1 vccd1 vccd1 _04279_ sky130_fd_sc_hd__a21o_1
XFILLER_92_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06655_ mmio.memload_or_instruction\[20\] net1049 datapath.ru.latched_instruction\[20\]
+ vssd1 vssd1 vccd1 vccd1 _01494_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11253__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09374_ _03525_ _03573_ _03524_ vssd1 vssd1 vccd1 vccd1 _04210_ sky130_fd_sc_hd__a21oi_1
X_06586_ button\[3\] vssd1 vssd1 vccd1 vccd1 _01427_ sky130_fd_sc_hd__inv_2
X_08325_ datapath.rf.registers\[24\]\[4\] net766 _03159_ _03160_ vssd1 vssd1 vccd1
+ vccd1 _03161_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout1160_A net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout516_A _05731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1258_A net1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08256_ datapath.rf.registers\[20\]\[5\] net839 net800 datapath.rf.registers\[15\]\[5\]
+ net873 vssd1 vssd1 vccd1 vccd1 _03092_ sky130_fd_sc_hd__a221o_1
XANTENNA__06871__A _01630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07207_ _02030_ _02031_ _02033_ vssd1 vssd1 vccd1 vccd1 _02043_ sky130_fd_sc_hd__or3_1
Xteam_04_1310 vssd1 vssd1 vccd1 vccd1 team_04_1310/HI gpio_oeb[19] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_119_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xteam_04_1321 vssd1 vssd1 vccd1 vccd1 team_04_1321/HI gpio_out[25] sky130_fd_sc_hd__conb_1
X_08187_ datapath.rf.registers\[23\]\[7\] net700 _03022_ net788 vssd1 vssd1 vccd1
+ vccd1 _03023_ sky130_fd_sc_hd__a211o_1
XANTENNA_clkbuf_leaf_81_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xteam_04_1332 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] team_04_1332/LO sky130_fd_sc_hd__conb_1
XFILLER_152_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xteam_04_1343 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] team_04_1343/LO sky130_fd_sc_hd__conb_1
X_07138_ datapath.rf.registers\[6\]\[28\] net825 _01760_ datapath.rf.registers\[23\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout885_A net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12812__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07069_ _01895_ _01901_ _01903_ _01904_ vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__or4_1
XFILLER_133_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1213_X net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09393__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11936__B net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_96_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10080_ _04714_ _04910_ _04915_ net224 vssd1 vssd1 vccd1 vccd1 _04916_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout673_X net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11428__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09193__C1 _02311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08535__A2 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07743__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout840_X net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout938_X net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13770_ clknet_leaf_82_clk _00579_ net1256 vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12095__A2 _05778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10982_ net1712 net257 net435 vssd1 vssd1 vccd1 vccd1 _00047_ sky130_fd_sc_hd__mux2_1
X_12721_ _05894_ _06543_ vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__nor2_1
XFILLER_15_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11163__S net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12652_ net498 _06489_ _06490_ net502 net2592 vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_26_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_34_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11603_ screen.counter.ct\[0\] _05293_ _05302_ _05795_ vssd1 vssd1 vccd1 vccd1 _05827_
+ sky130_fd_sc_hd__o31a_1
X_12583_ _06425_ _06427_ _06426_ vssd1 vssd1 vccd1 vccd1 _06433_ sky130_fd_sc_hd__o21bai_2
XFILLER_156_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14322_ clknet_leaf_33_clk _01027_ net1126 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11534_ _05750_ _05754_ vssd1 vssd1 vccd1 vccd1 _05758_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_152_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14253_ clknet_leaf_132_clk _00958_ net1113 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_49_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11465_ net1542 net217 net406 vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__mux2_1
XFILLER_139_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13204_ clknet_leaf_20_clk _00014_ net1118 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12555__B1 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10416_ net463 net452 _04304_ net457 vssd1 vssd1 vccd1 vccd1 _05252_ sky130_fd_sc_hd__o211a_1
X_14184_ clknet_leaf_51_clk _00939_ net1182 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11396_ net2243 net237 net412 vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__mux2_1
XANTENNA__08204__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13135_ net1723 net282 net384 vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__mux2_1
XANTENNA__08774__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10347_ net1039 _05180_ _05182_ vssd1 vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_55_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07982__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13066_ net1932 net299 net387 vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__mux2_1
X_10278_ _04851_ _05113_ vssd1 vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__nand2_1
XANTENNA__11338__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12017_ screen.register.currentYbus\[26\] _05786_ net995 screen.register.currentXbus\[2\]
+ _05779_ vssd1 vssd1 vccd1 vccd1 _06060_ sky130_fd_sc_hd__a221o_1
XANTENNA__14665__RESET_B net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_107_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07734__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13968_ clknet_leaf_106_clk _00746_ net1223 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06956__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12919_ net1808 net205 net484 vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__mux2_1
X_13899_ clknet_leaf_43_clk net1487 net1151 vssd1 vssd1 vccd1 vccd1 keypad.decode.sticky\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11833__A2 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06675__B _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11073__S net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08110_ datapath.rf.registers\[27\]\[8\] net809 net800 datapath.rf.registers\[15\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02946_ sky130_fd_sc_hd__a22o_1
X_09090_ _02025_ net554 net550 vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__or3_1
X_08041_ _01602_ _01784_ vssd1 vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__nor2_1
Xhold902 datapath.rf.registers\[26\]\[9\] vssd1 vssd1 vccd1 vccd1 net2250 sky130_fd_sc_hd__dlygate4sd3_1
Xhold913 datapath.rf.registers\[1\]\[11\] vssd1 vssd1 vccd1 vccd1 net2261 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold924 datapath.rf.registers\[17\]\[7\] vssd1 vssd1 vccd1 vccd1 net2272 sky130_fd_sc_hd__dlygate4sd3_1
Xhold935 datapath.rf.registers\[19\]\[30\] vssd1 vssd1 vccd1 vccd1 net2283 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_6_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09560__B1_N _04338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold946 datapath.rf.registers\[6\]\[6\] vssd1 vssd1 vccd1 vccd1 net2294 sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 datapath.rf.registers\[25\]\[23\] vssd1 vssd1 vccd1 vccd1 net2305 sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 datapath.rf.registers\[2\]\[22\] vssd1 vssd1 vccd1 vccd1 net2316 sky130_fd_sc_hd__dlygate4sd3_1
X_09992_ _04821_ _04822_ _04827_ _04721_ vssd1 vssd1 vccd1 vccd1 _04828_ sky130_fd_sc_hd__a31o_1
XANTENNA__10941__A net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06776__A1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold979 datapath.rf.registers\[27\]\[16\] vssd1 vssd1 vccd1 vccd1 net2327 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07973__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08943_ net575 _03777_ _03778_ _03769_ vssd1 vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__a22o_1
XFILLER_88_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07953__C net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_15_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_15_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_4_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11248__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10152__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08874_ _03708_ _03709_ net451 vssd1 vssd1 vccd1 vccd1 _03710_ sky130_fd_sc_hd__mux2_1
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07725__B1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07825_ _02660_ vssd1 vssd1 vccd1 vccd1 _02661_ sky130_fd_sc_hd__inv_2
XFILLER_151_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout466_A _01701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07756_ datapath.rf.registers\[5\]\[15\] net819 net813 datapath.rf.registers\[23\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__a22o_1
XANTENNA__06866__A net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06707_ datapath.ru.latched_instruction\[4\] datapath.ru.latched_instruction\[0\]
+ datapath.ru.latched_instruction\[1\] _01545_ vssd1 vssd1 vccd1 vccd1 _01546_ sky130_fd_sc_hd__nor4_1
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07687_ datapath.rf.registers\[0\]\[17\] net870 _02521_ vssd1 vssd1 vccd1 vccd1 _02523_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_13_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09426_ net327 _04033_ _04261_ net379 vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__a211o_1
X_06638_ mmio.memload_or_instruction\[31\] net1050 vssd1 vssd1 vccd1 vccd1 _01477_
+ sky130_fd_sc_hd__and2_2
XFILLER_12_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09357_ _04191_ _04192_ _03661_ net325 vssd1 vssd1 vccd1 vccd1 _04193_ sky130_fd_sc_hd__o2bb2a_1
X_06569_ datapath.ru.latched_instruction\[2\] vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout800_A _01772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12807__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout421_X net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout519_X net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08308_ datapath.rf.registers\[4\]\[4\] net864 net825 datapath.rf.registers\[6\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__a22o_1
XFILLER_60_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09288_ _02467_ _02523_ net443 vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__mux2_1
X_08239_ _03070_ _03071_ _03073_ _03074_ vssd1 vssd1 vccd1 vccd1 _03075_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_134_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12537__B1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07984__X _02820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07008__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11250_ net275 net2168 net420 vssd1 vssd1 vccd1 vccd1 _00299_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout790_X net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout888_X net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10201_ net1041 _05034_ _05036_ net640 vssd1 vssd1 vccd1 vccd1 _05037_ sky130_fd_sc_hd__a211o_1
XFILLER_106_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11181_ net284 net1611 net424 vssd1 vssd1 vccd1 vccd1 _00233_ sky130_fd_sc_hd__mux2_1
XFILLER_107_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06767__A1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10132_ _01702_ _04023_ _04967_ net1040 vssd1 vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__o211a_1
XFILLER_0_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11760__B2 _02385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11158__S net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10063_ _04898_ _04893_ vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__and2b_1
XFILLER_76_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07716__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input27_A DAT_I[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10997__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13822_ clknet_leaf_115_clk _00631_ net1189 vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12068__A2 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13753_ clknet_leaf_88_clk _00562_ net1253 vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__dfrtp_1
X_10965_ datapath.mulitply_result\[1\] net598 net621 vssd1 vssd1 vccd1 vccd1 _05702_
+ sky130_fd_sc_hd__a21o_1
XFILLER_16_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08141__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12704_ _06532_ _06533_ vssd1 vssd1 vccd1 vccd1 _00942_ sky130_fd_sc_hd__and2_1
X_13684_ clknet_leaf_94_clk _00494_ net1212 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10896_ net1264 _05636_ vssd1 vssd1 vccd1 vccd1 _05642_ sky130_fd_sc_hd__xnor2_1
X_12635_ _06471_ _06475_ vssd1 vssd1 vccd1 vccd1 _06476_ sky130_fd_sc_hd__and2_1
XFILLER_12_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07247__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12566_ _06416_ _06417_ _06415_ vssd1 vssd1 vccd1 vccd1 _06419_ sky130_fd_sc_hd__o21ai_1
XFILLER_8_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11517_ _05320_ _05741_ vssd1 vssd1 vccd1 vccd1 _05742_ sky130_fd_sc_hd__or2_1
X_14305_ clknet_leaf_64_clk _01010_ net1239 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[25\]
+ sky130_fd_sc_hd__dfrtp_4
X_12497_ net236 net1710 net507 vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__mux2_1
XFILLER_7_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14236_ clknet_leaf_122_clk datapath.multiplication_module.multiplier_i_n\[4\] net1214
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i\[4\] sky130_fd_sc_hd__dfrtp_1
Xhold209 datapath.rf.registers\[13\]\[25\] vssd1 vssd1 vccd1 vccd1 net1557 sky130_fd_sc_hd__dlygate4sd3_1
X_11448_ net1784 net300 net406 vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__mux2_1
XFILLER_137_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14167_ clknet_leaf_69_clk _00922_ net1245 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11379_ net1604 net289 net413 vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__mux2_1
XANTENNA__07955__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11751__B2 _02824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13118_ net205 net2061 net471 vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__mux2_1
X_14098_ clknet_leaf_122_clk _00864_ net1201 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11068__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13049_ net231 net1728 net475 vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__mux2_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07707__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1260 net1261 vssd1 vssd1 vccd1 vccd1 net1260 sky130_fd_sc_hd__clkbuf_4
Xfanout1271 screen.counter.ct\[15\] vssd1 vssd1 vccd1 vccd1 net1271 sky130_fd_sc_hd__buf_2
Xfanout1282 net1284 vssd1 vssd1 vccd1 vccd1 net1282 sky130_fd_sc_hd__buf_2
XFILLER_94_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1293 _01436_ vssd1 vssd1 vccd1 vccd1 net1293 sky130_fd_sc_hd__clkbuf_2
X_07610_ datapath.rf.registers\[9\]\[18\] net981 net943 vssd1 vssd1 vccd1 vccd1 _02446_
+ sky130_fd_sc_hd__and3_1
X_08590_ _03127_ _03173_ vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__nand2b_1
XFILLER_47_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07541_ datapath.rf.registers\[10\]\[20\] net706 net683 datapath.rf.registers\[27\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__a22o_1
XFILLER_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11806__A2 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08132__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07486__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07472_ datapath.rf.registers\[12\]\[21\] net826 net801 datapath.rf.registers\[3\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__a22o_1
XFILLER_34_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09211_ _03894_ _03895_ net341 vssd1 vssd1 vccd1 vccd1 _04047_ sky130_fd_sc_hd__mux2_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09142_ net556 _03976_ _03977_ _03952_ net632 vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__a32o_2
XANTENNA__07238__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09632__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07948__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09073_ _03906_ _03908_ net319 vssd1 vssd1 vccd1 vccd1 _03909_ sky130_fd_sc_hd__mux2_1
XFILLER_147_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12519__B1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08024_ datapath.rf.registers\[14\]\[10\] net776 net768 datapath.rf.registers\[24\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__a22o_1
XFILLER_151_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold710 datapath.rf.registers\[0\]\[8\] vssd1 vssd1 vccd1 vccd1 net2058 sky130_fd_sc_hd__dlygate4sd3_1
Xhold721 datapath.rf.registers\[12\]\[27\] vssd1 vssd1 vccd1 vccd1 net2069 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10942__Y _05682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold732 datapath.rf.registers\[30\]\[19\] vssd1 vssd1 vccd1 vccd1 net2080 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold743 datapath.rf.registers\[17\]\[10\] vssd1 vssd1 vccd1 vccd1 net2091 sky130_fd_sc_hd__dlygate4sd3_1
Xhold754 datapath.rf.registers\[16\]\[18\] vssd1 vssd1 vccd1 vccd1 net2102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold765 datapath.rf.registers\[1\]\[27\] vssd1 vssd1 vccd1 vccd1 net2113 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold776 datapath.rf.registers\[22\]\[23\] vssd1 vssd1 vccd1 vccd1 net2124 sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 datapath.rf.registers\[26\]\[6\] vssd1 vssd1 vccd1 vccd1 net2135 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11742__B2 _03292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08779__C _03613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07309__X _02145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09975_ _04735_ _04810_ vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__nand2_1
XANTENNA__07410__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold798 datapath.rf.registers\[10\]\[1\] vssd1 vssd1 vccd1 vccd1 net2146 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08926_ _03418_ net577 net546 _01889_ vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__o211a_1
X_08857_ _03689_ _03692_ net342 vssd1 vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout750_A _01804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout469_X net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout848_A _01737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07808_ datapath.rf.registers\[25\]\[14\] net842 net831 datapath.rf.registers\[14\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02644_ sky130_fd_sc_hd__a22o_1
XFILLER_44_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08788_ _01637_ net576 vssd1 vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__nand2_1
XFILLER_73_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07739_ datapath.rf.registers\[19\]\[16\] net730 _02574_ net786 vssd1 vssd1 vccd1
+ vccd1 _02575_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout636_X net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_886 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10750_ _01640_ _05516_ vssd1 vssd1 vccd1 vccd1 _05517_ sky130_fd_sc_hd__nor2_4
XANTENNA__07477__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06883__X _01719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09409_ _02660_ net553 net549 vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__or3_1
X_10681_ _05444_ _05498_ vssd1 vssd1 vccd1 vccd1 _05499_ sky130_fd_sc_hd__nand2_1
XANTENNA__07882__C1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09764__A1_N net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout803_X net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11441__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12420_ net1413 net130 _06357_ vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__a21o_1
XANTENNA__07229__A2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09623__B1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12351_ net230 _04891_ vssd1 vssd1 vccd1 vccd1 _06317_ sky130_fd_sc_hd__nor2_1
X_11302_ net177 net1993 net525 vssd1 vssd1 vccd1 vccd1 _00350_ sky130_fd_sc_hd__mux2_1
XANTENNA__10784__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12282_ datapath.PC\[7\] net309 _06265_ _06267_ vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__a22o_1
XFILLER_135_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14021_ clknet_leaf_78_clk _00790_ net1249 vssd1 vssd1 vccd1 vccd1 datapath.PC\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11233_ net196 net2474 net528 vssd1 vssd1 vccd1 vccd1 _00283_ sky130_fd_sc_hd__mux2_1
XFILLER_153_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10581__A _01934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11164_ net206 net1751 net530 vssd1 vssd1 vccd1 vccd1 _00217_ sky130_fd_sc_hd__mux2_1
XFILLER_106_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10115_ _04868_ _04869_ _04872_ vssd1 vssd1 vccd1 vccd1 _04951_ sky130_fd_sc_hd__o21ai_1
XFILLER_95_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11095_ net212 net1764 net535 vssd1 vssd1 vccd1 vccd1 _00152_ sky130_fd_sc_hd__mux2_1
XFILLER_122_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_147_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10046_ _04831_ _04881_ vssd1 vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__nor2_1
XANTENNA__06777__Y _01614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold70 net58 vssd1 vssd1 vccd1 vccd1 net1418 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07165__B2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold81 screen.controlBus\[25\] vssd1 vssd1 vccd1 vccd1 net1429 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 net120 vssd1 vssd1 vccd1 vccd1 net1440 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13805_ clknet_leaf_76_clk _00614_ net1247 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11997_ _05792_ _05832_ _06040_ vssd1 vssd1 vccd1 vccd1 _06041_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_67_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07889__X _02725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13736_ clknet_leaf_43_clk _00546_ net1150 vssd1 vssd1 vccd1 vccd1 keypad.decode.push
+ sky130_fd_sc_hd__dfrtp_1
X_10948_ datapath.mulitply_result\[31\] net597 net617 vssd1 vssd1 vccd1 vccd1 _05687_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__07468__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10879_ _01505_ net617 _05626_ _05627_ vssd1 vssd1 vccd1 vccd1 _05628_ sky130_fd_sc_hd__a22o_2
X_13667_ clknet_leaf_120_clk _00477_ net1193 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06953__B _01666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11351__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12618_ datapath.mulitply_result\[18\] datapath.multiplication_module.multiplicand_i\[18\]
+ vssd1 vssd1 vccd1 vccd1 _06462_ sky130_fd_sc_hd__or2_1
XFILLER_129_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13598_ clknet_leaf_146_clk _00408_ net1062 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_12549_ datapath.mulitply_result\[6\] net505 net501 _06404_ vssd1 vssd1 vccd1 vccd1
+ _00916_ sky130_fd_sc_hd__a22o_1
XFILLER_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_1 _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14219_ clknet_leaf_47_clk datapath.multiplication_module.multiplicand_i_n\[30\]
+ net1175 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07928__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout508 net509 vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__clkbuf_8
Xfanout519 net521 vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_111_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09760_ _03510_ _03718_ net623 _03512_ net642 vssd1 vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__o221a_1
XANTENNA__12910__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06972_ net912 net907 vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__and2_1
XFILLER_98_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06968__X _01804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08711_ net558 _03418_ vssd1 vssd1 vccd1 vccd1 _03547_ sky130_fd_sc_hd__nor2_1
X_09691_ net376 _04126_ _04526_ net331 vssd1 vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__o211a_1
Xfanout1090 net1091 vssd1 vssd1 vccd1 vccd1 net1090 sky130_fd_sc_hd__buf_2
XFILLER_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08642_ _01912_ _03476_ _01860_ vssd1 vssd1 vccd1 vccd1 _03478_ sky130_fd_sc_hd__o21ai_2
XFILLER_82_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08573_ datapath.rf.registers\[7\]\[0\] net968 _01820_ vssd1 vssd1 vccd1 vccd1 _03409_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout164_A net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07524_ datapath.rf.registers\[30\]\[20\] net834 net806 datapath.rf.registers\[28\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__a22o_1
XFILLER_81_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07459__A2 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07455_ datapath.rf.registers\[5\]\[21\] net945 net931 vssd1 vssd1 vccd1 vccd1 _02291_
+ sky130_fd_sc_hd__and3_1
XANTENNA__11261__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout429_A _05716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07386_ datapath.rf.registers\[29\]\[23\] net675 net660 datapath.rf.registers\[5\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__a22o_1
XFILLER_136_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09125_ _02169_ net553 net549 vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_98_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1240_A net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07092__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09056_ _03666_ _03890_ _03891_ _03880_ vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__a22o_1
XFILLER_124_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09908__A1 _01611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08007_ datapath.rf.registers\[14\]\[10\] net830 net809 datapath.rf.registers\[27\]\[10\]
+ _02831_ vssd1 vssd1 vccd1 vccd1 _02843_ sky130_fd_sc_hd__a221o_1
XANTENNA__13850__SET_B net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold540 datapath.rf.registers\[15\]\[12\] vssd1 vssd1 vccd1 vccd1 net1888 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold551 datapath.rf.registers\[18\]\[8\] vssd1 vssd1 vccd1 vccd1 net1899 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07919__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold562 datapath.rf.registers\[19\]\[10\] vssd1 vssd1 vccd1 vccd1 net1910 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold573 datapath.rf.registers\[24\]\[8\] vssd1 vssd1 vccd1 vccd1 net1921 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold584 datapath.rf.registers\[5\]\[4\] vssd1 vssd1 vccd1 vccd1 net1932 sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 datapath.rf.registers\[6\]\[29\] vssd1 vssd1 vccd1 vccd1 net1943 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout965_A net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12820__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09958_ _04767_ _04793_ _04766_ vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_129_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08909_ datapath.PC\[20\] _03744_ vssd1 vssd1 vccd1 vccd1 _03745_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout753_X net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06597__Y _00004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09889_ datapath.PC\[23\] net594 _04723_ _04724_ vssd1 vssd1 vccd1 vccd1 _04725_
+ sky130_fd_sc_hd__a211o_1
XANTENNA__11436__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1240 datapath.rf.registers\[17\]\[14\] vssd1 vssd1 vccd1 vccd1 net2588 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1251 datapath.rf.registers\[14\]\[14\] vssd1 vssd1 vccd1 vccd1 net2599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1262 datapath.rf.registers\[15\]\[11\] vssd1 vssd1 vccd1 vccd1 net2610 sky130_fd_sc_hd__dlygate4sd3_1
X_11920_ screen.register.currentYbus\[21\] net160 vssd1 vssd1 vccd1 vccd1 _05977_
+ sky130_fd_sc_hd__nand2_1
Xhold1273 datapath.rf.registers\[28\]\[26\] vssd1 vssd1 vccd1 vccd1 net2621 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07698__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1284 datapath.rf.registers\[20\]\[9\] vssd1 vssd1 vccd1 vccd1 net2632 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1295 datapath.rf.registers\[25\]\[27\] vssd1 vssd1 vccd1 vccd1 net2643 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11851_ net1010 _05910_ _05927_ _05928_ _05929_ vssd1 vssd1 vccd1 vccd1 _05930_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_142_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout920_X net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ _04561_ _05561_ net899 vssd1 vssd1 vccd1 vccd1 _05562_ sky130_fd_sc_hd__mux2_1
X_14570_ clknet_leaf_60_clk _01275_ net1169 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[21\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11782_ keypad.apps.app_c\[0\] keypad.apps.app_c\[1\] _05880_ _05895_ button\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05896_ sky130_fd_sc_hd__a2111o_1
XFILLER_14_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11675__A2_N _05885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10733_ net1544 net568 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[19\]
+ sky130_fd_sc_hd__and2_1
X_13521_ clknet_leaf_40_clk _00331_ net1140 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11171__S net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13452_ clknet_leaf_14_clk _00262_ net1103 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10664_ _05451_ _05482_ vssd1 vssd1 vccd1 vccd1 _05483_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_11_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07870__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_14_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10206__A1 _04600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12403_ _05960_ net156 vssd1 vssd1 vccd1 vccd1 _06349_ sky130_fd_sc_hd__nor2_1
XANTENNA__10863__X _05614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13383_ clknet_leaf_145_clk _00193_ net1087 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10595_ net1522 _01419_ _05291_ datapath.ru.n_memwrite vssd1 vssd1 vccd1 vccd1 _00002_
+ sky130_fd_sc_hd__a22o_1
X_12334_ _05002_ net307 _06304_ _06253_ _05631_ vssd1 vssd1 vccd1 vccd1 _06305_ sky130_fd_sc_hd__a32o_1
XANTENNA__07622__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13098__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12265_ _05002_ net307 _06251_ _06253_ _05276_ vssd1 vssd1 vccd1 vccd1 _06255_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_128_Right_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14004_ clknet_leaf_108_clk net1371 net1219 vssd1 vssd1 vccd1 vccd1 screen.counter.ack3
+ sky130_fd_sc_hd__dfrtp_1
X_11216_ net281 net1899 net529 vssd1 vssd1 vccd1 vccd1 _00266_ sky130_fd_sc_hd__mux2_1
XFILLER_123_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12196_ screen.counter.currentCt\[1\] _06205_ screen.counter.currentCt\[2\] vssd1
+ vssd1 vccd1 vccd1 _06208_ sky130_fd_sc_hd__a21oi_1
Xoutput60 net60 vssd1 vssd1 vccd1 vccd1 ADR_O[28] sky130_fd_sc_hd__buf_2
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 ADR_O[9] sky130_fd_sc_hd__buf_2
XANTENNA__08583__B1 _03384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14020__RESET_B net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput82 net82 vssd1 vssd1 vccd1 vccd1 DAT_O[18] sky130_fd_sc_hd__buf_2
X_11147_ net291 net2135 net530 vssd1 vssd1 vccd1 vccd1 _00200_ sky130_fd_sc_hd__mux2_1
Xoutput93 net93 vssd1 vssd1 vccd1 vccd1 DAT_O[28] sky130_fd_sc_hd__buf_2
XANTENNA__10390__A0 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11078_ net295 net2077 net534 vssd1 vssd1 vccd1 vccd1 _00135_ sky130_fd_sc_hd__mux2_1
XANTENNA__08335__A0 _03150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11346__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10029_ _04740_ _04808_ vssd1 vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__xnor2_2
XANTENNA__07689__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10142__B1 _01702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11870__A _03170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06964__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13719_ clknet_leaf_127_clk _00529_ net1209 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10445__B2 net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11081__S net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07310__A1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07240_ _02074_ _02075_ vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__or2_1
XANTENNA__07861__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07498__C net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07171_ datapath.rf.registers\[14\]\[27\] net983 net919 vssd1 vssd1 vccd1 vccd1 _02007_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12905__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07613__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08810__A1 _03228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12206__A _06168_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08403__B net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout305 _05523_ vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout316 _05905_ vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__clkbuf_2
Xfanout327 net328 vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__buf_2
X_09812_ _03484_ _03597_ _03482_ vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__a21oi_1
XFILLER_141_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout338 net339 vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__buf_2
Xfanout349 net350 vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__buf_2
X_06955_ net914 net911 vssd1 vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__nand2_1
X_09743_ net607 _04565_ _04578_ net555 vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__o211a_1
XANTENNA__08326__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout281_A _05554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11256__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10160__S net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09674_ _03539_ net629 net646 vssd1 vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__a21o_1
XFILLER_55_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06886_ net955 _01712_ vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__and2_1
X_08625_ _02241_ _03460_ _02242_ vssd1 vssd1 vccd1 vccd1 _03461_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_38_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1190_A net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout546_A _03759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08556_ datapath.rf.registers\[8\]\[0\] net697 _03389_ _03390_ _03391_ vssd1 vssd1
+ vccd1 vccd1 _03392_ sky130_fd_sc_hd__a2111o_1
X_07507_ datapath.rf.registers\[5\]\[20\] net945 net932 vssd1 vssd1 vccd1 vccd1 _02343_
+ sky130_fd_sc_hd__and3_1
X_08487_ _01663_ _01703_ vssd1 vssd1 vccd1 vccd1 _03323_ sky130_fd_sc_hd__and2_1
XFILLER_23_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout713_A _01817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07438_ datapath.rf.registers\[22\]\[22\] net734 net718 datapath.rf.registers\[20\]\[22\]
+ _02273_ vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__a221o_1
XANTENNA__07852__A2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07369_ datapath.rf.registers\[31\]\[23\] net794 _02200_ _02201_ _02202_ vssd1 vssd1
+ vccd1 vccd1 _02205_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout501_X net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1243_X net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12815__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09108_ _03495_ net627 net624 _03496_ net644 vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__a221o_1
XANTENNA__07065__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11939__B screen.counter.ack vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10380_ net558 _03418_ net623 vssd1 vssd1 vccd1 vccd1 _05216_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07604__A2 _02438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09039_ _02069_ _02125_ net442 vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__mux2_1
XFILLER_117_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12050_ screen.register.currentXbus\[28\] _05772_ _05837_ screen.register.currentYbus\[20\]
+ vssd1 vssd1 vccd1 vccd1 _06091_ sky130_fd_sc_hd__a22o_1
Xhold370 datapath.rf.registers\[21\]\[19\] vssd1 vssd1 vccd1 vccd1 net1718 sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 datapath.rf.registers\[29\]\[15\] vssd1 vssd1 vccd1 vccd1 net1729 sky130_fd_sc_hd__dlygate4sd3_1
Xhold392 datapath.rf.registers\[6\]\[5\] vssd1 vssd1 vccd1 vccd1 net1740 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_120_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11001_ _01649_ _03264_ vssd1 vssd1 vccd1 vccd1 _05707_ sky130_fd_sc_hd__nand2_1
XFILLER_77_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout850 _01735_ vssd1 vssd1 vccd1 vccd1 net850 sky130_fd_sc_hd__buf_2
Xfanout861 net863 vssd1 vssd1 vccd1 vccd1 net861 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_144_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout872 _01723_ vssd1 vssd1 vccd1 vccd1 net872 sky130_fd_sc_hd__buf_4
Xfanout883 _01719_ vssd1 vssd1 vccd1 vccd1 net883 sky130_fd_sc_hd__buf_6
Xfanout894 net896 vssd1 vssd1 vccd1 vccd1 net894 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11166__S net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08317__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06768__B _01603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12952_ net205 net1890 net394 vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__mux2_1
XANTENNA__08868__A1 _02857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1070 datapath.rf.registers\[20\]\[4\] vssd1 vssd1 vccd1 vccd1 net2418 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1081 datapath.rf.registers\[25\]\[12\] vssd1 vssd1 vccd1 vccd1 net2429 sky130_fd_sc_hd__dlygate4sd3_1
X_11903_ _02633_ screen.counter.ack vssd1 vssd1 vccd1 vccd1 _05966_ sky130_fd_sc_hd__or2_1
Xhold1092 screen.counter.currentCt\[19\] vssd1 vssd1 vccd1 vccd1 net2440 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10858__X _05610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ net233 net2003 net398 vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14622_ clknet_leaf_150_clk _01327_ net1061 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11834_ _05760_ _05816_ _05850_ _05819_ vssd1 vssd1 vccd1 vccd1 _05913_ sky130_fd_sc_hd__o31a_1
XANTENNA__09817__B1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06784__A _01611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10427__A1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13522__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11765_ net1482 net146 net140 _02145_ vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__a22o_1
X_14553_ clknet_leaf_31_clk _01258_ net1122 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13504_ clknet_leaf_135_clk _00314_ net1104 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10716_ net463 net573 _05510_ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[4\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_14_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11696_ _04932_ net155 net149 net1404 vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__a22o_1
X_14484_ clknet_leaf_128_clk _01189_ net1209 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10647_ _05450_ _05465_ _05431_ _05448_ vssd1 vssd1 vccd1 vccd1 _05467_ sky130_fd_sc_hd__o211ai_1
XANTENNA__10593__X _05416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13435_ clknet_leaf_38_clk _00245_ net1145 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_139_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07056__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13366_ clknet_leaf_142_clk _00176_ net1094 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10578_ net566 _01889_ _01981_ vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__nand3_1
XANTENNA__10753__B _04338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12317_ _05602_ _06253_ _06292_ net191 vssd1 vssd1 vccd1 vccd1 _06293_ sky130_fd_sc_hd__o2bb2a_1
X_13297_ clknet_leaf_38_clk _00107_ net1141 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12248_ screen.counter.currentCt\[20\] _06238_ screen.counter.currentCt\[21\] vssd1
+ vssd1 vccd1 vccd1 _06241_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_75_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12179_ _06159_ _06172_ _06178_ vssd1 vssd1 vccd1 vccd1 _06198_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06959__A _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09335__A net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11076__S net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08308__B1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06740_ net1004 net1020 _01578_ _01577_ vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__a31o_2
X_06671_ mmio.memload_or_instruction\[15\] net1048 vssd1 vssd1 vccd1 vccd1 _01510_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_35_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08410_ datapath.rf.registers\[24\]\[2\] _01712_ net930 vssd1 vssd1 vccd1 vccd1 _03246_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09341__Y _04177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09390_ _02418_ net440 _04151_ net363 vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_106_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08341_ datapath.rf.registers\[2\]\[3\] net988 net949 vssd1 vssd1 vccd1 vccd1 _03177_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08087__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07295__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08272_ datapath.rf.registers\[17\]\[5\] net747 net676 datapath.rf.registers\[29\]\[5\]
+ _03106_ vssd1 vssd1 vccd1 vccd1 _03108_ sky130_fd_sc_hd__a221o_1
XANTENNA__07834__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06981__X _01817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07223_ datapath.rf.registers\[23\]\[26\] net940 net921 vssd1 vssd1 vccd1 vccd1 _02059_
+ sky130_fd_sc_hd__and3_1
XFILLER_20_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout127_A _06369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07047__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12040__B1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07154_ datapath.rf.registers\[30\]\[28\] net760 net674 datapath.rf.registers\[7\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__a22o_1
XFILLER_145_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08795__B1 _01779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07085_ datapath.rf.registers\[28\]\[29\] net804 net801 datapath.rf.registers\[3\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__a22o_1
XFILLER_121_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout496_A _06550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12343__B2 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08011__A2 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout135 _05934_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1203_A net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06869__A _01579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout146 net147 vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__buf_1
XANTENNA_input1_A ACK_I vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout157 _06335_ vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__clkbuf_2
Xfanout168 net169 vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__clkbuf_2
Xfanout179 _05670_ vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__buf_1
X_07987_ _02809_ _02810_ _02817_ _02822_ vssd1 vssd1 vccd1 vccd1 _02823_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_126_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_126_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06938_ datapath.rf.registers\[15\]\[31\] net799 net796 datapath.rf.registers\[29\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__a22o_1
X_09726_ _04540_ _04560_ _04558_ vssd1 vssd1 vccd1 vccd1 _04562_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_2_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09899__B _04727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout830_A net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09657_ _03429_ _03563_ vssd1 vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__and2_1
X_06869_ _01579_ _01703_ vssd1 vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__and2_1
XFILLER_82_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout928_A _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08608_ _03439_ _03442_ _02773_ vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__o21bai_1
XFILLER_43_748 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09588_ _04422_ _04423_ _03642_ vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__a21oi_1
XFILLER_82_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07052__X _01888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10409__A1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10409__B2 _03604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08539_ datapath.rf.registers\[9\]\[0\] _01716_ _01756_ datapath.rf.registers\[5\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__a22o_1
XANTENNA__08078__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout716_X net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11550_ screen.counter.ct\[0\] screen.counter.ct\[1\] vssd1 vssd1 vccd1 vccd1 _05774_
+ sky130_fd_sc_hd__nand2b_1
XANTENNA__07987__X _02823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06891__X _01727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10501_ _05324_ _05330_ vssd1 vssd1 vccd1 vccd1 _05331_ sky130_fd_sc_hd__nor2_1
X_11481_ net303 net1974 net513 vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__mux2_1
XFILLER_137_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13220_ clknet_leaf_17_clk _00030_ net1109 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_137_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10432_ datapath.PC\[1\] _05267_ _05212_ vssd1 vssd1 vccd1 vccd1 _05268_ sky130_fd_sc_hd__mux2_1
XFILLER_136_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08786__A0 _01647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13151_ net1788 net203 net383 vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__mux2_1
X_10363_ datapath.PC\[8\] net1254 _05195_ _05198_ vssd1 vssd1 vccd1 vccd1 _05199_
+ sky130_fd_sc_hd__o22a_1
XFILLER_136_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08250__A2 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12102_ _06124_ _06139_ vssd1 vssd1 vccd1 vccd1 _06140_ sky130_fd_sc_hd__nor2_1
XFILLER_152_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13082_ net1863 net231 net386 vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__mux2_1
X_10294_ _03734_ _05129_ net1038 vssd1 vssd1 vccd1 vccd1 _05130_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12334__A1 _05002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08538__B1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12033_ _06021_ _06039_ _06074_ vssd1 vssd1 vccd1 vccd1 _06075_ sky130_fd_sc_hd__or3_1
XFILLER_151_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06779__A net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_8_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout680 _01828_ vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__clkbuf_4
Xfanout691 _01824_ vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13984_ clknet_leaf_108_clk _00761_ net1221 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08994__A net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12935_ net293 net2152 net394 vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__mux2_1
XFILLER_34_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12866_ net304 net1646 net401 vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__mux2_1
XANTENNA__07403__A net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14605_ clknet_leaf_131_clk _01310_ net1113 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11817_ _01527_ net1015 net313 net333 datapath.ru.latched_instruction\[23\] vssd1
+ vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__a32o_1
XANTENNA__08069__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12797_ net2385 net207 net493 vssd1 vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__mux2_1
XANTENNA__07122__B net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14536_ clknet_leaf_60_clk _01241_ net1169 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07816__A2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11748_ net1488 net144 net139 _02980_ vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__a22o_1
X_14467_ clknet_leaf_120_clk _01172_ net1200 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11679_ _05199_ net152 net151 net1407 vssd1 vssd1 vccd1 vccd1 _00564_ sky130_fd_sc_hd__a22o_1
XANTENNA__06961__B _01666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13418_ clknet_leaf_60_clk _00228_ net1169 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_77_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14398_ clknet_leaf_148_clk _01103_ net1061 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_127_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13349_ clknet_leaf_139_clk _00159_ net1191 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08521__X _03357_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08529__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07910_ _02731_ _02732_ _02744_ _02745_ vssd1 vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__or4_1
X_08890_ _03479_ net609 net605 _03725_ vssd1 vssd1 vccd1 vccd1 _03726_ sky130_fd_sc_hd__a211o_1
XANTENNA__10336__B1 _04239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07201__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07841_ datapath.rf.registers\[28\]\[14\] net751 net676 datapath.rf.registers\[29\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02677_ sky130_fd_sc_hd__a22o_1
XFILLER_29_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09741__A2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08400__C net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07772_ datapath.rf.registers\[24\]\[15\] net857 net833 datapath.rf.registers\[30\]\[15\]
+ _02593_ vssd1 vssd1 vccd1 vccd1 _02608_ sky130_fd_sc_hd__a221o_1
XANTENNA__06976__X _01812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06723_ _01461_ _01557_ _01559_ _01561_ vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__or4_1
X_09511_ _03263_ _03657_ _04346_ net460 vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_88_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09442_ _02750_ net554 net550 vssd1 vssd1 vccd1 vccd1 _04278_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_88_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06654_ mmio.memload_or_instruction\[20\] net1049 vssd1 vssd1 vccd1 vccd1 _01493_
+ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_4_2_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09373_ net630 _04208_ vssd1 vssd1 vccd1 vccd1 _04209_ sky130_fd_sc_hd__nor2_1
XANTENNA__11106__Y _05716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06585_ keypad.decode.q2 vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__inv_2
XFILLER_12_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08324_ datapath.rf.registers\[18\]\[4\] net722 net675 datapath.rf.registers\[29\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__a22o_1
XANTENNA__07807__A2 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08255_ datapath.rf.registers\[17\]\[5\] net850 net833 datapath.rf.registers\[30\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03091_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout411_A _05730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08480__A2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1153_A net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06871__B _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07206_ datapath.rf.registers\[12\]\[27\] net755 net684 datapath.rf.registers\[27\]\[27\]
+ _02027_ vssd1 vssd1 vccd1 vccd1 _02042_ sky130_fd_sc_hd__a221o_1
XFILLER_137_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xteam_04_1300 vssd1 vssd1 vccd1 vccd1 team_04_1300/HI gpio_oeb[9] sky130_fd_sc_hd__conb_1
X_08186_ datapath.rf.registers\[4\]\[7\] net716 net696 datapath.rf.registers\[8\]\[7\]
+ _03021_ vssd1 vssd1 vccd1 vccd1 _03022_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_119_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xteam_04_1311 vssd1 vssd1 vccd1 vccd1 team_04_1311/HI gpio_out[0] sky130_fd_sc_hd__conb_1
Xteam_04_1322 vssd1 vssd1 vccd1 vccd1 team_04_1322/HI gpio_out[26] sky130_fd_sc_hd__conb_1
Xteam_04_1333 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] team_04_1333/LO sky130_fd_sc_hd__conb_1
X_07137_ datapath.rf.registers\[5\]\[28\] _01756_ _01958_ _01960_ _01961_ vssd1 vssd1
+ vccd1 vccd1 _01973_ sky130_fd_sc_hd__a2111o_1
XFILLER_119_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xteam_04_1344 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] team_04_1344/LO sky130_fd_sc_hd__conb_1
XANTENNA__08232__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1039_X net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11776__Y _05894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07440__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07068_ datapath.rf.registers\[24\]\[30\] net768 net728 datapath.rf.registers\[25\]\[30\]
+ _01893_ vssd1 vssd1 vccd1 vccd1 _01904_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout780_A _01794_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09193__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout666_X net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09709_ net328 _04385_ _03623_ vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__o21ai_1
X_10981_ net2216 net262 net435 vssd1 vssd1 vccd1 vccd1 _00046_ sky130_fd_sc_hd__mux2_1
XANTENNA__08299__A2 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout833_X net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09496__A1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11444__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12720_ _06541_ _06542_ _06531_ vssd1 vssd1 vccd1 vccd1 _06543_ sky130_fd_sc_hd__o21a_1
X_12651_ _06481_ _06485_ _06488_ vssd1 vssd1 vccd1 vccd1 _06490_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_26_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09248__A1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11602_ _05773_ _05776_ _05778_ vssd1 vssd1 vccd1 vccd1 _05826_ sky130_fd_sc_hd__or3_1
XANTENNA__09799__A2 _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12582_ _06430_ _06431_ vssd1 vssd1 vccd1 vccd1 _06432_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_156_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14321_ clknet_leaf_35_clk _01026_ net1127 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11533_ _05294_ net1006 vssd1 vssd1 vccd1 vccd1 _05757_ sky130_fd_sc_hd__nor2_2
XANTENNA__10584__A _02824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08471__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12004__B1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14252_ clknet_leaf_16_clk _00957_ net1106 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11464_ net2369 net233 net406 vssd1 vssd1 vccd1 vccd1 _00502_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_152_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10415_ _03321_ net452 net457 vssd1 vssd1 vccd1 vccd1 _05251_ sky130_fd_sc_hd__a21oi_1
X_13203_ clknet_leaf_35_clk _00013_ net1130 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_137_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14183_ clknet_leaf_51_clk _00938_ net1182 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10871__X _05621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08223__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11395_ net1683 net220 net410 vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__mux2_1
X_10346_ _03737_ _05181_ net1039 vssd1 vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07431__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13134_ net2294 net290 net383 vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__mux2_1
XFILLER_98_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12307__B2 _04239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_72_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09708__C1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13065_ net1564 net302 net389 vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__mux2_1
X_10277_ _04848_ _04850_ vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__nand2b_1
XANTENNA__08501__B net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12016_ screen.register.currentYbus\[18\] _05773_ _05790_ screen.register.currentXbus\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06059_ sky130_fd_sc_hd__a22o_1
XFILLER_93_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13967_ clknet_leaf_106_clk _00745_ net1223 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09487__A1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06956__B net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11354__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12918_ net2459 net211 net482 vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__mux2_1
XFILLER_46_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07404__Y _02240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13898_ clknet_leaf_43_clk keypad.decode.sticky_n\[3\] net1151 vssd1 vssd1 vccd1
+ vccd1 keypad.decode.sticky\[3\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09239__A1 _03667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12849_ net236 net2080 net488 vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__mux2_1
XFILLER_15_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08998__A0 _01888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10254__C1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14519_ clknet_leaf_130_clk _01224_ net1114 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08040_ _02862_ _02865_ _02875_ net785 datapath.rf.registers\[0\]\[10\] vssd1 vssd1
+ vccd1 vccd1 _02876_ sky130_fd_sc_hd__o32a_4
Xhold903 datapath.rf.registers\[30\]\[5\] vssd1 vssd1 vccd1 vccd1 net2251 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14116__D datapath.ack_mul vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08214__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold914 datapath.rf.registers\[31\]\[12\] vssd1 vssd1 vccd1 vccd1 net2262 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12913__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold925 screen.register.currentYbus\[1\] vssd1 vssd1 vccd1 vccd1 net2273 sky130_fd_sc_hd__dlygate4sd3_1
Xhold936 datapath.rf.registers\[2\]\[14\] vssd1 vssd1 vccd1 vccd1 net2284 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07422__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold947 datapath.rf.registers\[8\]\[26\] vssd1 vssd1 vccd1 vccd1 net2295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold958 datapath.rf.registers\[20\]\[27\] vssd1 vssd1 vccd1 vccd1 net2306 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09991_ _04824_ _04826_ vssd1 vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__nor2_1
Xhold969 datapath.rf.registers\[27\]\[26\] vssd1 vssd1 vccd1 vccd1 net2317 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06776__A2 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08942_ net649 _03777_ net438 vssd1 vssd1 vccd1 vccd1 _03778_ sky130_fd_sc_hd__a21o_1
XANTENNA__10309__B1 net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12214__A _06168_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08411__B net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08873_ net464 net463 net446 vssd1 vssd1 vccd1 vccd1 _03709_ sky130_fd_sc_hd__mux2_1
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08922__B1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07824_ datapath.rf.registers\[0\]\[14\] net871 _02652_ _02659_ vssd1 vssd1 vccd1
+ vccd1 _02660_ sky130_fd_sc_hd__o22a_4
XANTENNA__07027__B net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07755_ datapath.rf.registers\[4\]\[15\] net958 net933 vssd1 vssd1 vccd1 vccd1 _02591_
+ sky130_fd_sc_hd__and3_1
XANTENNA__11264__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10088__A2 _01702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06706_ datapath.ru.latched_instruction\[3\] datapath.ru.latched_instruction\[5\]
+ datapath.ru.latched_instruction\[6\] datapath.ru.latched_instruction\[7\] vssd1
+ vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__or4_1
XANTENNA__07489__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07686_ datapath.rf.registers\[0\]\[17\] net870 _02521_ vssd1 vssd1 vccd1 vccd1 _02522_
+ sky130_fd_sc_hd__o21a_2
X_06637_ net1288 net1283 datapath.ru.latched_instruction\[11\] mmio.memload_or_instruction\[11\]
+ vssd1 vssd1 vccd1 vccd1 _01476_ sky130_fd_sc_hd__or4b_1
X_09425_ net327 _04260_ vssd1 vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_23_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout626_A net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06568_ datapath.ru.latched_instruction\[1\] vssd1 vssd1 vccd1 vccd1 _01409_ sky130_fd_sc_hd__inv_2
XFILLER_12_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09356_ net358 _04184_ _04190_ net325 vssd1 vssd1 vccd1 vccd1 _04192_ sky130_fd_sc_hd__o31a_1
XANTENNA__08426__X _03262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08307_ datapath.rf.registers\[8\]\[4\] net876 net856 datapath.rf.registers\[24\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__a22o_1
XFILLER_21_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09287_ _02365_ _03761_ _04089_ net368 vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout414_X net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09650__A1 _03667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08453__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08238_ datapath.rf.registers\[12\]\[6\] net754 net679 datapath.rf.registers\[6\]\[6\]
+ _03072_ vssd1 vssd1 vccd1 vccd1 _03074_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_134_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12537__A1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08169_ datapath.rf.registers\[9\]\[7\] _01716_ net854 datapath.rf.registers\[19\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03005_ sky130_fd_sc_hd__a22o_1
XANTENNA__12823__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08205__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09402__A1 _03673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10200_ _03747_ _05035_ net1043 vssd1 vssd1 vccd1 vccd1 _05036_ sky130_fd_sc_hd__o21a_1
XANTENNA__07413__B1 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_152_Left_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11180_ net292 net1924 net422 vssd1 vssd1 vccd1 vccd1 _00232_ sky130_fd_sc_hd__mux2_1
XFILLER_69_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout783_X net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10131_ net1265 net469 vssd1 vssd1 vccd1 vccd1 _04967_ sky130_fd_sc_hd__or2_1
XANTENNA__11439__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09166__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10062_ _04894_ _04897_ vssd1 vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__xor2_1
XFILLER_88_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07192__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13821_ clknet_leaf_141_clk _00630_ net1095 vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10579__A _02217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11174__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13752_ clknet_leaf_88_clk _00561_ net1252 vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__dfrtp_1
X_10964_ datapath.PC\[1\] _05267_ net897 vssd1 vssd1 vccd1 vccd1 _05701_ sky130_fd_sc_hd__mux2_1
XANTENNA__09720__X _04556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12703_ columns.count\[0\] _06531_ vssd1 vssd1 vccd1 vccd1 _06533_ sky130_fd_sc_hd__or2_1
XFILLER_44_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13683_ clknet_leaf_36_clk _00493_ net1129 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10895_ net206 net2007 net543 vssd1 vssd1 vccd1 vccd1 _00025_ sky130_fd_sc_hd__mux2_1
X_12634_ net498 _06474_ _06475_ net502 net2584 vssd1 vssd1 vccd1 vccd1 _00930_ sky130_fd_sc_hd__a32o_1
XFILLER_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12565_ _06415_ _06416_ _06417_ vssd1 vssd1 vccd1 vccd1 _06418_ sky130_fd_sc_hd__or3_1
XANTENNA__08444__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14304_ clknet_leaf_133_clk _01009_ net1112 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[24\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_129_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11516_ screen.controlBus\[1\] _05314_ _05318_ screen.controlBus\[0\] vssd1 vssd1
+ vccd1 vccd1 _05741_ sky130_fd_sc_hd__and4b_1
XANTENNA__07652__B1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12496_ net218 net1882 net506 vssd1 vssd1 vccd1 vccd1 _00896_ sky130_fd_sc_hd__mux2_1
XFILLER_8_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14235_ clknet_leaf_123_clk datapath.multiplication_module.multiplier_i_n\[3\] net1214
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i\[3\] sky130_fd_sc_hd__dfrtp_1
X_11447_ net2530 net304 net408 vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__mux2_1
XANTENNA__12733__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07404__B1 _01787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11378_ net1595 net258 net413 vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__mux2_1
X_14166_ clknet_leaf_70_clk _00921_ net1245 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11349__S net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10329_ _04864_ _05164_ vssd1 vssd1 vccd1 vccd1 _05165_ sky130_fd_sc_hd__nand2_1
X_13117_ net211 net2415 net470 vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__mux2_1
X_14097_ clknet_leaf_110_clk _00863_ net1201 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13048_ net237 net1718 net476 vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__mux2_1
XFILLER_121_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1250 net1251 vssd1 vssd1 vccd1 vccd1 net1250 sky130_fd_sc_hd__clkbuf_2
XFILLER_121_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1261 net1262 vssd1 vssd1 vccd1 vccd1 net1261 sky130_fd_sc_hd__buf_2
XANTENNA__11873__A _03123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1272 screen.counter.ct\[14\] vssd1 vssd1 vccd1 vccd1 net1272 sky130_fd_sc_hd__clkbuf_2
Xfanout1283 net1284 vssd1 vssd1 vccd1 vccd1 net1283 sky130_fd_sc_hd__buf_2
Xfanout1294 _01436_ vssd1 vssd1 vccd1 vccd1 net1294 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07183__A2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11084__S net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_80_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07540_ datapath.rf.registers\[13\]\[20\] net691 _02367_ net786 vssd1 vssd1 vccd1
+ vccd1 _02376_ sky130_fd_sc_hd__a211o_1
XFILLER_19_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07471_ datapath.rf.registers\[1\]\[21\] net845 net799 datapath.rf.registers\[15\]\[21\]
+ _02293_ vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__a221o_1
XANTENNA__12908__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09210_ _03666_ _04044_ _04045_ _04035_ vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__a22o_1
XANTENNA__07798__A _02633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_95_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09141_ _03604_ _03953_ _03954_ net608 _03952_ vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__o32a_1
XFILLER_147_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09632__A1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08406__B net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09072_ net343 _03907_ vssd1 vssd1 vccd1 vccd1 _03908_ sky130_fd_sc_hd__or2_1
XANTENNA__07643__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12519__A1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06997__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08023_ datapath.rf.registers\[25\]\[10\] net728 net689 datapath.rf.registers\[31\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_116_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold700 datapath.rf.registers\[20\]\[20\] vssd1 vssd1 vccd1 vccd1 net2048 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_146_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold711 datapath.rf.registers\[16\]\[11\] vssd1 vssd1 vccd1 vccd1 net2059 sky130_fd_sc_hd__dlygate4sd3_1
Xhold722 datapath.rf.registers\[14\]\[26\] vssd1 vssd1 vccd1 vccd1 net2070 sky130_fd_sc_hd__dlygate4sd3_1
Xhold733 datapath.mulitply_result\[8\] vssd1 vssd1 vccd1 vccd1 net2081 sky130_fd_sc_hd__dlygate4sd3_1
Xhold744 datapath.rf.registers\[15\]\[28\] vssd1 vssd1 vccd1 vccd1 net2092 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold755 datapath.rf.registers\[10\]\[18\] vssd1 vssd1 vccd1 vccd1 net2103 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11259__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold766 datapath.rf.registers\[3\]\[12\] vssd1 vssd1 vccd1 vccd1 net2114 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11742__A2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold777 datapath.mulitply_result\[5\] vssd1 vssd1 vccd1 vccd1 net2125 sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 datapath.rf.registers\[17\]\[2\] vssd1 vssd1 vccd1 vccd1 net2136 sky130_fd_sc_hd__dlygate4sd3_1
X_09974_ _04740_ _04743_ _04807_ _04739_ _04737_ vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__a311o_1
Xhold799 datapath.rf.registers\[0\]\[2\] vssd1 vssd1 vccd1 vccd1 net2147 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_33_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08925_ net557 net576 net546 vssd1 vssd1 vccd1 vccd1 _03761_ sky130_fd_sc_hd__o21ai_2
XANTENNA__09699__A1 _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09699__B2 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08856_ _03690_ _03691_ net449 vssd1 vssd1 vccd1 vccd1 _03692_ sky130_fd_sc_hd__mux2_1
XANTENNA__07174__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07807_ datapath.rf.registers\[10\]\[14\] net880 net833 datapath.rf.registers\[30\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02643_ sky130_fd_sc_hd__a22o_1
XFILLER_55_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout743_A net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08787_ _03617_ net378 vssd1 vssd1 vccd1 vccd1 _03623_ sky130_fd_sc_hd__or2_2
XANTENNA_clkbuf_leaf_48_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06921__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07738_ datapath.rf.registers\[22\]\[16\] net734 net694 datapath.rf.registers\[8\]\[16\]
+ _02573_ vssd1 vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__a221o_1
XFILLER_25_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout531_X net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_898 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12818__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07669_ datapath.rf.registers\[28\]\[17\] net929 net920 vssd1 vssd1 vccd1 vccd1 _02505_
+ sky130_fd_sc_hd__and3_1
XFILLER_41_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout629_X net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09408_ _04129_ _04132_ net349 vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__o21ai_1
X_10680_ _05483_ _05490_ _05492_ _05462_ _05497_ vssd1 vssd1 vccd1 vccd1 _05498_ sky130_fd_sc_hd__a221o_1
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09339_ _04167_ _04171_ _04174_ vssd1 vssd1 vccd1 vccd1 _04175_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_109_Right_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_106_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08316__B _01800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12350_ net1263 net310 _06316_ vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__a21o_1
XANTENNA__07634__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11301_ net186 net2643 net523 vssd1 vssd1 vccd1 vccd1 _00349_ sky130_fd_sc_hd__mux2_1
X_12281_ _05002_ net306 _06266_ _06253_ _05544_ vssd1 vssd1 vccd1 vccd1 _06267_ sky130_fd_sc_hd__a32o_1
X_14020_ clknet_leaf_79_clk _00789_ net1254 vssd1 vssd1 vccd1 vccd1 datapath.PC\[10\]
+ sky130_fd_sc_hd__dfrtp_4
X_11232_ net201 net1913 net527 vssd1 vssd1 vccd1 vccd1 _00282_ sky130_fd_sc_hd__mux2_1
XANTENNA__11169__S net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11163_ net211 net1835 net530 vssd1 vssd1 vccd1 vccd1 _00216_ sky130_fd_sc_hd__mux2_1
XFILLER_121_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08051__B net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10114_ net640 _04949_ _04948_ net225 vssd1 vssd1 vccd1 vccd1 _04950_ sky130_fd_sc_hd__a211o_1
X_11094_ net216 net1865 net535 vssd1 vssd1 vccd1 vccd1 _00151_ sky130_fd_sc_hd__mux2_1
XFILLER_49_924 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10045_ _04878_ _04880_ vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_4_10_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06787__A net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold60 net51 vssd1 vssd1 vccd1 vccd1 net1408 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 screen.controlBus\[19\] vssd1 vssd1 vccd1 vccd1 net1419 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 net56 vssd1 vssd1 vccd1 vccd1 net1430 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold93 net41 vssd1 vssd1 vccd1 vccd1 net1441 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13804_ clknet_leaf_74_clk _00613_ net1250 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11996_ _05788_ net998 _05790_ _05794_ vssd1 vssd1 vccd1 vccd1 _06040_ sky130_fd_sc_hd__or4b_1
XFILLER_17_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13735_ clknet_leaf_142_clk _00545_ net1086 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10947_ _03728_ _05685_ net902 vssd1 vssd1 vccd1 vccd1 _05686_ sky130_fd_sc_hd__mux2_2
X_13666_ clknet_leaf_151_clk _00476_ net1053 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07873__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10878_ datapath.mulitply_result\[21\] net615 net652 vssd1 vssd1 vccd1 vccd1 _05627_
+ sky130_fd_sc_hd__o21a_1
XFILLER_31_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12617_ datapath.mulitply_result\[18\] datapath.multiplication_module.multiplicand_i\[18\]
+ vssd1 vssd1 vccd1 vccd1 _06461_ sky130_fd_sc_hd__nand2_1
XFILLER_31_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08417__A2 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10248__S net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13861__RESET_B net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13597_ clknet_leaf_147_clk _00407_ net1088 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_4_14_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_14_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07625__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12548_ _06402_ _06403_ vssd1 vssd1 vccd1 vccd1 _06404_ sky130_fd_sc_hd__xor2_1
XANTENNA_2 _02466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ net258 net1789 net508 vssd1 vssd1 vccd1 vccd1 _00879_ sky130_fd_sc_hd__mux2_1
XFILLER_6_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14218_ clknet_leaf_51_clk datapath.multiplication_module.multiplicand_i_n\[29\]
+ net1175 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11724__A2 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11079__S net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14149_ clknet_leaf_20_clk _00906_ net1163 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_140_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_111_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout509 _06371_ vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_111_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06971_ net914 net909 vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__and2_1
XFILLER_39_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08710_ net559 _03359_ vssd1 vssd1 vccd1 vccd1 _03546_ sky130_fd_sc_hd__nor2_1
X_09690_ net327 _04525_ vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__or2_1
Xfanout1080 net1084 vssd1 vssd1 vccd1 vccd1 net1080 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07156__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07145__X _01981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1091 net1092 vssd1 vssd1 vccd1 vccd1 net1091 sky130_fd_sc_hd__clkbuf_2
X_08641_ _01860_ _01912_ _03476_ vssd1 vssd1 vccd1 vccd1 _03477_ sky130_fd_sc_hd__or3_1
XFILLER_67_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08572_ datapath.rf.registers\[29\]\[0\] net966 _01823_ vssd1 vssd1 vccd1 vccd1 _03408_
+ sky130_fd_sc_hd__and3_1
XFILLER_35_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07523_ datapath.rf.registers\[19\]\[20\] net854 net845 datapath.rf.registers\[1\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__a22o_1
XANTENNA__13949__RESET_B net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout157_A _06335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08510__D1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07454_ datapath.rf.registers\[21\]\[21\] net945 net921 vssd1 vssd1 vccd1 vccd1 _02290_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07864__B1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07385_ datapath.rf.registers\[4\]\[23\] net714 net679 datapath.rf.registers\[6\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__a22o_1
XFILLER_148_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09605__A1 _02961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1066_A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07616__B1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09124_ net356 net355 _03660_ vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__and3_1
XANTENNA__07040__B net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09055_ net649 _03890_ net439 vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_131_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12373__S net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1233_A net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08006_ datapath.rf.registers\[15\]\[10\] net984 net915 vssd1 vssd1 vccd1 vccd1 _02842_
+ sky130_fd_sc_hd__and3_1
Xhold530 datapath.mulitply_result\[16\] vssd1 vssd1 vccd1 vccd1 net1878 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold541 datapath.rf.registers\[13\]\[5\] vssd1 vssd1 vccd1 vccd1 net1889 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout693_A _01824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold552 datapath.rf.registers\[17\]\[1\] vssd1 vssd1 vccd1 vccd1 net1900 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11715__A2 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold563 datapath.rf.registers\[11\]\[17\] vssd1 vssd1 vccd1 vccd1 net1911 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold574 datapath.rf.registers\[25\]\[8\] vssd1 vssd1 vccd1 vccd1 net1922 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1021_X net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold585 datapath.rf.registers\[11\]\[28\] vssd1 vssd1 vccd1 vccd1 net1933 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold596 datapath.rf.registers\[15\]\[5\] vssd1 vssd1 vccd1 vccd1 net1944 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07395__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07991__A _02804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09957_ _04770_ _04792_ _04769_ vssd1 vssd1 vccd1 vccd1 _04793_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout860_A net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout481_X net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout958_A net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08908_ datapath.PC\[19\] _03743_ vssd1 vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_129_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09888_ net1265 net594 vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__and2_1
Xhold1230 datapath.mulitply_result\[31\] vssd1 vssd1 vccd1 vccd1 net2578 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09541__A0 _02913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07147__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1241 datapath.rf.registers\[15\]\[31\] vssd1 vssd1 vccd1 vccd1 net2589 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1252 screen.register.currentXbus\[6\] vssd1 vssd1 vccd1 vccd1 net2600 sky130_fd_sc_hd__dlygate4sd3_1
X_08839_ _01637_ _03671_ vssd1 vssd1 vccd1 vccd1 _03675_ sky130_fd_sc_hd__nand2_1
Xhold1263 datapath.ru.latched_instruction\[8\] vssd1 vssd1 vccd1 vccd1 net2611 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10151__B2 net1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1274 datapath.rf.registers\[3\]\[29\] vssd1 vssd1 vccd1 vccd1 net2622 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout746_X net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1285 datapath.rf.registers\[25\]\[1\] vssd1 vssd1 vccd1 vccd1 net2633 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1296 datapath.rf.registers\[8\]\[5\] vssd1 vssd1 vccd1 vccd1 net2644 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11850_ _05846_ _05913_ vssd1 vssd1 vccd1 vccd1 _05929_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_142_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06758__A2_N net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10439__C1 net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10801_ _05559_ _05560_ vssd1 vssd1 vccd1 vccd1 _05561_ sky130_fd_sc_hd__nor2_1
X_11781_ button\[0\] button\[2\] button\[1\] vssd1 vssd1 vccd1 vccd1 _05895_ sky130_fd_sc_hd__or3b_1
XANTENNA__11452__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13520_ clknet_leaf_24_clk _00330_ net1156 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[25\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10732_ net1572 net568 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[18\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_45_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13451_ clknet_leaf_56_clk _00261_ net1161 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10663_ _05443_ _05445_ vssd1 vssd1 vccd1 vccd1 _05482_ sky130_fd_sc_hd__nand2_1
XANTENNA__08046__B net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12402_ net1380 net131 _06348_ vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__a21o_1
XFILLER_127_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13382_ clknet_leaf_29_clk _00192_ net1133 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10594_ _05405_ _05416_ net615 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.zero_multi
+ sky130_fd_sc_hd__a21oi_2
XFILLER_127_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12333_ net640 _04833_ vssd1 vssd1 vccd1 vccd1 _06304_ sky130_fd_sc_hd__or2_1
XFILLER_5_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10592__A _02439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08280__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09158__A _02217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06830__A1 _01505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12264_ net229 net306 vssd1 vssd1 vccd1 vccd1 _06254_ sky130_fd_sc_hd__nand2_4
XFILLER_99_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06830__B2 datapath.ru.latched_instruction\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_147_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14003_ clknet_leaf_112_clk _00780_ net1198 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08032__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11215_ net284 net2285 net528 vssd1 vssd1 vccd1 vccd1 _00265_ sky130_fd_sc_hd__mux2_1
X_12195_ net2638 _06205_ _06207_ vssd1 vssd1 vccd1 vccd1 _00759_ sky130_fd_sc_hd__o21a_1
Xoutput50 net50 vssd1 vssd1 vccd1 vccd1 ADR_O[19] sky130_fd_sc_hd__buf_2
Xoutput61 net61 vssd1 vssd1 vccd1 vccd1 ADR_O[29] sky130_fd_sc_hd__buf_2
XFILLER_150_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07386__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 CYC_O sky130_fd_sc_hd__buf_2
Xoutput83 net83 vssd1 vssd1 vccd1 vccd1 DAT_O[19] sky130_fd_sc_hd__buf_2
X_11146_ net296 net2437 net531 vssd1 vssd1 vccd1 vccd1 _00199_ sky130_fd_sc_hd__mux2_1
Xoutput94 net94 vssd1 vssd1 vccd1 vccd1 DAT_O[29] sky130_fd_sc_hd__buf_2
XANTENNA__10390__A1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11077_ net299 net2182 net534 vssd1 vssd1 vccd1 vccd1 _00134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07138__A2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08335__A1 _03170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10028_ _04860_ _04861_ _04863_ vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__nand3_2
XANTENNA__09532__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07125__B net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11979_ _05741_ _05831_ vssd1 vssd1 vccd1 vccd1 _06024_ sky130_fd_sc_hd__and2_1
XANTENNA__06964__B net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11362__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13718_ clknet_leaf_141_clk _00528_ net1095 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14698_ clknet_leaf_60_clk _01403_ net1167 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07310__A2 _02145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13649_ clknet_leaf_39_clk _00459_ net1141 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07170_ datapath.rf.registers\[29\]\[27\] net975 net917 vssd1 vssd1 vccd1 vccd1 _02006_
+ sky130_fd_sc_hd__and3_1
XANTENNA__06980__A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08271__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_120_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_120_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_113_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08403__C net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08023__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12921__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout306 net307 vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__buf_4
XANTENNA__07377__A2 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09771__B1 _03978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout317 _03699_ vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__buf_2
X_09811_ net631 _04646_ vssd1 vssd1 vccd1 vccd1 _04647_ sky130_fd_sc_hd__and2_1
Xfanout328 _03622_ vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__buf_2
Xfanout339 _03683_ vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__clkbuf_2
XFILLER_101_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkload11_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10381__B2 _03673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09742_ net906 _03530_ _04575_ _04576_ _04577_ vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__a2111o_1
X_06954_ _01788_ net913 vssd1 vssd1 vccd1 vccd1 _01790_ sky130_fd_sc_hd__and2_1
XANTENNA__07129__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09673_ _02961_ _02983_ _03722_ vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__a21oi_1
X_06885_ net984 _01720_ vssd1 vssd1 vccd1 vccd1 _01721_ sky130_fd_sc_hd__and2_2
XFILLER_55_746 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07035__B net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08624_ _02285_ _03454_ _03457_ _02287_ vssd1 vssd1 vccd1 vccd1 _03460_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_38_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08555_ datapath.rf.registers\[22\]\[0\] net963 net909 _01809_ vssd1 vssd1 vccd1
+ vccd1 _03391_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout441_A net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09826__A1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1183_A net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11272__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout539_A net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07506_ datapath.rf.registers\[22\]\[20\] net954 net922 vssd1 vssd1 vccd1 vccd1 _02342_
+ sky130_fd_sc_hd__and3_1
X_08486_ _01591_ net897 _01665_ vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07301__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07437_ datapath.rf.registers\[11\]\[22\] net710 _02272_ net786 vssd1 vssd1 vccd1
+ vccd1 _02273_ sky130_fd_sc_hd__a211o_1
XFILLER_11_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout706_A net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06890__A net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07368_ datapath.rf.registers\[8\]\[23\] net876 net829 datapath.rf.registers\[14\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__a22o_1
XFILLER_108_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09107_ _03941_ _03942_ _03684_ vssd1 vssd1 vccd1 vccd1 _03943_ sky130_fd_sc_hd__mux2_1
XANTENNA__08262__B1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_111_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_111_clk
+ sky130_fd_sc_hd__clkbuf_8
X_07299_ datapath.rf.registers\[19\]\[25\] net732 net670 datapath.rf.registers\[21\]\[25\]
+ _02134_ vssd1 vssd1 vccd1 vccd1 _02135_ sky130_fd_sc_hd__a221o_1
X_09038_ _03873_ vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__inv_2
XFILLER_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout696_X net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold360 datapath.rf.registers\[15\]\[4\] vssd1 vssd1 vccd1 vccd1 net1708 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12831__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold371 datapath.rf.registers\[19\]\[23\] vssd1 vssd1 vccd1 vccd1 net1719 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06889__X _01725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07368__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold382 datapath.rf.registers\[16\]\[20\] vssd1 vssd1 vccd1 vccd1 net1730 sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 datapath.rf.registers\[21\]\[14\] vssd1 vssd1 vccd1 vccd1 net1741 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ net1699 net171 net434 vssd1 vssd1 vccd1 vccd1 _00065_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout863_X net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11447__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout840 _01740_ vssd1 vssd1 vccd1 vccd1 net840 sky130_fd_sc_hd__buf_6
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout851 _01735_ vssd1 vssd1 vccd1 vccd1 net851 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_144_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout862 net863 vssd1 vssd1 vccd1 vccd1 net862 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_144_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout873 _01723_ vssd1 vssd1 vccd1 vccd1 net873 sky130_fd_sc_hd__buf_2
Xfanout884 _01719_ vssd1 vssd1 vccd1 vccd1 net884 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09514__B1 _02750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout895 net896 vssd1 vssd1 vccd1 vccd1 net895 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06768__C _01604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12951_ net210 net2457 net394 vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__mux2_1
Xhold1060 datapath.rf.registers\[14\]\[22\] vssd1 vssd1 vccd1 vccd1 net2408 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1071 datapath.rf.registers\[19\]\[9\] vssd1 vssd1 vccd1 vccd1 net2419 sky130_fd_sc_hd__dlygate4sd3_1
X_11902_ net2523 net161 vssd1 vssd1 vccd1 vccd1 _05965_ sky130_fd_sc_hd__nand2_1
XFILLER_46_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1082 datapath.mulitply_result\[10\] vssd1 vssd1 vccd1 vccd1 net2430 sky130_fd_sc_hd__dlygate4sd3_1
X_12882_ net237 net2375 net400 vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__mux2_1
Xhold1093 datapath.rf.registers\[4\]\[10\] vssd1 vssd1 vccd1 vccd1 net2441 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_47_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07540__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14621_ clknet_leaf_146_clk _01326_ net1064 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11833_ _05303_ net1001 _05819_ _05911_ vssd1 vssd1 vccd1 vccd1 _05912_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_16_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09278__C1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06784__B net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11182__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07828__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14552_ clknet_leaf_6_clk _01257_ net1068 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11764_ net1470 net143 net138 _02189_ vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__a22o_1
XFILLER_14_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13503_ clknet_leaf_14_clk _00313_ net1079 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10715_ net2497 net573 vssd1 vssd1 vccd1 vccd1 _05510_ sky130_fd_sc_hd__nor2_1
X_14483_ clknet_leaf_39_clk _01188_ net1142 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11695_ _05019_ net155 net148 net1430 vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__a22o_1
XFILLER_146_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13434_ clknet_leaf_2_clk _00244_ net1065 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10646_ _05439_ _05440_ vssd1 vssd1 vccd1 vccd1 _05466_ sky130_fd_sc_hd__nor2_1
XFILLER_127_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13365_ clknet_leaf_129_clk _00175_ net1117 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10577_ _02025_ _02069_ _02125_ _02169_ vssd1 vssd1 vccd1 vccd1 _05400_ sky130_fd_sc_hd__or4_1
X_12316_ net635 _04867_ vssd1 vssd1 vccd1 vccd1 _06292_ sky130_fd_sc_hd__nor2_1
X_13296_ clknet_leaf_25_clk _00106_ net1159 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_114_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12247_ net1520 _06238_ _06240_ vssd1 vssd1 vccd1 vccd1 _00778_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12741__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_39_Left_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09616__A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12178_ _06197_ _06196_ net1270 vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__mux2_1
XFILLER_69_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11357__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06959__B net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11129_ net213 net1602 net426 vssd1 vssd1 vccd1 vccd1 _00184_ sky130_fd_sc_hd__mux2_1
XANTENNA__12104__A2 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06670_ _01492_ _01501_ _01508_ _01499_ vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__or4b_1
XANTENNA__06975__A _01797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07531__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07022__A_N net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_106_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06694__B net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11092__S net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07819__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08340_ datapath.rf.registers\[10\]\[3\] net986 net937 vssd1 vssd1 vccd1 vccd1 _03176_
+ sky130_fd_sc_hd__and3_1
X_08271_ datapath.rf.registers\[12\]\[5\] net755 net695 datapath.rf.registers\[8\]\[5\]
+ _03105_ vssd1 vssd1 vccd1 vccd1 _03107_ sky130_fd_sc_hd__a221o_1
XANTENNA__10784__X _05547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12916__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07222_ _02051_ _02053_ _02055_ _02057_ vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__or4_1
X_07153_ datapath.rf.registers\[26\]\[28\] net780 net678 datapath.rf.registers\[29\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_95_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08795__A1 _03419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12591__A2 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07084_ _01916_ _01917_ _01919_ vssd1 vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__nor3_1
XFILLER_154_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1029_A net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout391_A net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout136 _05934_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__buf_2
XANTENNA__11267__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout147 _05886_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__clkbuf_4
XFILLER_101_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout489_A _06552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout158 net159 vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__buf_2
XFILLER_87_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout169 net171 vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__clkbuf_2
X_07986_ datapath.rf.registers\[14\]\[11\] net776 net768 datapath.rf.registers\[24\]\[11\]
+ _02821_ vssd1 vssd1 vccd1 vccd1 _02822_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_126_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07770__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09725_ _04540_ _04560_ _04558_ vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__a21o_1
XFILLER_68_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06937_ net977 net917 vssd1 vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout656_A net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11854__A1 _05281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09656_ _03604_ _04491_ _04490_ net616 vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_2_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06885__A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06868_ _01703_ vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__inv_2
XFILLER_27_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07333__X _02169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08607_ _02727_ _02750_ _02772_ _03441_ vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__o31a_1
X_09587_ net326 _04072_ vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__or2_1
X_06799_ net1002 net1018 _01634_ vssd1 vssd1 vccd1 vccd1 _01635_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1186_X net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08538_ datapath.rf.registers\[1\]\[0\] net848 net828 datapath.rf.registers\[12\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__a22o_1
XANTENNA__12826__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08469_ datapath.rf.registers\[17\]\[1\] net852 net838 datapath.rf.registers\[26\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03305_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout611_X net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout709_X net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10500_ _05323_ _05328_ vssd1 vssd1 vccd1 vccd1 _05330_ sky130_fd_sc_hd__nand2b_1
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11480_ net288 net2275 net513 vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__mux2_1
XANTENNA__08605__A _02704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08235__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10431_ net631 _05243_ _05245_ _05266_ vssd1 vssd1 vccd1 vccd1 _05267_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_137_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_154_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07589__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13150_ net2025 net212 net383 vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__mux2_1
XFILLER_152_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout980_X net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10362_ net222 _05197_ net1292 vssd1 vssd1 vccd1 vccd1 _05198_ sky130_fd_sc_hd__a21o_1
XFILLER_128_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12101_ _06136_ _06138_ net1001 vssd1 vssd1 vccd1 vccd1 _06139_ sky130_fd_sc_hd__o21a_1
XFILLER_151_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13081_ net2443 net238 net388 vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__mux2_1
X_10293_ datapath.PC\[5\] _03733_ vssd1 vssd1 vccd1 vccd1 _05129_ sky130_fd_sc_hd__nand2_1
XFILLER_2_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12334__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12032_ _05343_ net998 _05824_ _05335_ _06073_ vssd1 vssd1 vccd1 vccd1 _06074_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_57_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09735__B1 _03770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold190 datapath.rf.registers\[0\]\[27\] vssd1 vssd1 vccd1 vccd1 net1538 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06779__B net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11177__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout670 _01832_ vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__buf_4
XANTENNA__07761__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout681 _01828_ vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__clkbuf_8
Xfanout692 _01824_ vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13983_ clknet_leaf_108_clk _00760_ net1221 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_18_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12934_ net294 net2005 net394 vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__mux2_1
XANTENNA__11845__B2 _05335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12865_ net286 net2355 net401 vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__mux2_1
X_14604_ clknet_leaf_133_clk _01309_ net1111 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11816_ net1047 net1015 net314 net334 datapath.ru.latched_instruction\[22\] vssd1
+ vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__a32o_1
X_12796_ _05515_ _05694_ vssd1 vssd1 vccd1 vccd1 _06551_ sky130_fd_sc_hd__nor2_4
X_14535_ clknet_leaf_144_clk _01240_ net1086 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11747_ net1461 net143 net138 _03028_ vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__a22o_1
XANTENNA__07122__C net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08474__B1 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12736__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09671__C1 _03614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14466_ clknet_leaf_150_clk _01171_ net1053 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11678_ _05126_ net154 net150 net1397 vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__a22o_1
X_13417_ clknet_leaf_21_clk _00227_ net1163 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10629_ net1037 _05447_ vssd1 vssd1 vccd1 vccd1 _05449_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_40_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14397_ clknet_leaf_144_clk _01102_ net1085 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_77_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12573__A2 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_47_Left_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13348_ clknet_leaf_18_clk _00158_ net1109 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11876__A _03076_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13279_ clknet_leaf_13_clk _00089_ net1078 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10336__A1 _04272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11087__S net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07840_ datapath.rf.registers\[22\]\[14\] net735 net669 datapath.rf.registers\[21\]\[14\]
+ _02675_ vssd1 vssd1 vccd1 vccd1 _02676_ sky130_fd_sc_hd__a221o_1
XANTENNA__07752__A2 _02587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07771_ datapath.rf.registers\[2\]\[15\] net888 net886 datapath.rf.registers\[9\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02607_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09510_ _03205_ net554 net550 vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__or3_1
X_06722_ _01554_ _01555_ _01556_ _01560_ vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__or4b_1
XPHY_EDGE_ROW_56_Left_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09441_ net349 _04188_ _04189_ vssd1 vssd1 vccd1 vccd1 _04277_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_88_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06653_ datapath.ru.latched_instruction\[12\] _01481_ _01489_ _01491_ vssd1 vssd1
+ vccd1 vccd1 _01492_ sky130_fd_sc_hd__a211o_1
XFILLER_24_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_121_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08409__B net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07313__B net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09372_ _03445_ _03524_ vssd1 vssd1 vccd1 vccd1 _04208_ sky130_fd_sc_hd__xnor2_1
X_06584_ screen.counter.ct\[16\] vssd1 vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__inv_2
XANTENNA__06992__X _01828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08323_ datapath.rf.registers\[11\]\[4\] net710 net699 datapath.rf.registers\[23\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03159_ sky130_fd_sc_hd__a22o_1
XANTENNA__08465__B1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout237_A _05616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10811__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08254_ datapath.rf.registers\[6\]\[5\] net825 net822 datapath.rf.registers\[22\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03090_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07205_ datapath.rf.registers\[10\]\[27\] net707 _02038_ _02040_ net787 vssd1 vssd1
+ vccd1 vccd1 _02041_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__08217__B1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_04_1301 vssd1 vssd1 vccd1 vccd1 team_04_1301/HI gpio_oeb[10] sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_65_Left_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08185_ datapath.rf.registers\[10\]\[7\] net708 net662 datapath.rf.registers\[5\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__a22o_1
Xteam_04_1312 vssd1 vssd1 vccd1 vccd1 team_04_1312/HI gpio_out[5] sky130_fd_sc_hd__conb_1
XANTENNA_fanout404_A _06549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xteam_04_1323 vssd1 vssd1 vccd1 vccd1 team_04_1323/HI gpio_out[27] sky130_fd_sc_hd__conb_1
Xteam_04_1334 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] team_04_1334/LO sky130_fd_sc_hd__conb_1
XFILLER_146_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07136_ datapath.rf.registers\[8\]\[28\] net878 net809 datapath.rf.registers\[27\]\[28\]
+ _01971_ vssd1 vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__a221o_1
Xteam_04_1345 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] team_04_1345/LO sky130_fd_sc_hd__conb_1
XANTENNA__11786__A net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07067_ datapath.rf.registers\[17\]\[30\] net748 net670 datapath.rf.registers\[21\]\[30\]
+ _01902_ vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__a221o_1
XANTENNA__10327__A1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout394_X net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10878__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07743__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout940_A _01717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_74_Left_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07969_ datapath.rf.registers\[0\]\[11\] net869 _02803_ vssd1 vssd1 vccd1 vccd1 _02805_
+ sky130_fd_sc_hd__o21ai_4
X_09708_ _03663_ _04541_ _04543_ net650 vssd1 vssd1 vccd1 vccd1 _04544_ sky130_fd_sc_hd__o211a_1
X_10980_ net2412 net266 net436 vssd1 vssd1 vccd1 vccd1 _00045_ sky130_fd_sc_hd__mux2_1
XFILLER_43_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09639_ _04396_ _04428_ _04454_ _04474_ vssd1 vssd1 vccd1 vccd1 _04475_ sky130_fd_sc_hd__or4b_1
XANTENNA_fanout826_X net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12650_ _06481_ _06485_ _06488_ vssd1 vssd1 vccd1 vccd1 _06489_ sky130_fd_sc_hd__a21o_1
XANTENNA__07223__B net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11601_ net997 _05824_ vssd1 vssd1 vccd1 vccd1 _05825_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_139_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12581_ datapath.mulitply_result\[12\] datapath.multiplication_module.multiplicand_i\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06431_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_156_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11460__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14320_ clknet_leaf_23_clk _01025_ net1155 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[23\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11532_ _01422_ screen.counter.ct\[5\] _05301_ vssd1 vssd1 vccd1 vccd1 _05756_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_83_Left_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10584__B _02876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14251_ clknet_leaf_55_clk _00956_ net1174 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_152_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11463_ net2258 net238 net408 vssd1 vssd1 vccd1 vccd1 _00501_ sky130_fd_sc_hd__mux2_1
XFILLER_7_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08054__B net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13202_ clknet_leaf_30_clk _00012_ net1132 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10414_ _03262_ _03657_ vssd1 vssd1 vccd1 vccd1 _05250_ sky130_fd_sc_hd__nand2_1
XANTENNA__12555__A2 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14182_ clknet_leaf_51_clk _00937_ net1182 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_124_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11394_ net1537 net240 net412 vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__mux2_1
X_13133_ net1740 net296 net382 vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__mux2_1
X_10345_ net1267 _03736_ datapath.PC\[10\] vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07893__B net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07982__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ net1686 net288 net388 vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__mux2_1
X_10276_ net892 _05107_ _05111_ net227 vssd1 vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12015_ net1007 _05758_ vssd1 vssd1 vccd1 vccd1 _06058_ sky130_fd_sc_hd__nor2_1
XANTENNA__08501__C _01816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07195__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07734__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11818__A1 datapath.ru.latched_instruction\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13966_ clknet_leaf_106_clk _00744_ net1223 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_62_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12917_ net2471 net214 net482 vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__mux2_1
XANTENNA__11207__Y _05721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13897_ clknet_leaf_44_clk keypad.decode.sticky_n\[2\] net1151 vssd1 vssd1 vccd1
+ vccd1 keypad.decode.sticky\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12848_ net219 net2269 net486 vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__mux2_1
XFILLER_62_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12779_ net247 net1948 net495 vssd1 vssd1 vccd1 vccd1 _01032_ sky130_fd_sc_hd__mux2_1
XANTENNA__11370__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06972__B net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08998__A1 _01934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14518_ clknet_leaf_142_clk _01223_ net1093 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08245__A net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14449_ clknet_leaf_35_clk _01154_ net1129 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_128_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold904 datapath.rf.registers\[10\]\[15\] vssd1 vssd1 vccd1 vccd1 net2252 sky130_fd_sc_hd__dlygate4sd3_1
Xhold915 datapath.rf.registers\[2\]\[24\] vssd1 vssd1 vccd1 vccd1 net2263 sky130_fd_sc_hd__dlygate4sd3_1
Xhold926 datapath.rf.registers\[23\]\[11\] vssd1 vssd1 vccd1 vccd1 net2274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold937 datapath.rf.registers\[18\]\[7\] vssd1 vssd1 vccd1 vccd1 net2285 sky130_fd_sc_hd__dlygate4sd3_1
Xhold948 datapath.rf.registers\[24\]\[29\] vssd1 vssd1 vccd1 vccd1 net2296 sky130_fd_sc_hd__dlygate4sd3_1
X_09990_ _04720_ _04825_ vssd1 vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__nand2_1
Xhold959 datapath.rf.registers\[22\]\[12\] vssd1 vssd1 vccd1 vccd1 net2307 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10714__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07973__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08941_ net347 _03776_ vssd1 vssd1 vccd1 vccd1 _03777_ sky130_fd_sc_hd__or2_1
XANTENNA__10309__A1 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08411__C net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08872_ _03009_ net560 net446 vssd1 vssd1 vccd1 vccd1 _03708_ sky130_fd_sc_hd__mux2_1
XANTENNA__07186__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06987__X _01823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07725__A2 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07823_ _02646_ _02654_ _02656_ _02658_ vssd1 vssd1 vccd1 vccd1 _02659_ sky130_fd_sc_hd__or4_1
XANTENNA__07027__C net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07754_ net561 _02588_ vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__nor2_1
XANTENNA__11809__B2 datapath.ru.latched_instruction\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_65_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06705_ datapath.ru.latched_instruction\[24\] datapath.ru.latched_instruction\[25\]
+ datapath.ru.latched_instruction\[26\] datapath.ru.latched_instruction\[27\] vssd1
+ vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__or4_1
X_07685_ _02513_ _02518_ _02520_ vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__or3_4
XFILLER_52_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_91_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_91_clk sky130_fd_sc_hd__clkbuf_8
X_09424_ _04125_ _04259_ net374 vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__mux2_1
X_06636_ net1288 net1283 mmio.memload_or_instruction\[11\] vssd1 vssd1 vccd1 vccd1
+ _01475_ sky130_fd_sc_hd__or3b_1
XFILLER_80_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09355_ _03965_ _03966_ net359 vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__a21o_1
X_06567_ datapath.ru.latched_instruction\[0\] vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout142_X net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11280__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06882__B _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08306_ _03139_ _03140_ _03141_ vssd1 vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__or3_1
XFILLER_139_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09286_ _03578_ _04119_ _04121_ vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07110__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_7_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08237_ datapath.rf.registers\[30\]\[6\] net758 net702 datapath.rf.registers\[9\]\[6\]
+ _03067_ vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__a221o_1
XFILLER_154_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1051_X net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout407_X net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08168_ datapath.rf.registers\[24\]\[7\] net858 net820 datapath.rf.registers\[5\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03004_ sky130_fd_sc_hd__a22o_1
XFILLER_107_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout890_A net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout988_A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07119_ net614 _01954_ net565 vssd1 vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__a21oi_1
X_08099_ _01594_ _01784_ vssd1 vssd1 vccd1 vccd1 _02935_ sky130_fd_sc_hd__nor2_1
XANTENNA__13000__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10130_ _04933_ _04943_ _04965_ _04932_ vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__a211o_1
XFILLER_122_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout776_X net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09166__A1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10061_ _04895_ _04896_ vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__nand2b_1
XANTENNA__07218__B net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07177__B1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07716__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_149_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout943_X net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10720__A1 _03057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11455__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13820_ clknet_leaf_98_clk _00629_ net1230 vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10579__B net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07234__A _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13751_ clknet_leaf_88_clk _00560_ net1253 vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__dfrtp_1
X_10963_ net1525 net208 net437 vssd1 vssd1 vccd1 vccd1 _00034_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_82_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08049__B net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12702_ columns.count\[0\] _06531_ vssd1 vssd1 vccd1 vccd1 _06532_ sky130_fd_sc_hd__nand2_1
XFILLER_44_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08141__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13682_ clknet_leaf_33_clk _00492_ net1125 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10894_ _01527_ net654 _05640_ vssd1 vssd1 vccd1 vccd1 _05641_ sky130_fd_sc_hd__o21a_4
XFILLER_44_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12633_ _06466_ _06473_ _06472_ _06471_ vssd1 vssd1 vccd1 vccd1 _06475_ sky130_fd_sc_hd__o211ai_1
XFILLER_31_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11190__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12564_ datapath.mulitply_result\[9\] datapath.multiplication_module.multiplicand_i\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06417_ sky130_fd_sc_hd__and2_1
XANTENNA__07101__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08065__A net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11984__B1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14303_ clknet_leaf_16_clk _01008_ net1106 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_11515_ _05338_ _05340_ _05347_ vssd1 vssd1 vccd1 vccd1 _05740_ sky130_fd_sc_hd__and3_1
XANTENNA__14014__RESET_B net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07652__A1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12495_ net241 net1862 net507 vssd1 vssd1 vccd1 vccd1 _00895_ sky130_fd_sc_hd__mux2_1
XFILLER_8_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14234_ clknet_leaf_123_clk datapath.multiplication_module.multiplier_i_n\[2\] net1215
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i\[2\] sky130_fd_sc_hd__dfrtp_1
X_11446_ net1668 net289 net409 vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__mux2_1
XFILLER_137_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07404__A1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14165_ clknet_leaf_70_clk _00920_ net1244 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11377_ net1829 net209 net413 vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__mux2_1
X_13116_ net214 net2499 net470 vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__mux2_1
XANTENNA__07955__A2 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10328_ _04860_ _04861_ _04863_ vssd1 vssd1 vccd1 vccd1 _05164_ sky130_fd_sc_hd__a21o_1
XFILLER_3_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14096_ clknet_leaf_122_clk _00862_ net1201 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13047_ net220 net1914 net475 vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__mux2_1
X_10259_ datapath.PC\[11\] net1249 _05091_ _05094_ vssd1 vssd1 vccd1 vccd1 _05095_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07707__A2 _02542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1240 net1241 vssd1 vssd1 vccd1 vccd1 net1240 sky130_fd_sc_hd__clkbuf_2
Xfanout1251 net1261 vssd1 vssd1 vccd1 vccd1 net1251 sky130_fd_sc_hd__buf_2
XANTENNA__11873__B net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1262 _00004_ vssd1 vssd1 vccd1 vccd1 net1262 sky130_fd_sc_hd__buf_4
Xfanout1273 screen.counter.ct\[13\] vssd1 vssd1 vccd1 vccd1 net1273 sky130_fd_sc_hd__clkbuf_2
XFILLER_94_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11365__S net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1284 net1285 vssd1 vssd1 vccd1 vccd1 net1284 sky130_fd_sc_hd__buf_1
Xfanout1295 _01436_ vssd1 vssd1 vccd1 vccd1 net1295 sky130_fd_sc_hd__clkbuf_2
XFILLER_94_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10489__B _05314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13949_ clknet_leaf_103_clk _00727_ net1225 vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_85_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_73_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08132__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_866 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07470_ _02303_ _02304_ _02305_ vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__or3_1
XFILLER_50_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06983__A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07340__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10227__B1 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09140_ _03970_ _03972_ _03975_ vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__or3b_1
XANTENNA__09093__A0 _02126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09071_ net451 _03712_ vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__or2_1
XANTENNA__12924__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10792__X _05554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08022_ datapath.rf.registers\[27\]\[10\] net685 net673 datapath.rf.registers\[7\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_116_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold701 datapath.rf.registers\[24\]\[15\] vssd1 vssd1 vccd1 vccd1 net2049 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08703__A _02961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold712 datapath.rf.registers\[23\]\[4\] vssd1 vssd1 vccd1 vccd1 net2060 sky130_fd_sc_hd__dlygate4sd3_1
Xhold723 datapath.rf.registers\[13\]\[26\] vssd1 vssd1 vccd1 vccd1 net2071 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold734 datapath.rf.registers\[12\]\[15\] vssd1 vssd1 vccd1 vccd1 net2082 sky130_fd_sc_hd__dlygate4sd3_1
Xhold745 datapath.rf.registers\[22\]\[14\] vssd1 vssd1 vccd1 vccd1 net2093 sky130_fd_sc_hd__dlygate4sd3_1
Xhold756 datapath.rf.registers\[13\]\[10\] vssd1 vssd1 vccd1 vccd1 net2104 sky130_fd_sc_hd__dlygate4sd3_1
Xhold767 datapath.rf.registers\[1\]\[23\] vssd1 vssd1 vccd1 vccd1 net2115 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold778 datapath.rf.registers\[25\]\[24\] vssd1 vssd1 vccd1 vccd1 net2126 sky130_fd_sc_hd__dlygate4sd3_1
X_09973_ _04740_ _04743_ _04807_ _04739_ vssd1 vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__a31o_1
Xhold789 datapath.rf.registers\[10\]\[31\] vssd1 vssd1 vccd1 vccd1 net2137 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08924_ net557 net577 _03759_ vssd1 vssd1 vccd1 vccd1 _03760_ sky130_fd_sc_hd__o21a_1
XANTENNA__07159__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1109_A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08855_ _02523_ net561 net444 vssd1 vssd1 vccd1 vccd1 _03691_ sky130_fd_sc_hd__mux2_1
XANTENNA__10702__A1 _03028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout471_A net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06906__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout569_A _05368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11275__S net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06877__B net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07806_ datapath.rf.registers\[9\]\[14\] net885 net811 datapath.rf.registers\[13\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02642_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08786_ _01647_ _03229_ _03615_ vssd1 vssd1 vccd1 vccd1 _03622_ sky130_fd_sc_hd__mux2_1
XFILLER_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07737_ datapath.rf.registers\[27\]\[16\] net683 net668 datapath.rf.registers\[21\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout736_A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_64_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_41_803 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07668_ datapath.rf.registers\[22\]\[17\] net952 net925 vssd1 vssd1 vccd1 vccd1 _02504_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07331__B1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09407_ _03572_ _04240_ _04242_ vssd1 vssd1 vccd1 vccd1 _04243_ sky130_fd_sc_hd__a21o_1
X_06619_ datapath.ru.latched_instruction\[4\] _01449_ _01455_ _01457_ _01447_ vssd1
+ vssd1 vccd1 vccd1 _01458_ sky130_fd_sc_hd__a2111o_1
XFILLER_41_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout524_X net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07599_ datapath.rf.registers\[30\]\[19\] net760 net752 datapath.rf.registers\[28\]\[19\]
+ _02433_ vssd1 vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__a221o_1
XFILLER_111_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07501__B net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09084__A0 _02125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09338_ net319 net317 _03942_ _04169_ _04173_ vssd1 vssd1 vccd1 vccd1 _04174_ sky130_fd_sc_hd__o311a_1
XANTENNA__10769__A1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08316__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09269_ _03963_ _03964_ net355 vssd1 vssd1 vccd1 vccd1 _04105_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12834__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11300_ net192 net2567 net522 vssd1 vssd1 vccd1 vccd1 _00348_ sky130_fd_sc_hd__mux2_1
XANTENNA__08172__X _03008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12280_ net892 _04845_ vssd1 vssd1 vccd1 vccd1 _06266_ sky130_fd_sc_hd__nand2_1
XFILLER_107_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11231_ net205 net2031 net526 vssd1 vssd1 vccd1 vccd1 _00281_ sky130_fd_sc_hd__mux2_1
XANTENNA__12135__A _06168_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07398__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11162_ net216 net1874 net530 vssd1 vssd1 vccd1 vccd1 _00215_ sky130_fd_sc_hd__mux2_1
XANTENNA__10792__A1_N _01467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09139__A1 _01620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08051__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10113_ _04118_ _04601_ vssd1 vssd1 vccd1 vccd1 _04949_ sky130_fd_sc_hd__xnor2_1
XFILLER_49_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11093_ net231 net1592 net535 vssd1 vssd1 vccd1 vccd1 _00150_ sky130_fd_sc_hd__mux2_1
XFILLER_103_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input32_A DAT_I[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10044_ _04819_ _04879_ vssd1 vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__xnor2_1
Xhold50 screen.controlBus\[18\] vssd1 vssd1 vccd1 vccd1 net1398 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11185__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold61 net65 vssd1 vssd1 vccd1 vccd1 net1409 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08362__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold72 net43 vssd1 vssd1 vccd1 vccd1 net1420 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 net115 vssd1 vssd1 vccd1 vccd1 net1431 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 net118 vssd1 vssd1 vccd1 vccd1 net1442 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07570__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13803_ clknet_leaf_75_clk _00612_ net1242 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[24\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_91_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10877__X _05626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11995_ _05330_ _05795_ _05842_ _06038_ vssd1 vssd1 vccd1 vccd1 _06039_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_67_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_55_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08114__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13734_ clknet_leaf_23_clk _00544_ net1154 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_11_Left_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10946_ datapath.PC\[31\] _05678_ vssd1 vssd1 vccd1 vccd1 _05685_ sky130_fd_sc_hd__xor2_1
XFILLER_17_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07322__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13665_ clknet_leaf_46_clk _00475_ net1172 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10877_ net898 _04057_ _05625_ net600 vssd1 vssd1 vccd1 vccd1 _05626_ sky130_fd_sc_hd__a211o_2
XANTENNA__08507__B net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12616_ net498 _06459_ _06460_ net502 net2509 vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_80_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07411__B net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13596_ clknet_leaf_8_clk _00406_ net1071 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12547_ _06395_ _06396_ _06397_ vssd1 vssd1 vccd1 vccd1 _06403_ sky130_fd_sc_hd__o21ba_1
XANTENNA__12744__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12478_ net208 net1565 net508 vssd1 vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__mux2_1
XANTENNA_3 _06551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14217_ clknet_leaf_50_clk datapath.multiplication_module.multiplicand_i_n\[28\]
+ net1182 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_144_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11429_ net237 net2526 net516 vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__mux2_1
XFILLER_6_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Left_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07389__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07928__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14148_ clknet_leaf_119_clk _00905_ net1191 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14079_ clknet_leaf_99_clk net1349 net1229 vssd1 vssd1 vccd1 vccd1 screen.register.cFill2
+ sky130_fd_sc_hd__dfrtp_1
X_06970_ _01800_ net907 vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__and2_1
XANTENNA__11095__S net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1070 net1075 vssd1 vssd1 vccd1 vccd1 net1070 sky130_fd_sc_hd__clkbuf_2
Xfanout1081 net1084 vssd1 vssd1 vccd1 vccd1 net1081 sky130_fd_sc_hd__clkbuf_2
X_08640_ _01957_ _02004_ _03470_ _03473_ _01910_ vssd1 vssd1 vccd1 vccd1 _03476_ sky130_fd_sc_hd__o311a_1
Xfanout1092 net1120 vssd1 vssd1 vccd1 vccd1 net1092 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07561__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08571_ datapath.rf.registers\[1\]\[0\] net764 net733 datapath.rf.registers\[19\]\[0\]
+ _03406_ vssd1 vssd1 vccd1 vccd1 _03407_ sky130_fd_sc_hd__a221o_1
XANTENNA__12919__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_46_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09302__A1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07522_ _02354_ _02355_ _02356_ _02357_ vssd1 vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__or4_1
XANTENNA__08510__C1 _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07453_ datapath.rf.registers\[9\]\[21\] net981 net943 vssd1 vssd1 vccd1 vccd1 _02289_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_33_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07384_ datapath.rf.registers\[12\]\[23\] net754 net702 datapath.rf.registers\[9\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_33_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09605__A2 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09123_ net379 _03958_ net312 vssd1 vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__o21ba_1
XFILLER_109_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07040__C net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09054_ net347 _03889_ vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__or2_1
XANTENNA__07092__A2 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08005_ datapath.rf.registers\[31\]\[10\] net976 net915 vssd1 vssd1 vccd1 vccd1 _02841_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09369__A1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold520 datapath.rf.registers\[14\]\[7\] vssd1 vssd1 vccd1 vccd1 net1868 sky130_fd_sc_hd__dlygate4sd3_1
Xhold531 datapath.rf.registers\[24\]\[23\] vssd1 vssd1 vccd1 vccd1 net1879 sky130_fd_sc_hd__dlygate4sd3_1
Xhold542 datapath.rf.registers\[3\]\[23\] vssd1 vssd1 vccd1 vccd1 net1890 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08152__B net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07919__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold553 datapath.rf.registers\[3\]\[30\] vssd1 vssd1 vccd1 vccd1 net1901 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold564 datapath.rf.registers\[10\]\[14\] vssd1 vssd1 vccd1 vccd1 net1912 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold575 datapath.rf.registers\[7\]\[6\] vssd1 vssd1 vccd1 vccd1 net1923 sky130_fd_sc_hd__dlygate4sd3_1
Xhold586 datapath.rf.registers\[23\]\[18\] vssd1 vssd1 vccd1 vccd1 net1934 sky130_fd_sc_hd__dlygate4sd3_1
Xhold597 datapath.rf.registers\[27\]\[31\] vssd1 vssd1 vccd1 vccd1 net1945 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout686_A _01827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09956_ _04774_ _04791_ _04772_ vssd1 vssd1 vccd1 vccd1 _04792_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06888__A _01707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08907_ datapath.PC\[17\] datapath.PC\[18\] _03742_ vssd1 vssd1 vccd1 vccd1 _03743_
+ sky130_fd_sc_hd__or3_1
XANTENNA__09264__A _02364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09887_ datapath.PC\[20\] datapath.PC\[21\] net596 vssd1 vssd1 vccd1 vccd1 _04723_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_129_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout474_X net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout853_A net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1220 datapath.rf.registers\[0\]\[11\] vssd1 vssd1 vccd1 vccd1 net2568 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1231 datapath.rf.registers\[26\]\[27\] vssd1 vssd1 vccd1 vccd1 net2579 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09541__A1 _02961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08838_ _03669_ _03672_ vssd1 vssd1 vccd1 vccd1 _03674_ sky130_fd_sc_hd__or2_1
Xhold1242 datapath.rf.registers\[28\]\[10\] vssd1 vssd1 vccd1 vccd1 net2590 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_142_Right_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1253 datapath.rf.registers\[0\]\[31\] vssd1 vssd1 vccd1 vccd1 net2601 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1264 datapath.mulitply_result\[26\] vssd1 vssd1 vccd1 vccd1 net2612 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1275 datapath.rf.registers\[25\]\[20\] vssd1 vssd1 vccd1 vccd1 net2623 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1286 datapath.rf.registers\[0\]\[16\] vssd1 vssd1 vccd1 vccd1 net2634 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1297 datapath.rf.registers\[2\]\[4\] vssd1 vssd1 vccd1 vccd1 net2645 sky130_fd_sc_hd__dlygate4sd3_1
X_08769_ _03602_ _03603_ vssd1 vssd1 vccd1 vccd1 _03605_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_142_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout739_X net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_37_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_8
X_10800_ net1267 _05548_ datapath.PC\[10\] vssd1 vssd1 vccd1 vccd1 _05560_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_49_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ net124 _05446_ _05894_ vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__mux2_1
XANTENNA__07304__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10731_ net1533 net569 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[17\]
+ sky130_fd_sc_hd__and2_1
XANTENNA_fanout906_X net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13450_ clknet_leaf_58_clk _00260_ net1168 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[18\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10662_ _05444_ _05474_ _05478_ _05480_ vssd1 vssd1 vccd1 vccd1 _05481_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_62_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12401_ _05958_ net158 vssd1 vssd1 vccd1 vccd1 _06348_ sky130_fd_sc_hd__nor2_1
XANTENNA__08046__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13381_ clknet_leaf_114_clk _00191_ net1190 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10593_ _05410_ _05413_ _05414_ _05415_ vssd1 vssd1 vccd1 vccd1 _05416_ sky130_fd_sc_hd__or4_2
XFILLER_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12332_ datapath.PC\[21\] _06303_ net306 vssd1 vssd1 vccd1 vccd1 _00800_ sky130_fd_sc_hd__mux2_1
XFILLER_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07083__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09439__A net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10592__B _02487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12263_ net224 net310 vssd1 vssd1 vccd1 vccd1 _06253_ sky130_fd_sc_hd__nor2_4
X_14002_ clknet_leaf_111_clk _00779_ net1198 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_107_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11214_ net291 net2024 net526 vssd1 vssd1 vccd1 vccd1 _00264_ sky130_fd_sc_hd__mux2_1
X_12194_ screen.counter.currentCt\[1\] _06205_ _06172_ vssd1 vssd1 vccd1 vccd1 _06207_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput40 net40 vssd1 vssd1 vccd1 vccd1 ADR_O[0] sky130_fd_sc_hd__buf_2
Xoutput51 net51 vssd1 vssd1 vccd1 vccd1 ADR_O[1] sky130_fd_sc_hd__buf_2
XANTENNA__08583__A2 _03417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput62 net62 vssd1 vssd1 vccd1 vccd1 ADR_O[2] sky130_fd_sc_hd__buf_2
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 DAT_O[0] sky130_fd_sc_hd__buf_2
X_11145_ net298 net1951 net530 vssd1 vssd1 vccd1 vccd1 _00198_ sky130_fd_sc_hd__mux2_1
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 DAT_O[1] sky130_fd_sc_hd__buf_2
XANTENNA__10812__S net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07791__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput95 net95 vssd1 vssd1 vccd1 vccd1 DAT_O[2] sky130_fd_sc_hd__buf_2
XFILLER_150_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_94_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11076_ net305 net2434 net536 vssd1 vssd1 vccd1 vccd1 _00133_ sky130_fd_sc_hd__mux2_1
XANTENNA__09532__A1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10027_ _04806_ _04862_ vssd1 vssd1 vccd1 vccd1 _04863_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10113__A _04118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07406__B _02240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07543__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07125__C net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12739__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_28_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_19_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11978_ screen.counter.ct\[8\] _05854_ _06020_ _06022_ vssd1 vssd1 vccd1 vccd1 _06023_
+ sky130_fd_sc_hd__o31a_1
XFILLER_16_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_152_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13717_ clknet_leaf_18_clk _00527_ net1116 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10929_ net176 net1908 net543 vssd1 vssd1 vccd1 vccd1 _00030_ sky130_fd_sc_hd__mux2_1
X_14697_ clknet_leaf_92_clk _01402_ net1232 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10850__A0 _04146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_32_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13648_ clknet_leaf_57_clk _00458_ net1160 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11879__A _03028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13579_ clknet_leaf_55_clk _00389_ net1173 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06980__B _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09349__A _02567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_47_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout307 _06247_ vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__clkbuf_4
X_09810_ _03475_ _03482_ vssd1 vssd1 vccd1 vccd1 _04646_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09771__A1 _03947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout318 _03699_ vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__buf_1
Xfanout329 _03622_ vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__buf_2
XFILLER_141_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10381__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09741_ _03527_ net629 net625 _03528_ net643 vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__a221o_1
X_06953_ net991 _01666_ vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__nor2_1
XFILLER_140_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14671__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08326__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_105_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07316__B net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09672_ net574 _04501_ _04502_ _04507_ vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__a22o_1
XANTENNA__06995__X _01831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06884_ _01630_ net961 _01639_ _01656_ vssd1 vssd1 vccd1 vccd1 _01720_ sky130_fd_sc_hd__and4bb_4
XANTENNA__07534__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09371__X _04207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08623_ _03454_ _03457_ vssd1 vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__nand2_1
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07035__C net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_19_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_38_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout267_A net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07603__Y _02439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08554_ datapath.rf.registers\[25\]\[0\] net965 net908 _01800_ vssd1 vssd1 vccd1
+ vccd1 _03390_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_124_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07505_ datapath.rf.registers\[21\]\[20\] net945 net922 vssd1 vssd1 vccd1 vccd1 _02341_
+ sky130_fd_sc_hd__and3_1
XFILLER_23_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08485_ net559 vssd1 vssd1 vccd1 vccd1 _03321_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout434_A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1176_A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09039__A0 _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07436_ datapath.rf.registers\[1\]\[22\] net762 net714 datapath.rf.registers\[4\]\[22\]
+ _02271_ vssd1 vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__a221o_1
XFILLER_149_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07367_ datapath.rf.registers\[16\]\[23\] net860 net810 datapath.rf.registers\[13\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout222_X net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13752__RESET_B net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06890__B net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09106_ net340 _03814_ vssd1 vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__or2_1
XFILLER_109_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07065__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07298_ datapath.rf.registers\[23\]\[25\] net700 net689 datapath.rf.registers\[31\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__a22o_1
X_09037_ net364 _03834_ _03872_ vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__o21ai_1
XFILLER_105_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold350 datapath.rf.registers\[6\]\[28\] vssd1 vssd1 vccd1 vccd1 net1698 sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 datapath.multiplication_module.multiplicand_i\[20\] vssd1 vssd1 vccd1 vccd1
+ net1709 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout970_A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout689_X net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold372 datapath.rf.registers\[9\]\[2\] vssd1 vssd1 vccd1 vccd1 net1720 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold383 datapath.rf.registers\[6\]\[1\] vssd1 vssd1 vccd1 vccd1 net1731 sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 datapath.rf.registers\[12\]\[16\] vssd1 vssd1 vccd1 vccd1 net1742 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07773__B1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout830 net831 vssd1 vssd1 vccd1 vccd1 net830 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10372__A2 net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout841 net844 vssd1 vssd1 vccd1 vccd1 net841 sky130_fd_sc_hd__clkbuf_8
Xfanout852 _01735_ vssd1 vssd1 vccd1 vccd1 net852 sky130_fd_sc_hd__clkbuf_4
X_09939_ datapath.PC\[4\] _03150_ vssd1 vssd1 vccd1 vccd1 _04775_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_144_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout856_X net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout863 _01728_ vssd1 vssd1 vccd1 vccd1 net863 sky130_fd_sc_hd__clkbuf_4
XFILLER_93_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout874 _01723_ vssd1 vssd1 vccd1 vccd1 net874 sky130_fd_sc_hd__buf_4
Xfanout885 net886 vssd1 vssd1 vccd1 vccd1 net885 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08317__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_13_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_13_0_clk sky130_fd_sc_hd__clkbuf_8
X_12950_ net214 net2496 net394 vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__mux2_1
Xfanout896 _01628_ vssd1 vssd1 vccd1 vccd1 net896 sky130_fd_sc_hd__buf_2
Xhold1050 datapath.rf.registers\[15\]\[14\] vssd1 vssd1 vccd1 vccd1 net2398 sky130_fd_sc_hd__dlygate4sd3_1
X_11901_ net135 _05964_ _05963_ vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__o21ai_1
Xhold1061 datapath.rf.registers\[14\]\[12\] vssd1 vssd1 vccd1 vccd1 net2409 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1072 datapath.rf.registers\[14\]\[27\] vssd1 vssd1 vccd1 vccd1 net2420 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09722__A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12881_ net220 net2029 net398 vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__mux2_1
Xhold1083 datapath.rf.registers\[25\]\[6\] vssd1 vssd1 vccd1 vccd1 net2431 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1094 mmio.memload_or_instruction\[5\] vssd1 vssd1 vccd1 vccd1 net2442 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11463__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11832_ _05302_ _05785_ _05794_ net1010 vssd1 vssd1 vccd1 vccd1 _05911_ sky130_fd_sc_hd__o211a_1
X_14620_ clknet_leaf_8_clk _01325_ net1071 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09278__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08338__A _03149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14551_ clknet_leaf_130_clk _01256_ net1113 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[4\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11763_ net1485 net145 net140 _02239_ vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__a22o_1
XANTENNA__08057__B _01712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13502_ clknet_leaf_147_clk _00312_ net1064 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[11\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10714_ net2364 _03204_ net573 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[3\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA__10832__B1 _05586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14482_ clknet_leaf_27_clk _01187_ net1132 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[3\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11694_ _05041_ net155 net148 net1414 vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__a22o_1
X_13433_ clknet_leaf_9_clk _00243_ net1072 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10645_ net1013 _05464_ vssd1 vssd1 vccd1 vccd1 _05465_ sky130_fd_sc_hd__nor2_1
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12585__B1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13364_ clknet_leaf_127_clk _00174_ net1211 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07056__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10576_ _05397_ _05398_ vssd1 vssd1 vccd1 vccd1 _05399_ sky130_fd_sc_hd__nand2_1
XFILLER_127_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12315_ datapath.PC\[16\] net307 _06291_ _04998_ vssd1 vssd1 vccd1 vccd1 _00795_
+ sky130_fd_sc_hd__o22a_1
X_13295_ clknet_leaf_28_clk _00105_ net1134 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[8\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12246_ screen.counter.currentCt\[20\] _06238_ net602 vssd1 vssd1 vccd1 vccd1 _06240_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__09202__B1 _02311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10348__C1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08801__A _03636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08556__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12177_ _06164_ net601 vssd1 vssd1 vccd1 vccd1 _06197_ sky130_fd_sc_hd__and2_1
XANTENNA__07764__B1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10363__A2 net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11128_ net216 net1987 net426 vssd1 vssd1 vccd1 vccd1 _00183_ sky130_fd_sc_hd__mux2_1
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08308__A2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11059_ net215 net2042 net430 vssd1 vssd1 vccd1 vccd1 _00119_ sky130_fd_sc_hd__mux2_1
XFILLER_37_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11373__S net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06975__B net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_103_Left_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10823__A0 _04272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08270_ datapath.rf.registers\[20\]\[5\] net719 net699 datapath.rf.registers\[23\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03106_ sky130_fd_sc_hd__a22o_1
XANTENNA__06991__A net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07295__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07221_ datapath.rf.registers\[2\]\[26\] net887 net885 datapath.rf.registers\[9\]\[26\]
+ _02056_ vssd1 vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__a221o_1
XFILLER_9_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07047__A2 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07152_ datapath.rf.registers\[24\]\[28\] net768 net696 datapath.rf.registers\[8\]\[28\]
+ _01987_ vssd1 vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__a221o_1
XANTENNA__12040__A2 _05778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12932__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07083_ datapath.rf.registers\[17\]\[29\] net850 _01918_ net872 vssd1 vssd1 vccd1
+ vccd1 _01919_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_8_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08711__A net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09744__A1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout126 net127 vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08430__B net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout137 _05934_ vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__clkbuf_2
Xfanout148 net150 vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__buf_2
Xfanout159 _06335_ vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__buf_2
X_07985_ datapath.rf.registers\[26\]\[11\] net780 net728 datapath.rf.registers\[25\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__a22o_1
XFILLER_75_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout384_A net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09724_ _04552_ _04556_ _04559_ net555 vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_126_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06936_ net982 net915 vssd1 vssd1 vccd1 vccd1 _01772_ sky130_fd_sc_hd__and2_2
XFILLER_86_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09655_ _03562_ _03563_ vssd1 vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__xor2_1
X_06867_ _01576_ _01588_ vssd1 vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__nor2_4
XFILLER_28_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1293_A _01436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08180__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06885__B _01720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11283__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout649_A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08606_ _02750_ _02772_ vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__nor2_1
X_09586_ _04416_ _04421_ net326 vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__o21ai_1
XFILLER_83_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06798_ datapath.ru.latched_instruction\[22\] _01456_ net1014 vssd1 vssd1 vccd1 vccd1
+ _01634_ sky130_fd_sc_hd__mux2_2
X_08537_ datapath.rf.registers\[29\]\[0\] net797 _03372_ net875 vssd1 vssd1 vccd1
+ vccd1 _03373_ sky130_fd_sc_hd__a211o_1
XANTENNA__13933__RESET_B net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout437_X net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08468_ datapath.rf.registers\[2\]\[1\] _01713_ _01772_ datapath.rf.registers\[15\]\[1\]
+ _03302_ vssd1 vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__a221o_1
XANTENNA__07286__A2 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07419_ net872 _02250_ _02252_ _02254_ vssd1 vssd1 vccd1 vccd1 _02255_ sky130_fd_sc_hd__or4_1
XFILLER_149_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08399_ datapath.rf.registers\[27\]\[2\] net980 net939 vssd1 vssd1 vccd1 vccd1 _03235_
+ sky130_fd_sc_hd__and3_1
XANTENNA__13003__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12567__B1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10430_ _05264_ _05265_ _05249_ vssd1 vssd1 vccd1 vccd1 _05266_ sky130_fd_sc_hd__a21o_1
XANTENNA__07038__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10361_ _04848_ _05196_ vssd1 vssd1 vccd1 vccd1 _05197_ sky130_fd_sc_hd__or2_1
XANTENNA__12842__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12100_ screen.register.currentXbus\[15\] _05768_ _05772_ screen.register.currentXbus\[31\]
+ _06137_ vssd1 vssd1 vccd1 vccd1 _06138_ sky130_fd_sc_hd__a221o_1
XANTENNA__07994__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13080_ net1935 net219 net386 vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__mux2_1
XFILLER_124_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10292_ datapath.PC\[5\] _04454_ net468 vssd1 vssd1 vccd1 vccd1 _05128_ sky130_fd_sc_hd__mux2_1
XFILLER_152_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout973_X net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11458__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12031_ _05328_ _06003_ vssd1 vssd1 vccd1 vccd1 _06073_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_57_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09735__A1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08538__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold180 screen.controlBus\[5\] vssd1 vssd1 vccd1 vccd1 net1528 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold191 datapath.rf.registers\[4\]\[24\] vssd1 vssd1 vccd1 vccd1 net1539 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08340__B net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout660 net663 vssd1 vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__buf_4
Xfanout671 net674 vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__buf_4
Xfanout682 _01828_ vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__buf_2
X_13982_ clknet_leaf_107_clk _00759_ net1221 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_70_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout693 _01824_ vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__buf_4
XFILLER_19_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_831 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12933_ net300 net1978 net395 vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__mux2_1
XANTENNA__11193__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12864_ net258 net1794 net400 vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__mux2_1
XFILLER_33_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14603_ clknet_leaf_56_clk _01308_ net1161 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[5\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11815_ datapath.ru.latched_instruction\[21\] net334 net314 _01505_ vssd1 vssd1 vccd1
+ vccd1 _00681_ sky130_fd_sc_hd__a22o_1
X_12795_ net170 net2245 net495 vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__mux2_1
X_11746_ net1493 net144 net138 _03076_ vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__a22o_1
X_14534_ clknet_leaf_28_clk _01239_ net1133 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07277__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12270__A2 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11677_ _05157_ net154 net150 net1396 vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__a22o_1
X_14465_ clknet_leaf_37_clk _01170_ net1171 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10628_ net1037 _05447_ vssd1 vssd1 vccd1 vccd1 _05448_ sky130_fd_sc_hd__nor2_1
X_13416_ clknet_leaf_65_clk _00226_ net1238 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[10\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_139_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12022__A2 _06018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14396_ clknet_leaf_8_clk _01101_ net1072 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_40_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13347_ clknet_leaf_139_clk _00157_ net1099 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[22\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_143_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10559_ screen.register.currentXbus\[21\] screen.register.currentXbus\[20\] screen.register.currentXbus\[23\]
+ screen.register.currentXbus\[22\] vssd1 vssd1 vccd1 vccd1 _05383_ sky130_fd_sc_hd__or4_1
XANTENNA__12752__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07985__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13278_ clknet_leaf_150_clk _00088_ net1059 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[27\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11368__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08529__A2 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12229_ _06228_ _06229_ vssd1 vssd1 vccd1 vccd1 _00771_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_90_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07737__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07201__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07770_ datapath.rf.registers\[12\]\[15\] net827 _02603_ _02604_ _02605_ vssd1 vssd1
+ vccd1 vccd1 _02606_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_108_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06986__A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06721_ _01534_ _01551_ _01558_ vssd1 vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__and3_1
XANTENNA__13880__Q datapath.ru.latched_instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08162__B1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09440_ _03569_ _04273_ vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__xnor2_1
X_06652_ datapath.ru.latched_instruction\[10\] _01490_ vssd1 vssd1 vccd1 vccd1 _01491_
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_88_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_121_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09371_ net555 _04183_ _04206_ _04180_ net631 vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__a32o_2
XANTENNA__08409__C _01720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06583_ net1273 vssd1 vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__inv_2
XANTENNA__07313__C net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10795__X _05556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12927__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08322_ datapath.rf.registers\[13\]\[4\] net691 net683 datapath.rf.registers\[27\]\[4\]
+ _03152_ vssd1 vssd1 vccd1 vccd1 _03158_ sky130_fd_sc_hd__a221o_1
XANTENNA__08706__A net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08253_ datapath.rf.registers\[18\]\[5\] net792 _03086_ _03088_ vssd1 vssd1 vccd1
+ vccd1 _03089_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout132_A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07204_ datapath.rf.registers\[23\]\[27\] net699 net680 datapath.rf.registers\[6\]\[27\]
+ _02039_ vssd1 vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__a221o_1
XANTENNA__12549__B1 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08184_ datapath.rf.registers\[20\]\[7\] net720 net670 datapath.rf.registers\[21\]\[7\]
+ _03010_ vssd1 vssd1 vccd1 vccd1 _03020_ sky130_fd_sc_hd__a221o_1
Xteam_04_1302 vssd1 vssd1 vccd1 vccd1 team_04_1302/HI gpio_oeb[11] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_119_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xteam_04_1313 vssd1 vssd1 vccd1 vccd1 team_04_1313/HI gpio_out[6] sky130_fd_sc_hd__conb_1
Xteam_04_1324 vssd1 vssd1 vccd1 vccd1 team_04_1324/HI gpio_out[28] sky130_fd_sc_hd__conb_1
X_07135_ datapath.rf.registers\[11\]\[28\] net883 net802 datapath.rf.registers\[3\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__a22o_1
XFILLER_145_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xteam_04_1335 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] team_04_1335/LO sky130_fd_sc_hd__conb_1
XANTENNA_fanout1041_A net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xteam_04_1346 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] team_04_1346/LO sky130_fd_sc_hd__conb_1
XANTENNA__07976__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1139_A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11786__B datapath.ack_mul vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07066_ datapath.rf.registers\[23\]\[30\] net700 net693 datapath.rf.registers\[13\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__a22o_1
XANTENNA__07440__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11278__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09178__C1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout599_A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07728__B1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout766_A net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout387_X net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07968_ datapath.rf.registers\[0\]\[11\] net868 _02803_ vssd1 vssd1 vccd1 vccd1 _02804_
+ sky130_fd_sc_hd__o21a_2
XFILLER_102_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_52_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06919_ net954 net923 vssd1 vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__and2_1
X_09707_ net358 _04361_ _04542_ net345 vssd1 vssd1 vccd1 vccd1 _04543_ sky130_fd_sc_hd__a211o_1
XFILLER_74_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout933_A _01725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07899_ _02733_ _02734_ vssd1 vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__or2_1
XFILLER_28_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07504__B _01707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09638_ _04470_ _04473_ _04472_ net630 vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__07900__B1 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09569_ _04376_ _04378_ net362 vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout721_X net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07223__C net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12837__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout819_X net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11600_ _05758_ _05823_ vssd1 vssd1 vccd1 vccd1 _05824_ sky130_fd_sc_hd__nor2_1
XFILLER_12_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_139_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12580_ datapath.mulitply_result\[12\] datapath.multiplication_module.multiplicand_i\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06430_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_156_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_156_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11531_ net1009 _05753_ _05754_ vssd1 vssd1 vccd1 vccd1 _05755_ sky130_fd_sc_hd__nor3_2
XFILLER_7_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10584__C _02934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14250_ clknet_leaf_59_clk _00955_ net1169 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[15\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11462_ net1637 net221 net406 vssd1 vssd1 vccd1 vccd1 _00500_ sky130_fd_sc_hd__mux2_1
XANTENNA__12004__A2 _05786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13201_ clknet_leaf_35_clk _00011_ net1130 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_59_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10413_ net643 _05247_ _05248_ vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__or3_1
XANTENNA__08054__C net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14181_ clknet_leaf_50_clk _00936_ net1175 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11393_ net2524 net244 net410 vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__mux2_1
XFILLER_137_696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13132_ net1953 net298 net382 vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__mux2_1
X_10344_ datapath.PC\[10\] _04561_ net466 vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__mux2_1
XFILLER_136_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07431__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07893__C net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11188__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_72_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13063_ net1896 net259 net389 vssd1 vssd1 vccd1 vccd1 _01306_ sky130_fd_sc_hd__mux2_1
XFILLER_79_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10275_ net1044 _05110_ _05109_ net639 vssd1 vssd1 vccd1 vccd1 _05111_ sky130_fd_sc_hd__a211o_1
XFILLER_2_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07719__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12014_ _06057_ net1435 _06017_ vssd1 vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__mux2_1
XFILLER_105_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06927__D1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout490 _06551_ vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__buf_6
XANTENNA__07254__X _02090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13965_ clknet_leaf_106_clk _00743_ net1223 vssd1 vssd1 vccd1 vccd1 screen.counter.ct\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08144__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload8_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12916_ net1730 net233 net484 vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__mux2_1
X_13896_ clknet_leaf_44_clk net1484 net1152 vssd1 vssd1 vccd1 vccd1 keypad.decode.sticky\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06774__A1_N _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12747__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12847_ net239 net2229 net488 vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__mux2_1
X_12778_ net253 net1666 net494 vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__mux2_1
XANTENNA__08447__B2 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10254__A1 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14517_ clknet_leaf_130_clk _01222_ net1115 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[29\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11729_ net16 net1033 net1023 net1436 vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__o22a_1
XANTENNA__10494__C _05314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08960__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14448_ clknet_leaf_24_clk _01153_ net1158 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[16\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_128_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12482__S net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold905 datapath.rf.registers\[26\]\[28\] vssd1 vssd1 vccd1 vccd1 net2253 sky130_fd_sc_hd__dlygate4sd3_1
X_14379_ clknet_leaf_55_clk _01084_ net1179 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[30\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold916 datapath.rf.registers\[8\]\[11\] vssd1 vssd1 vccd1 vccd1 net2264 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11754__B2 _02680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold927 datapath.rf.registers\[19\]\[2\] vssd1 vssd1 vccd1 vccd1 net2275 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_142_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07422__A2 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold938 datapath.rf.registers\[27\]\[4\] vssd1 vssd1 vccd1 vccd1 net2286 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13875__Q datapath.ru.latched_instruction\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold949 datapath.rf.registers\[18\]\[18\] vssd1 vssd1 vccd1 vccd1 net2297 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11098__S net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08940_ net357 _03775_ vssd1 vssd1 vccd1 vccd1 _03776_ sky130_fd_sc_hd__or2_1
XFILLER_143_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08871_ _03703_ _03706_ net342 vssd1 vssd1 vccd1 vccd1 _03707_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08383__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07822_ datapath.rf.registers\[6\]\[14\] net824 _02641_ _02647_ _02657_ vssd1 vssd1
+ vccd1 vccd1 _02658_ sky130_fd_sc_hd__a2111o_1
XFILLER_85_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07605__A _02418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07753_ net561 _02588_ vssd1 vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__and2_1
XANTENNA__08135__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06704_ datapath.ru.latched_instruction\[28\] datapath.ru.latched_instruction\[29\]
+ datapath.ru.latched_instruction\[30\] datapath.ru.latched_instruction\[31\] vssd1
+ vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__or4_1
XFILLER_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07489__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07684_ _02508_ _02509_ _02519_ vssd1 vssd1 vccd1 vccd1 _02520_ sky130_fd_sc_hd__or3b_1
XFILLER_25_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09423_ net367 _04257_ _04258_ vssd1 vssd1 vccd1 vccd1 _04259_ sky130_fd_sc_hd__a21o_1
X_06635_ mmio.memload_or_instruction\[11\] net1051 vssd1 vssd1 vccd1 vccd1 _01474_
+ sky130_fd_sc_hd__and2_1
X_09354_ net353 _04188_ _04189_ vssd1 vssd1 vccd1 vccd1 _04190_ sky130_fd_sc_hd__and3_1
X_06566_ datapath.pc_module.i_ack1 vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_23_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08305_ datapath.rf.registers\[3\]\[4\] net802 net800 datapath.rf.registers\[15\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__a22o_1
XANTENNA__06882__C _01656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09285_ _03578_ _04119_ _03604_ vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout135_X net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout514_A _05731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1256_A net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08236_ datapath.rf.registers\[26\]\[6\] net778 net671 datapath.rf.registers\[7\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_134_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08167_ datapath.rf.registers\[13\]\[7\] net812 _02991_ _02992_ _03002_ vssd1 vssd1
+ vccd1 vccd1 _03003_ sky130_fd_sc_hd__a2111oi_1
XANTENNA_fanout1044_X net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07118_ datapath.rf.registers\[0\]\[29\] net784 _01950_ _01953_ vssd1 vssd1 vccd1
+ vccd1 _01954_ sky130_fd_sc_hd__o22a_4
XANTENNA__11745__B2 _03123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07413__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08098_ datapath.rf.registers\[0\]\[9\] net783 _02933_ vssd1 vssd1 vccd1 vccd1 _02934_
+ sky130_fd_sc_hd__o21ba_4
XANTENNA_fanout883_A _01719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07049_ datapath.rf.registers\[27\]\[30\] net809 net806 datapath.rf.registers\[28\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__a22o_1
XFILLER_134_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10060_ datapath.PC\[29\] net595 vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__nand2_1
XFILLER_87_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07218__C net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout671_X net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout769_X net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08374__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11308__Y _05726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08126__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout936_X net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10579__C _02311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13750_ clknet_leaf_88_clk _00559_ net1252 vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__dfrtp_1
X_10962_ _01500_ net655 _05698_ _05699_ vssd1 vssd1 vccd1 vccd1 _05700_ sky130_fd_sc_hd__o22a_1
X_12701_ _01432_ _01434_ vssd1 vssd1 vccd1 vccd1 _06531_ sky130_fd_sc_hd__or2_1
XANTENNA__08049__C net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10893_ datapath.mulitply_result\[23\] net599 _05635_ _05639_ net618 vssd1 vssd1
+ vccd1 vccd1 _05640_ sky130_fd_sc_hd__a221o_1
X_13681_ clknet_leaf_41_clk _00491_ net1142 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[14\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11471__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12632_ _06471_ _06472_ _06473_ _06466_ vssd1 vssd1 vccd1 vccd1 _06474_ sky130_fd_sc_hd__a211o_1
XANTENNA__06792__C _01585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12563_ datapath.mulitply_result\[9\] datapath.multiplication_module.multiplicand_i\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06416_ sky130_fd_sc_hd__nor2_1
X_14302_ clknet_leaf_147_clk _01007_ net1064 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[0\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11514_ _05336_ _05342_ _05738_ vssd1 vssd1 vccd1 vccd1 _05739_ sky130_fd_sc_hd__a21o_1
XFILLER_145_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12494_ net245 net2472 net506 vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__mux2_1
XANTENNA__07652__A2 _02487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14233_ clknet_leaf_123_clk datapath.multiplication_module.multiplier_i_n\[1\] net1215
+ vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplier_i\[1\] sky130_fd_sc_hd__dfrtp_1
X_11445_ datapath.rf.registers\[14\]\[1\] net260 net409 vssd1 vssd1 vccd1 vccd1 _00483_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__10815__S net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14164_ clknet_leaf_66_clk _00919_ net1237 vssd1 vssd1 vccd1 vccd1 datapath.mulitply_result\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_124_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14054__RESET_B net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07404__A2 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11376_ _05696_ _05729_ vssd1 vssd1 vccd1 vccd1 _05730_ sky130_fd_sc_hd__nor2_4
XANTENNA__08512__C _01831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_156_Right_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10327_ net896 _04584_ _05162_ _05161_ net228 vssd1 vssd1 vccd1 vccd1 _05163_ sky130_fd_sc_hd__o311a_1
X_13115_ net232 net2519 net471 vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__mux2_1
X_14095_ clknet_leaf_110_clk _00861_ net1222 vssd1 vssd1 vccd1 vccd1 screen.register.currentXbus\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07409__B net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09905__A _01585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13046_ net239 net1965 net476 vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__mux2_1
X_10258_ net223 _05093_ net1292 vssd1 vssd1 vccd1 vccd1 _05094_ sky130_fd_sc_hd__a21o_1
XFILLER_140_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1230 net1231 vssd1 vssd1 vccd1 vccd1 net1230 sky130_fd_sc_hd__clkbuf_2
XFILLER_94_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08365__B1 _01753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1241 net1251 vssd1 vssd1 vccd1 vccd1 net1241 sky130_fd_sc_hd__clkbuf_4
X_10189_ datapath.PC\[17\] net467 net1040 vssd1 vssd1 vccd1 vccd1 _05025_ sky130_fd_sc_hd__o21ai_1
Xfanout1252 net1261 vssd1 vssd1 vccd1 vccd1 net1252 sky130_fd_sc_hd__clkbuf_4
Xfanout1263 datapath.PC\[26\] vssd1 vssd1 vccd1 vccd1 net1263 sky130_fd_sc_hd__buf_2
Xfanout1274 screen.counter.ct\[12\] vssd1 vssd1 vccd1 vccd1 net1274 sky130_fd_sc_hd__buf_2
XFILLER_120_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1285 mmio.key_en2 vssd1 vssd1 vccd1 vccd1 net1285 sky130_fd_sc_hd__clkbuf_2
XFILLER_66_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13110__A0 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08117__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13948_ clknet_leaf_103_clk _00726_ net1225 vssd1 vssd1 vccd1 vccd1 screen.dcx sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_85_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06679__B1 _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11672__B1 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13879_ clknet_leaf_53_clk _00683_ net1183 vssd1 vssd1 vccd1 vccd1 datapath.ru.latched_instruction\[23\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_35_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11381__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09617__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09093__A1 _02170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09070_ _03903_ _03905_ net340 vssd1 vssd1 vccd1 vccd1 _03906_ sky130_fd_sc_hd__mux2_1
XANTENNA__07643__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08840__A1 _03296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08021_ datapath.rf.registers\[0\]\[10\] net868 _02855_ vssd1 vssd1 vccd1 vccd1 _02857_
+ sky130_fd_sc_hd__o21ai_4
XANTENNA__06851__B1 _01598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold702 datapath.rf.registers\[20\]\[18\] vssd1 vssd1 vccd1 vccd1 net2050 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13101__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold713 datapath.rf.registers\[28\]\[23\] vssd1 vssd1 vccd1 vccd1 net2061 sky130_fd_sc_hd__dlygate4sd3_1
Xhold724 datapath.rf.registers\[9\]\[1\] vssd1 vssd1 vccd1 vccd1 net2072 sky130_fd_sc_hd__dlygate4sd3_1
Xhold735 datapath.rf.registers\[19\]\[12\] vssd1 vssd1 vccd1 vccd1 net2083 sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 datapath.rf.registers\[29\]\[2\] vssd1 vssd1 vccd1 vccd1 net2094 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold757 datapath.rf.registers\[1\]\[1\] vssd1 vssd1 vccd1 vccd1 net2105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold768 mmio.memload_or_instruction\[11\] vssd1 vssd1 vccd1 vccd1 net2116 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09972_ _04743_ _04807_ vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__nand2_1
XFILLER_131_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12940__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold779 datapath.rf.registers\[11\]\[26\] vssd1 vssd1 vccd1 vccd1 net2127 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_123_Right_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08923_ net991 net576 vssd1 vssd1 vccd1 vccd1 _03759_ sky130_fd_sc_hd__nand2_1
XFILLER_58_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08356__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout297_A _05536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09553__C1 _03613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08854_ _02419_ _02467_ net444 vssd1 vssd1 vccd1 vccd1 _03690_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1004_A net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_894 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07805_ datapath.rf.registers\[21\]\[14\] net946 net923 vssd1 vssd1 vccd1 vccd1 _02641_
+ sky130_fd_sc_hd__and3_1
X_08785_ net990 _03228_ _03615_ vssd1 vssd1 vccd1 vccd1 _03621_ sky130_fd_sc_hd__mux2_1
XANTENNA__08108__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout464_A _03104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09305__C1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07736_ datapath.rf.registers\[12\]\[16\] net754 net698 datapath.rf.registers\[23\]\[16\]
+ _02569_ vssd1 vssd1 vccd1 vccd1 _02572_ sky130_fd_sc_hd__a221o_1
XFILLER_44_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07667_ datapath.rf.registers\[5\]\[17\] net947 net935 vssd1 vssd1 vccd1 vccd1 _02503_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout631_A net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11291__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout729_A _01812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06618_ datapath.ru.latched_instruction\[22\] _01456_ vssd1 vssd1 vccd1 vccd1 _01457_
+ sky130_fd_sc_hd__xor2_1
X_09406_ _03572_ _04240_ net580 vssd1 vssd1 vccd1 vccd1 _04242_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07882__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07598_ _02422_ _02424_ _02430_ _02432_ vssd1 vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__or4_1
XFILLER_139_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09084__A1 _02169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09337_ _03516_ _03718_ _04170_ net642 vssd1 vssd1 vccd1 vccd1 _04173_ sky130_fd_sc_hd__o211a_1
XANTENNA__07501__C net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout517_X net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1259_X net1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07095__B1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09268_ _04102_ _04103_ net349 vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07634__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08219_ datapath.rf.registers\[3\]\[6\] net801 net799 datapath.rf.registers\[15\]\[6\]
+ _03054_ vssd1 vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__a221o_1
XFILLER_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09199_ net380 _04034_ net312 vssd1 vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__o21bai_1
XANTENNA__13011__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11230_ net211 net2463 net526 vssd1 vssd1 vccd1 vccd1 _00280_ sky130_fd_sc_hd__mux2_1
XFILLER_107_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12135__B net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout886_X net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11161_ net233 net1743 net530 vssd1 vssd1 vccd1 vccd1 _00214_ sky130_fd_sc_hd__mux2_1
XFILLER_136_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12850__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10112_ net1041 _04945_ _04947_ net640 vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11092_ net238 net2313 net536 vssd1 vssd1 vccd1 vccd1 _00149_ sky130_fd_sc_hd__mux2_1
XFILLER_110_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11466__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10043_ _04818_ _04832_ _04724_ vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__a21o_1
XFILLER_76_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10154__B1 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12449__A1_N net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold40 mmio.memload_or_instruction\[28\] vssd1 vssd1 vccd1 vccd1 net1388 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold51 screen.controlBus\[26\] vssd1 vssd1 vccd1 vccd1 net1399 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 screen.controlBus\[17\] vssd1 vssd1 vccd1 vccd1 net1410 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input25_A DAT_I[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold73 net62 vssd1 vssd1 vccd1 vccd1 net1421 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 net45 vssd1 vssd1 vccd1 vccd1 net1432 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 net50 vssd1 vssd1 vccd1 vccd1 net1443 sky130_fd_sc_hd__dlygate4sd3_1
X_13802_ clknet_leaf_52_clk _00611_ net1183 vssd1 vssd1 vccd1 vccd1 mmio.memload_or_instruction\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11994_ _05325_ _05752_ vssd1 vssd1 vccd1 vccd1 _06038_ sky130_fd_sc_hd__nor2_1
XFILLER_91_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10457__A1 _04909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13733_ clknet_leaf_116_clk _00543_ net1188 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12297__S net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10945_ net174 net2438 net543 vssd1 vssd1 vccd1 vccd1 _00032_ sky130_fd_sc_hd__mux2_1
X_13664_ clknet_leaf_138_clk _00474_ net1112 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10876_ net898 _05624_ vssd1 vssd1 vccd1 vccd1 _05625_ sky130_fd_sc_hd__nor2_1
XANTENNA__07873__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08507__C _01831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12615_ _06457_ _06458_ _06456_ vssd1 vssd1 vccd1 vccd1 _06460_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07411__C net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13595_ clknet_leaf_38_clk _00405_ net1145 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07209__A2_N net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07086__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07625__A2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12546_ _06400_ _06401_ vssd1 vssd1 vccd1 vccd1 _06402_ sky130_fd_sc_hd__nand2_1
XFILLER_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12477_ _05518_ _06370_ vssd1 vssd1 vccd1 vccd1 _06371_ sky130_fd_sc_hd__or2_1
XANTENNA_4 datapath.multiplication_module.multiplicand_i_n\[15\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14216_ clknet_leaf_50_clk datapath.multiplication_module.multiplicand_i_n\[27\]
+ net1175 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11428_ net218 net1815 net514 vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__mux2_1
XFILLER_141_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12760__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14147_ clknet_leaf_150_clk _00904_ net1053 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[31\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11359_ net244 net2602 net519 vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__mux2_1
XFILLER_4_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06611__X _01450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14078_ clknet_leaf_111_clk _00845_ net1199 vssd1 vssd1 vccd1 vccd1 screen.controlBus\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_140_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09535__C1 _02857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13029_ net207 net2340 net477 vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__mux2_1
XFILLER_79_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08889__A1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1060 net1061 vssd1 vssd1 vccd1 vccd1 net1060 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07010__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1071 net1072 vssd1 vssd1 vccd1 vccd1 net1071 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10696__A1 _03357_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_6_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1082 net1084 vssd1 vssd1 vccd1 vccd1 net1082 sky130_fd_sc_hd__clkbuf_4
Xfanout1093 net1096 vssd1 vssd1 vccd1 vccd1 net1093 sky130_fd_sc_hd__clkbuf_4
XFILLER_67_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08570_ datapath.rf.registers\[4\]\[0\] _01636_ net990 net968 net913 vssd1 vssd1
+ vccd1 vccd1 _03406_ sky130_fd_sc_hd__o2111a_1
X_07521_ datapath.rf.registers\[6\]\[20\] net824 _02342_ _02343_ _02344_ vssd1 vssd1
+ vccd1 vccd1 _02357_ sky130_fd_sc_hd__a2111o_1
XFILLER_23_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07452_ datapath.rf.registers\[2\]\[21\] net981 net949 vssd1 vssd1 vccd1 vccd1 _02288_
+ sky130_fd_sc_hd__and3_1
XFILLER_22_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07864__A2 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07383_ datapath.rf.registers\[11\]\[23\] net710 net698 datapath.rf.registers\[23\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__a22o_1
XANTENNA__12935__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09122_ _03633_ _03957_ net378 vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__mux2_1
XFILLER_148_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12070__B1 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07616__A2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08714__A _03263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09053_ net356 _03888_ vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_98_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08004_ datapath.rf.registers\[28\]\[10\] net806 net797 datapath.rf.registers\[29\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02840_ sky130_fd_sc_hd__a22o_1
Xhold510 datapath.rf.registers\[12\]\[8\] vssd1 vssd1 vccd1 vccd1 net1858 sky130_fd_sc_hd__dlygate4sd3_1
Xhold521 datapath.rf.registers\[20\]\[21\] vssd1 vssd1 vccd1 vccd1 net1869 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold532 datapath.rf.registers\[4\]\[4\] vssd1 vssd1 vccd1 vccd1 net1880 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08152__C _01720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold543 datapath.rf.registers\[11\]\[4\] vssd1 vssd1 vccd1 vccd1 net1891 sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 datapath.rf.registers\[23\]\[3\] vssd1 vssd1 vccd1 vccd1 net1902 sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 datapath.rf.registers\[18\]\[24\] vssd1 vssd1 vccd1 vccd1 net1913 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1121_A _00004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold576 datapath.rf.registers\[10\]\[6\] vssd1 vssd1 vccd1 vccd1 net1924 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1219_A net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold587 datapath.rf.registers\[5\]\[18\] vssd1 vssd1 vccd1 vccd1 net1935 sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 datapath.rf.registers\[30\]\[25\] vssd1 vssd1 vccd1 vccd1 net1946 sky130_fd_sc_hd__dlygate4sd3_1
X_09955_ _04788_ _04789_ _04775_ vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__a21oi_1
XFILLER_131_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08329__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11286__S net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06888__B net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout679_A _01828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08906_ datapath.PC\[16\] _03741_ vssd1 vssd1 vccd1 vccd1 _03742_ sky130_fd_sc_hd__or2_1
X_09886_ datapath.PC\[24\] net594 vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__xnor2_1
XFILLER_112_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1210 datapath.rf.registers\[5\]\[6\] vssd1 vssd1 vccd1 vccd1 net2558 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1221 screen.register.currentYbus\[28\] vssd1 vssd1 vccd1 vccd1 net2569 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07001__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1232 datapath.rf.registers\[16\]\[29\] vssd1 vssd1 vccd1 vccd1 net2580 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1243 datapath.rf.registers\[17\]\[31\] vssd1 vssd1 vccd1 vccd1 net2591 sky130_fd_sc_hd__dlygate4sd3_1
X_08837_ _03669_ _03672_ vssd1 vssd1 vccd1 vccd1 _03673_ sky130_fd_sc_hd__nor2_2
XFILLER_85_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout846_A _01737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1254 datapath.rf.registers\[20\]\[16\] vssd1 vssd1 vccd1 vccd1 net2602 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1265 datapath.rf.registers\[31\]\[31\] vssd1 vssd1 vccd1 vccd1 net2613 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1276 datapath.rf.registers\[0\]\[24\] vssd1 vssd1 vccd1 vccd1 net2624 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1287 screen.register.currentYbus\[10\] vssd1 vssd1 vccd1 vccd1 net2635 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1298 mmio.key_data\[2\] vssd1 vssd1 vccd1 vccd1 net2646 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12428__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_748 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08768_ _03602_ _03603_ vssd1 vssd1 vccd1 vccd1 _03604_ sky130_fd_sc_hd__and2_4
XTAP_TAPCELL_ROW_49_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10439__A1 _01702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07719_ datapath.rf.registers\[31\]\[16\] net793 net790 datapath.rf.registers\[18\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__a22o_1
XFILLER_82_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout634_X net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08699_ _02857_ _02879_ vssd1 vssd1 vccd1 vccd1 _03535_ sky130_fd_sc_hd__and2_1
XANTENNA__13006__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07512__B net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10730_ net1546 net569 vssd1 vssd1 vccd1 vccd1 datapath.multiplication_module.multiplicand_i_n\[16\]
+ sky130_fd_sc_hd__and2_1
XFILLER_53_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07855__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10661_ _05428_ _05445_ _05479_ vssd1 vssd1 vccd1 vccd1 _05480_ sky130_fd_sc_hd__or3_1
XFILLER_13_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout801_X net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12845__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12400_ net1382 net131 _06347_ vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__a21o_1
XANTENNA__07068__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_149_Left_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13380_ clknet_leaf_17_clk _00190_ net1109 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[9\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10592_ _02439_ _02487_ _02542_ _02587_ vssd1 vssd1 vccd1 vccd1 _05415_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_11_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12331_ net640 _06302_ _04960_ vssd1 vssd1 vccd1 vccd1 _06303_ sky130_fd_sc_hd__o21bai_1
XANTENNA__08280__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10592__C _02542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08343__B net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12262_ _05002_ net306 vssd1 vssd1 vccd1 vccd1 _06252_ sky130_fd_sc_hd__nand2_1
X_14001_ clknet_leaf_114_clk _00778_ net1196 vssd1 vssd1 vccd1 vccd1 screen.counter.currentCt\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11213_ net296 net1959 net526 vssd1 vssd1 vccd1 vccd1 _00263_ sky130_fd_sc_hd__mux2_1
X_12193_ _06205_ _06206_ net567 vssd1 vssd1 vccd1 vccd1 _00758_ sky130_fd_sc_hd__and3b_1
XANTENNA__08032__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput41 net41 vssd1 vssd1 vccd1 vccd1 ADR_O[10] sky130_fd_sc_hd__buf_2
Xoutput52 net52 vssd1 vssd1 vccd1 vccd1 ADR_O[20] sky130_fd_sc_hd__buf_2
XANTENNA__07527__X _02363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11144_ net302 net2329 net533 vssd1 vssd1 vccd1 vccd1 _00197_ sky130_fd_sc_hd__mux2_1
XFILLER_1_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput63 net63 vssd1 vssd1 vccd1 vccd1 ADR_O[30] sky130_fd_sc_hd__buf_2
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 DAT_O[10] sky130_fd_sc_hd__buf_2
XFILLER_122_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput85 net85 vssd1 vssd1 vccd1 vccd1 DAT_O[20] sky130_fd_sc_hd__buf_2
XFILLER_122_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11196__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput96 net96 vssd1 vssd1 vccd1 vccd1 DAT_O[30] sky130_fd_sc_hd__buf_2
XFILLER_110_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11075_ net286 net1736 net537 vssd1 vssd1 vccd1 vccd1 _00132_ sky130_fd_sc_hd__mux2_1
XANTENNA__10127__B1 net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10026_ _04742_ _04743_ vssd1 vssd1 vccd1 vccd1 _04862_ sky130_fd_sc_hd__and2b_1
XANTENNA__10888__X _05635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11977_ _05846_ _05860_ vssd1 vssd1 vccd1 vccd1 _06022_ sky130_fd_sc_hd__nor2_1
XANTENNA__08077__Y _02913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08518__B net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13716_ clknet_leaf_128_clk _00526_ net1210 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[19\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10928_ net1045 net653 _05668_ _05669_ vssd1 vssd1 vccd1 vccd1 _05670_ sky130_fd_sc_hd__o22a_2
XFILLER_32_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14696_ clknet_leaf_64_clk _01401_ net1233 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[17\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12755__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13647_ clknet_leaf_26_clk _00457_ net1135 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[24\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10859_ net218 net2478 net542 vssd1 vssd1 vccd1 vccd1 _00020_ sky130_fd_sc_hd__mux2_1
XFILLER_31_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07059__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08256__C1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13578_ clknet_leaf_21_clk _00388_ net1164 vssd1 vssd1 vccd1 vccd1 datapath.rf.registers\[20\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06980__C _01647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12529_ _06381_ _06383_ _06380_ vssd1 vssd1 vccd1 vccd1 _06388_ sky130_fd_sc_hd__o21ba_1
XANTENNA__08271__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12490__S net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08023__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09220__A1 _03607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06989__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07231__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09365__A _03613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout308 _06246_ vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__clkbuf_4
XFILLER_87_807 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout319 _03684_ vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__buf_2
XFILLER_87_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06952_ _01636_ net990 net970 vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__and3_1
X_09740_ net324 _03818_ vssd1 vssd1 vccd1 vccd1 _04576_ sky130_fd_sc_hd__nor2_1
.ends

