module t07_display(
    input logic clk, nrst,
    
    output logic [15:0] out
    //output logic delay 
);

    logic [17:0] counter, next_ctr;

    always_ff @(posedge clk, negedge nrst) begin 
        if (~nrst) begin
            counter <= '0;
        end else begin
            counter <= next_ctr;
        end
    end

  always_comb begin
    next_ctr = counter + 1;
    //delay = 0;
    // out = '0;
    case (counter) 
        18'd0: out = 16'h80_00; 
        18'd3: out = 16'h40_00;
        18'd6: out = 16'h80_88;
        18'd9: out = 16'h00_0B;

        18'd139: out = 16'h80_89;
        18'd143: out = 16'h00_02;

        18'd273: out = 16'h80_10;
        18'd276: out = 16'h00_0C;
        18'd279: out = 16'h80_04;
        18'd282: out = 16'h00_81;

        18'd412: out = 16'h80_14;
        18'd415: out = 16'h00_63;
        18'd418: out = 16'h80_15;
        18'd421: out = 16'h00_00;
        18'd424: out = 16'h80_16;
        18'd427: out = 16'h00_03;
        18'd430: out = 16'h80_17;
        18'd433: out = 16'h00_03;
        18'd436: out = 16'h80_18;
        18'd439: out = 16'h00_0B;
        18'd442: out = 16'h80_19;
        18'd445: out = 16'h00_DF;
        18'd458: out = 16'h80_1A;
        18'd461: out = 16'h00_01;
        18'd464: out = 16'h80_1B;
        18'd467: out = 16'h00_1F;
        18'd470: out = 16'h80_1C;
        18'd473: out = 16'h00_00;
        18'd476: out = 16'h80_1D;
        18'd479: out = 16'h00_16;
        18'd482: out = 16'h80_1E;
        18'd485: out = 16'h00_00;
        18'd488: out = 16'h80_1F;
        18'd491: out = 16'h00_01;
        18'd494: out = 16'h80_30;
        18'd497: out = 16'h00_00;
        18'd500: out = 16'h80_31;
        18'd503: out = 16'h00_00;
        18'd506: out = 16'h80_34;
        18'd509: out = 16'h00_1F;
        18'd512: out = 16'h80_35;
        18'd515: out = 16'h00_03;
        18'd518: out = 16'h80_32;
        18'd521: out = 16'h00_00;
        18'd524: out = 16'h80_33;
        18'd527: out = 16'h00_00;
        18'd530: out = 16'h80_36;
        18'd533: out = 16'h00_DF;
        18'd536: out = 16'h80_37;
        18'd539: out = 16'h00_01;
        18'd542: out = 16'h80_8E;
        18'd545: out = 16'h00_80;


        18'd63045: out = 16'h80_01;
        18'd63048: out = 16'h00_80;
        18'd63051: out = 16'h80_C7;
        18'd63054: out = 16'h00_01;
        18'd63057: out = 16'h80_8A;
        18'd63060: out = 16'h00_8A;
        18'd63063: out = 16'h80_8B;
        18'd63066: out = 16'h00_80;
        18'd63069: out = 16'h80_91;
        18'd63072: out = 16'h00_00;
        18'd63075: out = 16'h80_92;
        18'd63078: out = 16'h00_00;
        18'd63081: out = 16'h80_93;
        18'd63084: out = 16'h00_00;
        18'd63087: out = 16'h80_94;
        18'd63090: out = 16'h00_00;
        18'd63093: out = 16'h80_95;
        18'd63096: out = 16'h00_1F;
        18'd63099: out = 16'h80_96;
        18'd63102: out = 16'h00_03;
        18'd63105: out = 16'h80_97;
        18'd63108: out = 16'h00_DF;
        18'd63111: out = 16'h80_98;
        18'd63114: out = 16'h00_01;
        18'd63117: out = 16'h80_63;
        18'd63120: out = 16'h00_00;
        18'd63123: out = 16'h80_64;
        18'd63126: out = 16'h00_00;
        18'd63129: out = 16'h80_65;
        18'd63132: out = 16'h00_00;
        18'd63135: out = 16'h80_90;
        18'd63138: out = 16'h00_B0;
        18'd63141: out = 16'h80_90;
        18'd63144: out = 16'h40_00;
        18'd63147: out = 16'h80_90;
        18'd63150: out = 16'h40_00;
        18'd63153: out = 16'h80_90;
        18'd63156: out = 16'h40_00;
        18'd63159: out = 16'h80_90;
        18'd63162: out = 16'h40_00;
        18'd63165: out = 16'h80_90;
        18'd63168: out = 16'h40_00;
        18'd63171: out = 16'h80_90;
        18'd63174: out = 16'h40_00;
        18'd63177: out = 16'h80_90;
        18'd63180: out = 16'h40_00;
        18'd63183: out = 16'h80_90;
        18'd63186: out = 16'h40_00;
        18'd63189: out = 16'h80_90;
        18'd63192: out = 16'h40_00;
        18'd63195: out = 16'h80_90;
        18'd63198: out = 16'h40_00;
        18'd63201: out = 16'h80_90;
        18'd63204: out = 16'h40_00;
        18'd63207: out = 16'h80_90;
        18'd63210: out = 16'h40_00;
        18'd63213: out = 16'h80_90;
        18'd63216: out = 16'h40_00;
        18'd63219: out = 16'h80_90;
        18'd63222: out = 16'h40_00;
        18'd63225: out = 16'h80_90;
        18'd63228: out = 16'h40_00;
        18'd63231: out = 16'h80_90;
        18'd63234: out = 16'h40_00;
        18'd63237: out = 16'h80_90;
        18'd63240: out = 16'h40_00;
        18'd63243: out = 16'h80_90;
        18'd63246: out = 16'h40_00;
        18'd63249: out = 16'h80_90;
        18'd63252: out = 16'h40_00;
        18'd63255: out = 16'h80_90;
        18'd63258: out = 16'h40_00;
        18'd63261: out = 16'h80_90;
        18'd63264: out = 16'h40_00;
        18'd63267: out = 16'h80_90;
        18'd63270: out = 16'h40_00;
        18'd63273: out = 16'h80_90;
        18'd63276: out = 16'h40_00;
        18'd63279: out = 16'h80_90;
        18'd63282: out = 16'h40_00;
        18'd63285: out = 16'h80_90;
        18'd63288: out = 16'h40_00;
        18'd63291: out = 16'h80_90;
        18'd63294: out = 16'h40_00;
        18'd63297: out = 16'h80_90;
        18'd63300: out = 16'h40_00;
        18'd63303: out = 16'h80_90;
        18'd63306: out = 16'h40_00;
        18'd63309: out = 16'h80_90;
        18'd63312: out = 16'h40_00;
        18'd63315: out = 16'h80_90;
        18'd63318: out = 16'h40_00;
        18'd63321: out = 16'h80_90;
        18'd63324: out = 16'h40_00;
        18'd63327: out = 16'h80_90;
        18'd63330: out = 16'h40_00;
        18'd63333: out = 16'h80_90;
        18'd63336: out = 16'h40_00;
        18'd63339: out = 16'h80_90;
        18'd63342: out = 16'h40_00;
        18'd63345: out = 16'h80_90;
        18'd63348: out = 16'h40_00;
        18'd63351: out = 16'h80_90;
        18'd63354: out = 16'h40_00;
        18'd63357: out = 16'h80_90;
        18'd63360: out = 16'h40_00;
        18'd63363: out = 16'h80_90;
        18'd63366: out = 16'h40_00;
        18'd63369: out = 16'h80_90;
        18'd63372: out = 16'h40_00;
        18'd63375: out = 16'h80_90;
        18'd63378: out = 16'h40_00;
        18'd63381: out = 16'h80_90;
        18'd63384: out = 16'h40_00;
        18'd63387: out = 16'h80_90;
        18'd63390: out = 16'h40_00;
        18'd63393: out = 16'h80_90;
        18'd63396: out = 16'h40_00;
        18'd63399: out = 16'h80_90;
        18'd63402: out = 16'h40_00;
        18'd63405: out = 16'h80_90;
        18'd63408: out = 16'h40_00;
        18'd63411: out = 16'h80_90;
        18'd63414: out = 16'h40_00;
        18'd63417: out = 16'h80_90;
        18'd63420: out = 16'h40_00;
        18'd63423: out = 16'h80_90;
        18'd63426: out = 16'h40_00;
        18'd63429: out = 16'h80_90;
        18'd63432: out = 16'h40_00;
        18'd63435: out = 16'h80_90;
        18'd63438: out = 16'h40_00;
        18'd63441: out = 16'h80_90;
        18'd63444: out = 16'h40_00;
        18'd63447: out = 16'h80_90;
        18'd63450: out = 16'h40_00;
        18'd63453: out = 16'h80_90;
        18'd63456: out = 16'h40_00;
        18'd63459: out = 16'h80_90;
        18'd63462: out = 16'h40_00;
        18'd63465: out = 16'h80_90;
        18'd63468: out = 16'h40_00;
        18'd63471: out = 16'h80_90;
        18'd63474: out = 16'h40_00;
        18'd63477: out = 16'h80_90;
        18'd63480: out = 16'h40_00;
        18'd63483: out = 16'h80_90;
        18'd63486: out = 16'h40_00;
        18'd63489: out = 16'h80_90;
        18'd63492: out = 16'h40_00;
        18'd63495: out = 16'h80_90;
        18'd63498: out = 16'h40_00;
        18'd63501: out = 16'h80_90;
        18'd63504: out = 16'h40_00;
        18'd63507: out = 16'h80_90;
        18'd63510: out = 16'h40_00;
        18'd63513: out = 16'h80_90;
        18'd63516: out = 16'h40_00;
        18'd63519: out = 16'h80_90;
        18'd63522: out = 16'h40_00;
        18'd63525: out = 16'h80_90;
        18'd63528: out = 16'h40_00;
        18'd63531: out = 16'h80_90;
        18'd63534: out = 16'h40_00;
        18'd63537: out = 16'h80_90;
        18'd63540: out = 16'h40_00;
        18'd63543: out = 16'h80_90;
        18'd63546: out = 16'h40_00;
        18'd63549: out = 16'h80_90;
        18'd63552: out = 16'h40_00;
        18'd63555: out = 16'h80_90;
        18'd63558: out = 16'h40_00;
        18'd63561: out = 16'h80_90;
        18'd63564: out = 16'h40_00;
        18'd63567: out = 16'h80_90;
        18'd63570: out = 16'h40_00;
        18'd63573: out = 16'h80_90;
        18'd63576: out = 16'h40_00;
        18'd63579: out = 16'h80_90;
        18'd63582: out = 16'h40_00;
        18'd63585: out = 16'h80_90;
        18'd63588: out = 16'h40_00;
        18'd63591: out = 16'h80_90;
        18'd63594: out = 16'h40_00;
        18'd63597: out = 16'h80_90;
        18'd63600: out = 16'h40_00;
        18'd63603: out = 16'h80_90;
        18'd63606: out = 16'h40_00;
        18'd63609: out = 16'h80_90;
        18'd63612: out = 16'h40_00;
        18'd63615: out = 16'h80_90;
        18'd63618: out = 16'h40_00;
        18'd63621: out = 16'h80_90;
        18'd63624: out = 16'h40_00;
        18'd63627: out = 16'h80_90;
        18'd63630: out = 16'h40_00;
        18'd63633: out = 16'h80_90;
        18'd63636: out = 16'h40_00;
        18'd63639: out = 16'h80_90;
        18'd63642: out = 16'h40_00;
        18'd63645: out = 16'h80_90;
        18'd63648: out = 16'h40_00;
        18'd63651: out = 16'h80_90;
        18'd63654: out = 16'h40_00;
        18'd63657: out = 16'h80_90;
        18'd63660: out = 16'h40_00;
        18'd63663: out = 16'h80_90;
        18'd63666: out = 16'h40_00;
        18'd63669: out = 16'h80_90;
        18'd63672: out = 16'h40_00;
        18'd63675: out = 16'h80_90;
        18'd63678: out = 16'h40_00;
        18'd63681: out = 16'h80_90;
        18'd63684: out = 16'h40_00;
        18'd63687: out = 16'h80_90;
        18'd63690: out = 16'h40_00;
        18'd63693: out = 16'h80_90;
        18'd63696: out = 16'h40_00;
        18'd63699: out = 16'h80_90;
        18'd63702: out = 16'h40_00;
        18'd63705: out = 16'h80_90;
        18'd63708: out = 16'h40_00;
        18'd63711: out = 16'h80_90;
        18'd63714: out = 16'h40_00;
        18'd63717: out = 16'h80_90;
        18'd63720: out = 16'h40_00;
        18'd63723: out = 16'h80_90;
        18'd63726: out = 16'h40_00;
        18'd63729: out = 16'h80_90;
        18'd63732: out = 16'h40_00;
        18'd63735: out = 16'h80_90;
        18'd63738: out = 16'h40_00;
        18'd63741: out = 16'h80_90;
        18'd63744: out = 16'h40_00;
        18'd63747: out = 16'h80_90;
        18'd63750: out = 16'h40_00;
        18'd63753: out = 16'h80_90;
        18'd63756: out = 16'h40_00;
        18'd63759: out = 16'h80_90;
        18'd63762: out = 16'h40_00;
        18'd63765: out = 16'h80_90;
        18'd63768: out = 16'h40_00;
        18'd63771: out = 16'h80_90;
        18'd63774: out = 16'h40_00;
        18'd63777: out = 16'h80_90;
        18'd63780: out = 16'h40_00;
        18'd63783: out = 16'h80_90;
        18'd63786: out = 16'h40_00;
        18'd63789: out = 16'h80_90;
        18'd63792: out = 16'h40_00;
        18'd63795: out = 16'h80_90;
        18'd63798: out = 16'h40_00;
        18'd63801: out = 16'h80_90;
        18'd63804: out = 16'h40_00;
        18'd63807: out = 16'h80_90;
        18'd63810: out = 16'h40_00;
        18'd63813: out = 16'h80_90;
        18'd63816: out = 16'h40_00;
        18'd63819: out = 16'h80_90;
        18'd63822: out = 16'h40_00;
        18'd63825: out = 16'h80_90;
        18'd63828: out = 16'h40_00;
        18'd63831: out = 16'h80_90;
        18'd63834: out = 16'h40_00;
        18'd63837: out = 16'h80_90;
        18'd63840: out = 16'h40_00;
        18'd63843: out = 16'h80_90;
        18'd63846: out = 16'h40_00;
        18'd63849: out = 16'h80_90;
        18'd63852: out = 16'h40_00;
        18'd63855: out = 16'h80_90;
        18'd63858: out = 16'h40_00;
        18'd63861: out = 16'h80_90;
        18'd63864: out = 16'h40_00;
        18'd63867: out = 16'h80_90;
        18'd63870: out = 16'h40_00;
        18'd63873: out = 16'h80_90;
        18'd63876: out = 16'h40_00;
        18'd63879: out = 16'h80_90;
        18'd63882: out = 16'h40_00;
        18'd63885: out = 16'h80_90;
        18'd63888: out = 16'h40_00;
        18'd63891: out = 16'h80_90;
        18'd63894: out = 16'h40_00;
        18'd63897: out = 16'h80_90;
        18'd63900: out = 16'h40_00;
        18'd63903: out = 16'h80_90;
        18'd63906: out = 16'h40_00;
        18'd63909: out = 16'h80_90;
        18'd63912: out = 16'h40_00;
        18'd63915: out = 16'h80_90;
        18'd63918: out = 16'h40_00;
        18'd63921: out = 16'h80_90;
        18'd63924: out = 16'h40_00;
        18'd63927: out = 16'h80_90;
        18'd63930: out = 16'h40_00;
        18'd63933: out = 16'h80_90;
        18'd63936: out = 16'h40_00;
        18'd63939: out = 16'h80_90;
        18'd63942: out = 16'h40_00;
        18'd63945: out = 16'h80_90;
        18'd63948: out = 16'h40_00;
        18'd63951: out = 16'h80_90;
        18'd63954: out = 16'h40_00;
        18'd63957: out = 16'h80_90;
        18'd63960: out = 16'h40_00;
        18'd63963: out = 16'h80_90;
        18'd63966: out = 16'h40_00;
        18'd63969: out = 16'h80_90;
        18'd63972: out = 16'h40_00;
        18'd63975: out = 16'h80_90;
        18'd63978: out = 16'h40_00;
        18'd63981: out = 16'h80_90;
        18'd63984: out = 16'h40_00;
        18'd63987: out = 16'h80_90;
        18'd63990: out = 16'h40_00;
        18'd63993: out = 16'h80_90;
        18'd63996: out = 16'h40_00;
        18'd63999: out = 16'h80_90;
        18'd64002: out = 16'h40_00;
        18'd64005: out = 16'h80_90;
        18'd64008: out = 16'h40_00;
        18'd64011: out = 16'h80_90;
        18'd64014: out = 16'h40_00;
        18'd64017: out = 16'h80_90;
        18'd64020: out = 16'h40_00;
        18'd64023: out = 16'h80_90;
        18'd64026: out = 16'h40_00;
        18'd64029: out = 16'h80_90;
        18'd64032: out = 16'h40_00;
        18'd64035: out = 16'h80_90;
        18'd64038: out = 16'h40_00;
        18'd64041: out = 16'h80_90;
        18'd64044: out = 16'h40_00;
        18'd64047: out = 16'h80_90;
        18'd64050: out = 16'h40_00;
        18'd64053: out = 16'h80_90;
        18'd64056: out = 16'h40_00;
        18'd64059: out = 16'h80_90;
        18'd64062: out = 16'h40_00;
        18'd64065: out = 16'h80_90;
        18'd64068: out = 16'h40_00;
        18'd64071: out = 16'h80_90;
        18'd64074: out = 16'h40_00;
        18'd64077: out = 16'h80_90;
        18'd64080: out = 16'h40_00;
        18'd64083: out = 16'h80_90;
        18'd64086: out = 16'h40_00;
        18'd64089: out = 16'h80_90;
        18'd64092: out = 16'h40_00;
        18'd64095: out = 16'h80_90;
        18'd64098: out = 16'h40_00;
        18'd64101: out = 16'h80_90;
        18'd64104: out = 16'h40_00;
        18'd64107: out = 16'h80_90;
        18'd64110: out = 16'h40_00;
        18'd64113: out = 16'h80_90;
        18'd64116: out = 16'h40_00;
        18'd64119: out = 16'h80_90;
        18'd64122: out = 16'h40_00;
        18'd64125: out = 16'h80_90;
        18'd64128: out = 16'h40_00;
        18'd64131: out = 16'h80_90;
        18'd64134: out = 16'h40_00;
        18'd64137: out = 16'h80_90;
        18'd64140: out = 16'h40_00;
        18'd64143: out = 16'h80_90;
        18'd64146: out = 16'h40_00;
        18'd64149: out = 16'h80_90;
        18'd64152: out = 16'h40_00;
        18'd64155: out = 16'h80_90;
        18'd64158: out = 16'h40_00;
        18'd64161: out = 16'h80_90;
        18'd64164: out = 16'h40_00;
        18'd64167: out = 16'h80_90;
        18'd64170: out = 16'h40_00;
        18'd64173: out = 16'h80_90;
        18'd64176: out = 16'h40_00;
        18'd64179: out = 16'h80_90;
        18'd64182: out = 16'h40_00;
        18'd64185: out = 16'h80_90;
        18'd64188: out = 16'h40_00;
        18'd64191: out = 16'h80_90;
        18'd64194: out = 16'h40_00;
        18'd64197: out = 16'h80_90;
        18'd64200: out = 16'h40_00;
        18'd64203: out = 16'h80_90;
        18'd64206: out = 16'h40_00;
        18'd64209: out = 16'h80_90;
        18'd64212: out = 16'h40_00;
        18'd64215: out = 16'h80_90;
        18'd64218: out = 16'h40_00;
        18'd64221: out = 16'h80_90;
        18'd64224: out = 16'h40_00;
        18'd64227: out = 16'h80_90;
        18'd64230: out = 16'h40_00;
        18'd64233: out = 16'h80_90;
        18'd64236: out = 16'h40_00;
        18'd64239: out = 16'h80_90;
        18'd64242: out = 16'h40_00;
        18'd64245: out = 16'h80_90;
        18'd64248: out = 16'h40_00;
        18'd64251: out = 16'h80_90;
        18'd64254: out = 16'h40_00;
        18'd64257: out = 16'h80_90;
        18'd64260: out = 16'h40_00;
        18'd64263: out = 16'h80_90;
        18'd64266: out = 16'h40_00;
        18'd64269: out = 16'h80_90;
        18'd64272: out = 16'h40_00;
        18'd64275: out = 16'h80_90;
        18'd64278: out = 16'h40_00;
        18'd64281: out = 16'h80_90;
        18'd64284: out = 16'h40_00;
        18'd64287: out = 16'h80_90;
        18'd64290: out = 16'h40_00;
        18'd64293: out = 16'h80_90;
        18'd64296: out = 16'h40_00;
        18'd64299: out = 16'h80_90;
        18'd64302: out = 16'h40_00;
        18'd64305: out = 16'h80_90;
        18'd64308: out = 16'h40_00;
        18'd64311: out = 16'h80_90;
        18'd64314: out = 16'h40_00;
        18'd64317: out = 16'h80_90;
        18'd64320: out = 16'h40_00;
        18'd64323: out = 16'h80_90;
        18'd64326: out = 16'h40_00;
        18'd64329: out = 16'h80_90;
        18'd64332: out = 16'h40_00;
        18'd64335: out = 16'h80_90;
        18'd64338: out = 16'h40_00;
        18'd64341: out = 16'h80_90;
        18'd64344: out = 16'h40_00;
        18'd64347: out = 16'h80_90;
        18'd64350: out = 16'h40_00;
        18'd64353: out = 16'h80_90;
        18'd64356: out = 16'h40_00;
        18'd64359: out = 16'h80_90;
        18'd64362: out = 16'h40_00;
        18'd64365: out = 16'h80_90;
        18'd64368: out = 16'h40_00;
        18'd64371: out = 16'h80_90;
        18'd64374: out = 16'h40_00;
        18'd64377: out = 16'h80_90;
        18'd64380: out = 16'h40_00;
        18'd64383: out = 16'h80_90;
        18'd64386: out = 16'h40_00;
        18'd64389: out = 16'h80_90;
        18'd64392: out = 16'h40_00;
        18'd64395: out = 16'h80_90;
        18'd64398: out = 16'h40_00;
        18'd64401: out = 16'h80_90;
        18'd64404: out = 16'h40_00;
        18'd64407: out = 16'h80_90;
        18'd64410: out = 16'h40_00;
        18'd64413: out = 16'h80_90;
        18'd64416: out = 16'h40_00;
        18'd64419: out = 16'h80_90;
        18'd64422: out = 16'h40_00;
        18'd64425: out = 16'h80_90;
        18'd64428: out = 16'h40_00;
        18'd64431: out = 16'h80_90;
        18'd64434: out = 16'h40_00;
        18'd64437: out = 16'h80_90;
        18'd64440: out = 16'h40_00;
        18'd64443: out = 16'h80_90;
        18'd64446: out = 16'h40_00;
        18'd64449: out = 16'h80_90;
        18'd64452: out = 16'h40_00;
        18'd64455: out = 16'h80_90;
        18'd64458: out = 16'h40_00;
        18'd64461: out = 16'h80_90;
        18'd64464: out = 16'h40_00;
        18'd64467: out = 16'h80_90;
        18'd64470: out = 16'h40_00;
        18'd64473: out = 16'h80_90;
        18'd64476: out = 16'h40_00;
        18'd64479: out = 16'h80_90;
        18'd64482: out = 16'h40_00;
        18'd64485: out = 16'h80_90;
        18'd64488: out = 16'h40_00;
        18'd64491: out = 16'h80_90;
        18'd64494: out = 16'h40_00;
        18'd64497: out = 16'h80_90;
        18'd64500: out = 16'h40_00;
        18'd64503: out = 16'h80_90;
        18'd64506: out = 16'h40_00;
        18'd64509: out = 16'h80_90;
        18'd64512: out = 16'h40_00;
        18'd64515: out = 16'h80_90;
        18'd64518: out = 16'h40_00;
        18'd64521: out = 16'h80_90;
        18'd64524: out = 16'h40_00;
        18'd64527: out = 16'h80_90;
        18'd64530: out = 16'h40_00;
        18'd64533: out = 16'h80_90;
        18'd64536: out = 16'h40_00;
        18'd64539: out = 16'h80_90;
        18'd64542: out = 16'h40_00;
        18'd64545: out = 16'h80_90;
        18'd64548: out = 16'h40_00;
        18'd64551: out = 16'h80_90;
        18'd64554: out = 16'h40_00;
        18'd64557: out = 16'h80_90;
        18'd64560: out = 16'h40_00;
        18'd64563: out = 16'h80_90;
        18'd64566: out = 16'h40_00;
        18'd64569: out = 16'h80_90;
        18'd64572: out = 16'h40_00;
        18'd64575: out = 16'h80_90;
        18'd64578: out = 16'h40_00;
        18'd64581: out = 16'h80_90;
        18'd64584: out = 16'h40_00;
        18'd64587: out = 16'h80_90;
        18'd64590: out = 16'h40_00;
        18'd64593: out = 16'h80_90;
        18'd64596: out = 16'h40_00;
        18'd64599: out = 16'h80_90;
        18'd64602: out = 16'h40_00;
        18'd64605: out = 16'h80_90;
        18'd64608: out = 16'h40_00;
        18'd64611: out = 16'h80_90;
        18'd64614: out = 16'h40_00;
        18'd64617: out = 16'h80_90;
        18'd64620: out = 16'h40_00;
        18'd64623: out = 16'h80_90;
        18'd64626: out = 16'h40_00;
        18'd64629: out = 16'h80_90;
        18'd64632: out = 16'h40_00;
        18'd64635: out = 16'h80_90;
        18'd64638: out = 16'h40_00;
        18'd64641: out = 16'h80_90;
        18'd64644: out = 16'h40_00;
        18'd64647: out = 16'h80_90;
        18'd64650: out = 16'h40_00;
        18'd64653: out = 16'h80_90;
        18'd64656: out = 16'h40_00;
        18'd64659: out = 16'h80_90;
        18'd64662: out = 16'h40_00;
        18'd64665: out = 16'h80_90;
        18'd64668: out = 16'h40_00;
        18'd64671: out = 16'h80_90;
        18'd64674: out = 16'h40_00;
        18'd64677: out = 16'h80_90;
        18'd64680: out = 16'h40_00;
        18'd64683: out = 16'h80_90;
        18'd64686: out = 16'h40_00;
        18'd64689: out = 16'h80_90;
        18'd64692: out = 16'h40_00;
        18'd64695: out = 16'h80_90;
        18'd64698: out = 16'h40_00;
        18'd64701: out = 16'h80_90;
        18'd64704: out = 16'h40_00;
        18'd64707: out = 16'h80_90;
        18'd64710: out = 16'h40_00;
        18'd64713: out = 16'h80_90;
        18'd64716: out = 16'h40_00;
        18'd64719: out = 16'h80_90;
        18'd64722: out = 16'h40_00;
        18'd64725: out = 16'h80_90;
        18'd64728: out = 16'h40_00;
        18'd64731: out = 16'h80_90;
        18'd64734: out = 16'h40_00;
        18'd64737: out = 16'h80_90;
        18'd64740: out = 16'h40_00;
        18'd64743: out = 16'h80_90;
        18'd64746: out = 16'h40_00;
        18'd64749: out = 16'h80_90;
        18'd64752: out = 16'h40_00;
        18'd64755: out = 16'h80_90;
        18'd64758: out = 16'h40_00;
        18'd64761: out = 16'h80_90;
        18'd64764: out = 16'h40_00;
        18'd64767: out = 16'h80_90;
        18'd64770: out = 16'h40_00;
        18'd64773: out = 16'h80_90;
        18'd64776: out = 16'h40_00;
        18'd64779: out = 16'h80_90;
        18'd64782: out = 16'h40_00;
        18'd64785: out = 16'h80_90;
        18'd64788: out = 16'h40_00;
        18'd64791: out = 16'h80_90;
        18'd64794: out = 16'h40_00;
        18'd64797: out = 16'h80_90;
        18'd64800: out = 16'h40_00;
        18'd64803: out = 16'h80_90;
        18'd64806: out = 16'h40_00;
        18'd64809: out = 16'h80_90;
        18'd64812: out = 16'h40_00;
        18'd64815: out = 16'h80_90;
        18'd64818: out = 16'h40_00;
        18'd64821: out = 16'h80_90;
        18'd64824: out = 16'h40_00;
        18'd64827: out = 16'h80_90;
        18'd64830: out = 16'h40_00;
        18'd64833: out = 16'h80_90;
        18'd64836: out = 16'h40_00;
        18'd64839: out = 16'h80_90;
        18'd64842: out = 16'h40_00;
        18'd64845: out = 16'h80_90;
        18'd64848: out = 16'h40_00;
        18'd64851: out = 16'h80_90;
        18'd64854: out = 16'h40_00;
        18'd64857: out = 16'h80_90;
        18'd64860: out = 16'h40_00;
        18'd64863: out = 16'h80_90;
        18'd64866: out = 16'h40_00;
        18'd64869: out = 16'h80_90;
        18'd64872: out = 16'h40_00;
        18'd64875: out = 16'h80_90;
        18'd64878: out = 16'h40_00;
        18'd64881: out = 16'h80_90;
        18'd64884: out = 16'h40_00;
        18'd64887: out = 16'h80_90;
        18'd64890: out = 16'h40_00;
        18'd64893: out = 16'h80_90;
        18'd64896: out = 16'h40_00;
        18'd64899: out = 16'h80_90;
        18'd64902: out = 16'h40_00;
        18'd64905: out = 16'h80_90;
        18'd64908: out = 16'h40_00;
        18'd64911: out = 16'h80_90;
        18'd64914: out = 16'h40_00;
        18'd64917: out = 16'h80_90;
        18'd64920: out = 16'h40_00;
        18'd64923: out = 16'h80_90;
        18'd64926: out = 16'h40_00;
        18'd64929: out = 16'h80_90;
        18'd64932: out = 16'h40_00;
        18'd64935: out = 16'h80_90;
        18'd64938: out = 16'h40_00;
        18'd64941: out = 16'h80_90;
        18'd64944: out = 16'h40_00;
        18'd64947: out = 16'h80_90;
        18'd64950: out = 16'h40_00;
        18'd64953: out = 16'h80_90;
        18'd64956: out = 16'h40_00;
        18'd64959: out = 16'h80_90;
        18'd64962: out = 16'h40_00;
        18'd64965: out = 16'h80_90;
        18'd64968: out = 16'h40_00;
        18'd64971: out = 16'h80_90;
        18'd64974: out = 16'h40_00;
        18'd64977: out = 16'h80_90;
        18'd64980: out = 16'h40_00;
        18'd64983: out = 16'h80_90;
        18'd64986: out = 16'h40_00;
        18'd64989: out = 16'h80_90;
        18'd64992: out = 16'h40_00;
        18'd64995: out = 16'h80_90;
        18'd64998: out = 16'h40_00;
        18'd65001: out = 16'h80_90;
        18'd65004: out = 16'h40_00;
        18'd65007: out = 16'h80_90;
        18'd65010: out = 16'h40_00;
        18'd65013: out = 16'h80_90;
        18'd65016: out = 16'h40_00;
        18'd65019: out = 16'h80_90;
        18'd65022: out = 16'h40_00;
        18'd65025: out = 16'h80_90;
        18'd65028: out = 16'h40_00;
        18'd65031: out = 16'h80_90;
        18'd65034: out = 16'h40_00;
        18'd65037: out = 16'h80_90;
        18'd65040: out = 16'h40_00;
        18'd65043: out = 16'h80_90;
        18'd65046: out = 16'h40_00;
        18'd65049: out = 16'h80_90;
        18'd65052: out = 16'h40_00;
        18'd65055: out = 16'h80_90;
        18'd65058: out = 16'h40_00;
        18'd65061: out = 16'h80_90;
        18'd65064: out = 16'h40_00;
        18'd65067: out = 16'h80_90;
        18'd65070: out = 16'h40_00;
        18'd65073: out = 16'h80_90;
        18'd65076: out = 16'h40_00;
        18'd65079: out = 16'h80_90;
        18'd65082: out = 16'h40_00;
        18'd65085: out = 16'h80_90;
        18'd65088: out = 16'h40_00;
        18'd65091: out = 16'h80_90;
        18'd65094: out = 16'h40_00;
        18'd65097: out = 16'h80_90;
        18'd65100: out = 16'h40_00;
        18'd65103: out = 16'h80_90;
        18'd65106: out = 16'h40_00;
        18'd65109: out = 16'h80_90;
        18'd65112: out = 16'h40_00;
        18'd65115: out = 16'h80_90;
        18'd65118: out = 16'h40_00;
        18'd65121: out = 16'h80_90;
        18'd65124: out = 16'h40_00;
        18'd65127: out = 16'h80_90;
        18'd65130: out = 16'h40_00;
        18'd65133: out = 16'h80_90;
        18'd65136: out = 16'h40_00;
        18'd65139: out = 16'h80_90;
        18'd65142: out = 16'h40_00;
        18'd65145: out = 16'h80_90;
        18'd65148: out = 16'h40_00;
        18'd65151: out = 16'h80_90;
        18'd65154: out = 16'h40_00;
        18'd65157: out = 16'h80_90;
        18'd65160: out = 16'h40_00;
        18'd65163: out = 16'h80_90;
        18'd65166: out = 16'h40_00;
        18'd65169: out = 16'h80_90;
        18'd65172: out = 16'h40_00;
        18'd65175: out = 16'h80_90;
        18'd65178: out = 16'h40_00;
        18'd65181: out = 16'h80_90;
        18'd65184: out = 16'h40_00;
        18'd65187: out = 16'h80_90;
        18'd65190: out = 16'h40_00;
        18'd65193: out = 16'h80_90;
        18'd65196: out = 16'h40_00;
        18'd65199: out = 16'h80_90;
        18'd65202: out = 16'h40_00;
        18'd65205: out = 16'h80_90;
        18'd65208: out = 16'h40_00;
        18'd65211: out = 16'h80_90;
        18'd65214: out = 16'h40_00;
        18'd65217: out = 16'h80_90;
        18'd65220: out = 16'h40_00;
        18'd65223: out = 16'h80_90;
        18'd65226: out = 16'h40_00;
        18'd65229: out = 16'h80_90;
        18'd65232: out = 16'h40_00;
        18'd65235: out = 16'h80_90;
        18'd65238: out = 16'h40_00;
        18'd65241: out = 16'h80_90;
        18'd65244: out = 16'h40_00;
        18'd65247: out = 16'h80_90;
        18'd65250: out = 16'h40_00;
        18'd65253: out = 16'h80_90;
        18'd65256: out = 16'h40_00;
        18'd65259: out = 16'h80_90;
        18'd65262: out = 16'h40_00;
        18'd65265: out = 16'h80_90;
        18'd65268: out = 16'h40_00;
        18'd65271: out = 16'h80_90;
        18'd65274: out = 16'h40_00;
        18'd65277: out = 16'h80_90;
        18'd65280: out = 16'h40_00;
        18'd65283: out = 16'h80_90;
        18'd65286: out = 16'h40_00;
        18'd65289: out = 16'h80_40;
        18'd65292: out = 16'h40_00;
        18'd65295: out = 16'h00_00;
        18'd65298: out = 16'h80_99;
        18'd65301: out = 16'h00_90;
        18'd65304: out = 16'h80_9A;
        18'd65307: out = 16'h00_01;
        18'd65310: out = 16'h80_9B;
        18'd65313: out = 16'h00_F0;
        18'd65316: out = 16'h80_9C;
        18'd65319: out = 16'h00_00;
        18'd65322: out = 16'h80_9D;
        18'd65325: out = 16'h00_32;
        18'd65328: out = 16'h80_63;
        18'd65331: out = 16'h00_1F;
        18'd65334: out = 16'h80_64;
        18'd65337: out = 16'h00_00;
        18'd65340: out = 16'h80_65;
        18'd65343: out = 16'h00_1F;
        18'd65346: out = 16'h80_90;
        18'd65349: out = 16'h00_60;
        18'd65352: out = 16'h80_90;
        18'd65355: out = 16'h40_00;
        18'd65358: out = 16'h80_90;
        18'd65361: out = 16'h40_00;
        18'd65364: out = 16'h80_90;
        18'd65367: out = 16'h40_00;
        18'd65370: out = 16'h80_90;
        18'd65373: out = 16'h40_00;
        18'd65376: out = 16'h80_90;
        18'd65379: out = 16'h40_00;
        18'd65382: out = 16'h80_90;
        18'd65385: out = 16'h40_00;
        18'd65388: out = 16'h80_90;
        18'd65391: out = 16'h40_00;
        18'd65394: out = 16'h80_90;
        18'd65397: out = 16'h40_00;
        18'd65400: out = 16'h80_90;
        18'd65403: out = 16'h40_00;
        18'd65406: out = 16'h80_90;
        18'd65409: out = 16'h40_00;
        18'd65412: out = 16'h80_90;
        18'd65415: out = 16'h40_00;
        18'd65418: out = 16'h80_90;
        18'd65421: out = 16'h40_00;
        18'd65424: out = 16'h80_90;
        18'd65427: out = 16'h40_00;
        18'd65430: out = 16'h80_90;
        18'd65433: out = 16'h40_00;
        18'd65436: out = 16'h80_90;
        18'd65439: out = 16'h40_00;
        18'd65442: out = 16'h80_90;
        18'd65445: out = 16'h40_00;
        18'd65448: out = 16'h80_90;
        18'd65451: out = 16'h40_00;
        18'd65454: out = 16'h80_90;
        18'd65457: out = 16'h40_00;
        18'd65460: out = 16'h80_90;
        18'd65463: out = 16'h40_00;
        18'd65466: out = 16'h80_90;
        18'd65469: out = 16'h40_00;
        18'd65472: out = 16'h80_90;
        18'd65475: out = 16'h40_00;
        18'd65478: out = 16'h80_90;
        18'd65481: out = 16'h40_00;
        18'd65484: out = 16'h80_90;
        18'd65487: out = 16'h40_00;
        18'd65490: out = 16'h80_90;
        18'd65493: out = 16'h40_00;
        18'd65496: out = 16'h80_90;
        18'd65499: out = 16'h40_00;
        18'd65502: out = 16'h80_90;
        18'd65505: out = 16'h40_00;
        18'd65508: out = 16'h80_90;
        18'd65511: out = 16'h40_00;
        18'd65514: out = 16'h80_90;
        18'd65517: out = 16'h40_00;
        18'd65520: out = 16'h80_90;
        18'd65523: out = 16'h40_00;
        18'd65526: out = 16'h80_90;
        18'd65529: out = 16'h40_00;
        18'd65532: out = 16'h80_90;
        18'd65535: out = 16'h40_00;
        18'd65538: out = 16'h80_90;
        18'd65541: out = 16'h40_00;
        18'd65544: out = 16'h80_90;
        18'd65547: out = 16'h40_00;
        18'd65550: out = 16'h80_90;
        18'd65553: out = 16'h40_00;
        18'd65556: out = 16'h80_90;
        18'd65559: out = 16'h40_00;
        18'd65562: out = 16'h80_90;
        18'd65565: out = 16'h40_00;
        18'd65568: out = 16'h80_90;
        18'd65571: out = 16'h40_00;
        18'd65574: out = 16'h80_90;
        18'd65577: out = 16'h40_00;
        18'd65580: out = 16'h80_90;
        18'd65583: out = 16'h40_00;
        18'd65586: out = 16'h80_90;
        18'd65589: out = 16'h40_00;
        18'd65592: out = 16'h80_90;
        18'd65595: out = 16'h40_00;
        18'd65598: out = 16'h80_90;
        18'd65601: out = 16'h40_00;
        18'd65604: out = 16'h80_90;
        18'd65607: out = 16'h40_00;
        18'd65610: out = 16'h80_90;
        18'd65613: out = 16'h40_00;
        18'd65616: out = 16'h80_90;
        18'd65619: out = 16'h40_00;
        18'd65622: out = 16'h80_90;
        18'd65625: out = 16'h40_00;
        18'd65628: out = 16'h80_90;
        18'd65631: out = 16'h40_00;
        18'd65634: out = 16'h80_90;
        18'd65637: out = 16'h40_00;
        18'd65640: out = 16'h80_90;
        18'd65643: out = 16'h40_00;
        18'd65646: out = 16'h80_90;
        18'd65649: out = 16'h40_00;
        18'd65652: out = 16'h80_90;
        18'd65655: out = 16'h40_00;
        18'd65658: out = 16'h80_90;
        18'd65661: out = 16'h40_00;
        18'd65664: out = 16'h80_90;
        18'd65667: out = 16'h40_00;
        18'd65670: out = 16'h80_90;
        18'd65673: out = 16'h40_00;
        18'd65676: out = 16'h80_90;
        18'd65679: out = 16'h40_00;
        18'd65682: out = 16'h80_90;
        18'd65685: out = 16'h40_00;
        18'd65688: out = 16'h80_90;
        18'd65691: out = 16'h40_00;
        18'd65694: out = 16'h80_90;
        18'd65697: out = 16'h40_00;
        18'd65700: out = 16'h80_90;
        18'd65703: out = 16'h40_00;
        18'd65706: out = 16'h80_90;
        18'd65709: out = 16'h40_00;



        default: begin
            delay = 1;
            out = 0;
        end 
    endcase
  end
endmodule