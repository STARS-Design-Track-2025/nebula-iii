`timescale 1ns / 1ps
module request_unit_tb;
logic clk, rst, i_ack, d_ack, freeze;
logic [31:0] PC, mem_address,

















endmodule