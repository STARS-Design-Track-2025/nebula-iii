* NGSPICE file created from team_08.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_16 abstract view
.subckt sky130_fd_sc_hd__clkinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_1 abstract view
.subckt sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_2 abstract view
.subckt sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

.subckt team_08 ACK_I ADR_O[0] ADR_O[10] ADR_O[11] ADR_O[12] ADR_O[13] ADR_O[14] ADR_O[15]
+ ADR_O[16] ADR_O[17] ADR_O[18] ADR_O[19] ADR_O[1] ADR_O[20] ADR_O[21] ADR_O[22] ADR_O[23]
+ ADR_O[24] ADR_O[25] ADR_O[26] ADR_O[27] ADR_O[28] ADR_O[29] ADR_O[2] ADR_O[30] ADR_O[31]
+ ADR_O[3] ADR_O[4] ADR_O[5] ADR_O[6] ADR_O[7] ADR_O[8] ADR_O[9] CYC_O DAT_I[0] DAT_I[10]
+ DAT_I[11] DAT_I[12] DAT_I[13] DAT_I[14] DAT_I[15] DAT_I[16] DAT_I[17] DAT_I[18]
+ DAT_I[19] DAT_I[1] DAT_I[20] DAT_I[21] DAT_I[22] DAT_I[23] DAT_I[24] DAT_I[25] DAT_I[26]
+ DAT_I[27] DAT_I[28] DAT_I[29] DAT_I[2] DAT_I[30] DAT_I[31] DAT_I[3] DAT_I[4] DAT_I[5]
+ DAT_I[6] DAT_I[7] DAT_I[8] DAT_I[9] DAT_O[0] DAT_O[10] DAT_O[11] DAT_O[12] DAT_O[13]
+ DAT_O[14] DAT_O[15] DAT_O[16] DAT_O[17] DAT_O[18] DAT_O[19] DAT_O[1] DAT_O[20] DAT_O[21]
+ DAT_O[22] DAT_O[23] DAT_O[24] DAT_O[25] DAT_O[26] DAT_O[27] DAT_O[28] DAT_O[29]
+ DAT_O[2] DAT_O[30] DAT_O[31] DAT_O[3] DAT_O[4] DAT_O[5] DAT_O[6] DAT_O[7] DAT_O[8]
+ DAT_O[9] SEL_O[0] SEL_O[1] SEL_O[2] SEL_O[3] STB_O WE_O clk en gpio_in[0] gpio_in[10]
+ gpio_in[11] gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17]
+ gpio_in[18] gpio_in[19] gpio_in[1] gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23]
+ gpio_in[24] gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2]
+ gpio_in[30] gpio_in[31] gpio_in[32] gpio_in[33] gpio_in[3] gpio_in[4] gpio_in[5]
+ gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9] gpio_oeb[0] gpio_oeb[10] gpio_oeb[11]
+ gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15] gpio_oeb[16] gpio_oeb[17] gpio_oeb[18]
+ gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21] gpio_oeb[22] gpio_oeb[23] gpio_oeb[24]
+ gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28] gpio_oeb[29] gpio_oeb[2] gpio_oeb[30]
+ gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[3] gpio_oeb[4] gpio_oeb[5] gpio_oeb[6]
+ gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12]
+ gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19]
+ gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25]
+ gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31]
+ gpio_out[32] gpio_out[33] gpio_out[3] gpio_out[4] gpio_out[5] gpio_out[6] gpio_out[7]
+ gpio_out[8] gpio_out[9] nrst vccd1 vssd1
XFILLER_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09523__A2 net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11866__A0 _05771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09671_ top.CPU.registers.data\[57\] top.CPU.registers.data\[25\] net837 vssd1 vssd1
+ vccd1 vccd1 _05310_ sky130_fd_sc_hd__mux2_1
XANTENNA__11330__A2 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08622_ top.CPU.registers.data\[558\] top.CPU.registers.data\[526\] net819 vssd1
+ vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__mux2_1
X_13882__52 clknet_leaf_161_clk vssd1 vssd1 vccd1 vccd1 net1521 sky130_fd_sc_hd__inv_2
XFILLER_54_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10958__B net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11618__A0 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08553_ _04158_ _04190_ vssd1 vssd1 vccd1 vccd1 _04192_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout162_A _06760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08484_ top.CPU.control_unit.instruction\[17\] _03160_ _03985_ vssd1 vssd1 vccd1
+ vccd1 _04123_ sky130_fd_sc_hd__o21a_2
XANTENNA__08495__C1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09039__A1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1071_A net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12892__C _07322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout427_A _06756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1169_A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07759__S net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09105_ net712 _04742_ _04743_ vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__or3_1
XANTENNA__13791__B1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout215_X net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1336_A net1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09036_ top.CPU.registers.data\[968\] net1314 net845 top.CPU.registers.data\[1000\]
+ net716 vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__a221o_1
XFILLER_164_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout796_A net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13543__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14352__522 clknet_leaf_200_clk vssd1 vssd1 vccd1 vccd1 net1991 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_57_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold340 top.CPU.registers.data\[686\] vssd1 vssd1 vccd1 vccd1 net2897 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold351 top.CPU.registers.data\[309\] vssd1 vssd1 vccd1 vccd1 net2908 sky130_fd_sc_hd__dlygate4sd3_1
X_14649__819 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 net2288 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_92_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold362 top.CPU.handler.toreg\[30\] vssd1 vssd1 vccd1 vccd1 net2919 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold373 top.CPU.registers.data\[513\] vssd1 vssd1 vccd1 vccd1 net2930 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold384 top.CPU.registers.data\[786\] vssd1 vssd1 vccd1 vccd1 net2941 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold395 _02599_ vssd1 vssd1 vccd1 vccd1 net2952 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout820 net822 vssd1 vssd1 vccd1 vccd1 net820 sky130_fd_sc_hd__clkbuf_4
XFILLER_117_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout831 net839 vssd1 vssd1 vccd1 vccd1 net831 sky130_fd_sc_hd__buf_4
X_09938_ _04193_ _05576_ vssd1 vssd1 vccd1 vccd1 _05577_ sky130_fd_sc_hd__or2_1
Xfanout842 net843 vssd1 vssd1 vccd1 vccd1 net842 sky130_fd_sc_hd__clkbuf_4
Xfanout853 net854 vssd1 vssd1 vccd1 vccd1 net853 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_70_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout864 net870 vssd1 vssd1 vccd1 vccd1 net864 sky130_fd_sc_hd__clkbuf_4
Xfanout875 net876 vssd1 vssd1 vccd1 vccd1 net875 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_70_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout886 net887 vssd1 vssd1 vccd1 vccd1 net886 sky130_fd_sc_hd__buf_2
XANTENNA__11029__B net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11857__B1 net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09869_ _05432_ _05502_ _05504_ _05507_ _05434_ vssd1 vssd1 vccd1 vccd1 _05508_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout751_X net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1040 top.CPU.registers.data\[847\] vssd1 vssd1 vccd1 vccd1 net3597 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08722__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11321__A2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1051 top.CPU.registers.data\[622\] vssd1 vssd1 vccd1 vccd1 net3608 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13525__A _03783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11900_ net457 _06601_ vssd1 vssd1 vccd1 vccd1 _06770_ sky130_fd_sc_hd__nor2_2
Xhold1062 top.CPU.registers.data\[509\] vssd1 vssd1 vccd1 vccd1 net3619 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10501__X _06126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12880_ top.CPU.alu.program_counter\[24\] _03646_ vssd1 vssd1 vccd1 vccd1 _07326_
+ sky130_fd_sc_hd__and2_1
Xhold1073 top.CPU.registers.data\[101\] vssd1 vssd1 vccd1 vccd1 net3630 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08619__A _04225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1084 net97 vssd1 vssd1 vccd1 vccd1 net3641 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1095 top.CPU.registers.data\[652\] vssd1 vssd1 vccd1 vccd1 net3652 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11609__A0 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10868__B _06467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11831_ net1404 net540 _06754_ vssd1 vssd1 vccd1 vccd1 _06766_ sky130_fd_sc_hd__or3_1
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11762_ net469 _06605_ net241 net163 net3395 vssd1 vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__a32o_1
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13501_ top.CPU.data_out\[9\] net587 _02969_ _02970_ vssd1 vssd1 vccd1 vccd1 _02507_
+ sky130_fd_sc_hd__o22a_1
X_10713_ _04859_ _05275_ _05541_ vssd1 vssd1 vccd1 vccd1 _06328_ sky130_fd_sc_hd__a21oi_1
X_11693_ _06521_ net208 net167 net3013 vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__a22o_1
X_16220_ net2554 _02430_ net1194 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[1020\]
+ sky130_fd_sc_hd__dfrtp_1
X_13432_ net3627 _02867_ net121 vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__mux2_1
XANTENNA__12034__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10644_ _06217_ _06261_ net306 vssd1 vssd1 vccd1 vccd1 _06262_ sky130_fd_sc_hd__mux2_1
XFILLER_167_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11388__A2 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13960__130 clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 net1599 sky130_fd_sc_hd__inv_2
X_16151_ net2485 _02361_ net1180 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[951\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10575_ net408 _06023_ vssd1 vssd1 vccd1 vccd1 _06196_ sky130_fd_sc_hd__nand2_1
X_13363_ top.I2C.data_out\[15\] net554 _02890_ net597 vssd1 vssd1 vccd1 vccd1 _02891_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09450__A1 _05087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15102_ net1484 _01315_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r2_prev\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_12314_ net2605 _05498_ net1253 vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__mux2_1
XFILLER_5_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16082_ net2416 _02292_ net1101 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[882\]
+ sky130_fd_sc_hd__dfrtp_1
X_14903__1073 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 net2542 sky130_fd_sc_hd__inv_2
X_13294_ top.mmio.mem_data_i\[21\] top.mmio.mem_data_i\[20\] top.mmio.mem_data_i\[23\]
+ top.mmio.mem_data_i\[22\] vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__and4b_1
XFILLER_170_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12337__A1 _05018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15033_ clknet_leaf_91_clk _01278_ net1270 vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__dfrtp_1
XFILLER_114_219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14095__265 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 net1734 sky130_fd_sc_hd__inv_2
XANTENNA__09202__A1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12245_ net2921 _05934_ net434 vssd1 vssd1 vccd1 vccd1 _01435_ sky130_fd_sc_hd__mux2_1
X_12176_ top.CPU.registers.data\[64\] net172 vssd1 vssd1 vccd1 vccd1 _06856_ sky130_fd_sc_hd__and2_1
XFILLER_150_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07764__A1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11560__A2 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11127_ net481 net458 _06621_ net301 net3528 vssd1 vssd1 vccd1 vccd1 _02289_ sky130_fd_sc_hd__a32o_1
XANTENNA__10124__A _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09913__A net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14831__1001 clknet_leaf_179_clk vssd1 vssd1 vccd1 vccd1 net2470 sky130_fd_sc_hd__inv_2
XANTENNA__11848__B1 net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15935_ net2269 _02145_ net1221 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[735\]
+ sky130_fd_sc_hd__dfrtp_1
X_11058_ net325 net140 net536 net367 net2808 vssd1 vssd1 vccd1 vccd1 _02323_ sky130_fd_sc_hd__a32o_1
XFILLER_77_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09505__A2 net1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09061__S0 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11312__A2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10009_ _03683_ _03755_ net375 vssd1 vssd1 vccd1 vccd1 _05648_ sky130_fd_sc_hd__mux2_1
XFILLER_77_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15866_ net2200 _02076_ net1250 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[666\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10520__B1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15797_ net2131 _02007_ net1211 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[597\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_91_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11076__B2 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10780__C_N net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14793__963 clknet_leaf_184_clk vssd1 vssd1 vccd1 vccd1 net2432 sky130_fd_sc_hd__inv_2
XANTENNA__10794__A net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08492__A2 net1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16418_ clknet_leaf_55_clk net2595 net1142 vssd1 vssd1 vccd1 vccd1 top.I2C.I2C_state\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_165_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08229__C1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11379__A2 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16349_ clknet_leaf_68_clk _02558_ net1167 vssd1 vssd1 vccd1 vccd1 top.CPU.addressnew\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_146_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14336__506 clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 net1975 sky130_fd_sc_hd__inv_2
XFILLER_8_170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11000__B2 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12233__B net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout127 net129 vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__buf_2
Xfanout138 _05692_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__buf_2
XFILLER_86_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout149 _06412_ vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__clkbuf_2
X_07984_ top.CPU.registers.data\[760\] net1378 net983 top.CPU.registers.data\[728\]
+ net907 vssd1 vssd1 vccd1 vccd1 _03623_ sky130_fd_sc_hd__a221o_1
XFILLER_101_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13828__B2 top.CPU.data_out\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09382__X _05021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09723_ top.CPU.control_unit.instruction\[25\] net1046 net899 vssd1 vssd1 vccd1 vccd1
+ _05362_ sky130_fd_sc_hd__o21a_1
XANTENNA__11839__B1 net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10969__A net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11303__A2 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout377_A net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08704__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13345__A _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09654_ _04125_ _05291_ vssd1 vssd1 vccd1 vccd1 _05293_ sky130_fd_sc_hd__and2b_1
XANTENNA__08439__A net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08605_ top.CPU.registers.data\[943\] top.CPU.registers.data\[911\] top.CPU.registers.data\[815\]
+ top.CPU.registers.data\[783\] net974 net1281 vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__mux4_1
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09585_ net673 _05223_ _05222_ net928 vssd1 vssd1 vccd1 vccd1 _05224_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout544_A _06523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout165_X net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1286_A net1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11067__A1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08468__C1 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08536_ net933 _04160_ _04161_ net953 vssd1 vssd1 vccd1 vccd1 _04175_ sky130_fd_sc_hd__o211a_1
XFILLER_23_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12803__A2 _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10814__A1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout332_X net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout711_A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08467_ top.CPU.registers.data\[593\] net1296 net1016 top.CPU.registers.data\[625\]
+ net938 vssd1 vssd1 vccd1 vccd1 _04106_ sky130_fd_sc_hd__a221o_1
X_13944__114 clknet_leaf_169_clk vssd1 vssd1 vccd1 vccd1 net1583 sky130_fd_sc_hd__inv_2
XANTENNA_fanout809_A net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1074_X net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08398_ top.CPU.registers.data\[850\] net1287 net1006 top.CPU.registers.data\[882\]
+ net930 vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__a221o_1
XFILLER_11_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_93_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08235__A2 net1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10042__A2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10360_ net1406 net577 net518 net133 vssd1 vssd1 vccd1 vccd1 _05991_ sky130_fd_sc_hd__and4_1
X_14079__249 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 net1718 sky130_fd_sc_hd__inv_2
XFILLER_136_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12319__A1 _03783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout799_X net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11790__A2 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09019_ top.CPU.registers.data_out_r2_prev\[9\] net685 _04657_ vssd1 vssd1 vccd1
+ vccd1 _04658_ sky130_fd_sc_hd__o21ai_2
X_10291_ _05780_ _05788_ net387 vssd1 vssd1 vccd1 vccd1 _05924_ sky130_fd_sc_hd__mux2_1
XANTENNA__10643__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08180__Y _03819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12030_ net141 net3282 net150 vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10870__C net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold170 top.CPU.registers.data\[399\] vssd1 vssd1 vccd1 vccd1 net2727 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 top.CPU.registers.data\[257\] vssd1 vssd1 vccd1 vccd1 net2738 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 net81 vssd1 vssd1 vccd1 vccd1 net2749 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_151_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout966_X net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11542__A2 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_31_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout650 net658 vssd1 vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__clkbuf_4
Xfanout661 net662 vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__clkbuf_8
Xfanout672 net673 vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__clkbuf_4
Xfanout683 net684 vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__buf_4
XANTENNA__10879__A net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout694 net701 vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__clkbuf_4
X_15720_ net2054 _01930_ net1099 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[520\]
+ sky130_fd_sc_hd__dfrtp_1
X_12932_ _07365_ _07373_ net129 vssd1 vssd1 vccd1 vccd1 _07374_ sky130_fd_sc_hd__mux2_1
XFILLER_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_166_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08171__A1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15651_ net1985 _01861_ net1206 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[451\]
+ sky130_fd_sc_hd__dfrtp_1
X_12863_ _07307_ _07309_ vssd1 vssd1 vccd1 vccd1 _07311_ sky130_fd_sc_hd__nor2_1
X_14480__650 clknet_leaf_198_clk vssd1 vssd1 vccd1 vccd1 net2119 sky130_fd_sc_hd__inv_2
XFILLER_74_887 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_46_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08068__B net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11058__A1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14777__947 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 net2416 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_87_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11814_ net571 _06654_ net236 _06765_ vssd1 vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__a31o_1
XANTENNA__13598__A3 _06081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11206__C net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08459__C1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15582_ net1916 _01792_ net1201 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[382\]
+ sky130_fd_sc_hd__dfrtp_1
X_12794_ top.CPU.alu.program_counter\[15\] _07240_ vssd1 vssd1 vccd1 vccd1 _07249_
+ sky130_fd_sc_hd__xor2_1
XFILLER_57_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_164_Left_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09120__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11745_ _06587_ net498 net192 net2727 vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__a22o_1
XFILLER_18_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14521__691 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 net2160 sky130_fd_sc_hd__inv_2
XANTENNA__11503__A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12007__B1 net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07700__B _03331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14818__988 clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 net2457 sky130_fd_sc_hd__inv_2
X_11676_ net461 _06493_ net236 net165 net3620 vssd1 vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__a32o_1
XFILLER_128_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16203_ net2537 _02413_ net1057 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[1003\]
+ sky130_fd_sc_hd__dfrtp_1
X_13415_ net890 _02928_ vssd1 vssd1 vccd1 vccd1 _02929_ sky130_fd_sc_hd__and2_1
XFILLER_146_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11222__B net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10627_ net406 _06071_ _06245_ net415 vssd1 vssd1 vccd1 vccd1 _06246_ sky130_fd_sc_hd__a211o_1
XANTENNA__10119__A net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08226__A2 net1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_104_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16134_ net2468 _02344_ net1080 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[934\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_155_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13346_ net1402 _02878_ net667 vssd1 vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__mux2_1
X_10558_ _05999_ _06179_ net403 vssd1 vssd1 vccd1 vccd1 _06180_ sky130_fd_sc_hd__mux2_1
XFILLER_142_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11781__A2 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16065_ net2399 _02275_ net1243 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[865\]
+ sky130_fd_sc_hd__dfrtp_1
X_13277_ _03101_ _03137_ _07060_ _07061_ vssd1 vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__a31o_1
XFILLER_170_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10489_ _05913_ _06113_ net405 vssd1 vssd1 vccd1 vccd1 _06114_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_149_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_173_Left_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15016_ clknet_leaf_93_clk _01261_ net1268 vssd1 vssd1 vccd1 vccd1 top.SPI.parameters\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09119__S net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12228_ net3695 net645 _06880_ vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__o21a_1
XFILLER_64_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_119_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12159_ net3777 net172 _06847_ vssd1 vssd1 vccd1 vccd1 _01483_ sky130_fd_sc_hd__a21o_1
XANTENNA__12988__B _06945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08698__C1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15918_ net2252 _02128_ net1106 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[718\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_83_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11297__B2 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08162__A1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11836__A3 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16249__Q top.CPU.control_unit.instruction\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_92_662 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15849_ net2183 _02059_ net1060 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[649\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_80_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13852__22 clknet_leaf_138_clk vssd1 vssd1 vccd1 vccd1 net1491 sky130_fd_sc_hd__inv_2
XFILLER_52_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10301__B _05933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09370_ net956 _05008_ _05007_ net613 vssd1 vssd1 vccd1 vccd1 _05009_ sky130_fd_sc_hd__a211o_1
XANTENNA__11116__C net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09111__B1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08321_ top.CPU.registers.data\[947\] top.CPU.registers.data\[915\] top.CPU.registers.data\[819\]
+ top.CPU.registers.data\[787\] net989 net914 vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__mux4_1
XANTENNA__08465__A2 net1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08252_ top.CPU.registers.data\[406\] net1300 net1021 top.CPU.registers.data\[438\]
+ net917 vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__a221o_1
XANTENNA__10955__C _05808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10526__C_N net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08183_ net1035 _03819_ _03821_ vssd1 vssd1 vccd1 vccd1 _03822_ sky130_fd_sc_hd__a21oi_4
XANTENNA__11132__B net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15290__RESET_B net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_08_1450 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] team_08_1450/LO sky130_fd_sc_hd__conb_1
XANTENNA__12943__S net1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09414__A1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_12_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_12_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout125_A net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_08_1461 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] team_08_1461/LO sky130_fd_sc_hd__conb_1
XANTENNA__11221__B2 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10971__B _06010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11772__A2 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1034_A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09029__S net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07728__A1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout494_A net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11524__A2 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12531__X _07040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout661_A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout282_X net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07967_ net706 _03600_ _03601_ net720 vssd1 vssd1 vccd1 vccd1 _03606_ sky130_fd_sc_hd__o211a_1
XFILLER_102_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13277__A2 _03137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout759_A net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09706_ top.CPU.registers.data\[185\] net1384 net1001 top.CPU.registers.data\[153\]
+ net682 vssd1 vssd1 vccd1 vccd1 _05345_ sky130_fd_sc_hd__a221o_1
XFILLER_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14464__634 clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 net2103 sky130_fd_sc_hd__inv_2
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07898_ net801 _03532_ _03533_ net730 vssd1 vssd1 vccd1 vccd1 _03537_ sky130_fd_sc_hd__o211a_1
X_09637_ _04862_ _04923_ _05274_ _04859_ _04796_ vssd1 vssd1 vccd1 vccd1 _05276_ sky130_fd_sc_hd__o311a_1
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14902__1072 clknet_leaf_182_clk vssd1 vssd1 vccd1 vccd1 net2541 sky130_fd_sc_hd__inv_2
XANTENNA_fanout926_A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1191_X net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1289_X net1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14505__675 clknet_leaf_157_clk vssd1 vssd1 vccd1 vccd1 net2144 sky130_fd_sc_hd__inv_2
X_09568_ net673 _05197_ _05198_ _05201_ net626 vssd1 vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__a311o_1
XANTENNA__09102__B1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08519_ net880 _04155_ _04157_ vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_65_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout714_X net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09499_ top.CPU.registers.data\[929\] top.CPU.registers.data\[897\] top.CPU.registers.data\[801\]
+ top.CPU.registers.data\[769\] net1000 net921 vssd1 vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__mux4_1
X_11530_ net3793 net250 _06734_ _06497_ vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__a22o_1
XFILLER_12_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_137_Right_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11042__B _05694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11461_ _06253_ net3518 net264 vssd1 vssd1 vccd1 vccd1 _02061_ sky130_fd_sc_hd__mux2_1
XANTENNA__08208__A2 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14830__1000 clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 net2469 sky130_fd_sc_hd__inv_2
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13200_ _02773_ _02778_ _02779_ net3571 vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__a22o_1
XANTENNA__07947__S net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10412_ _05997_ _06039_ net310 vssd1 vssd1 vccd1 vccd1 _06040_ sky130_fd_sc_hd__mux2_1
XANTENNA__11212__B2 _03190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11392_ _06514_ net281 net273 net3843 vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__a22o_1
XANTENNA__08613__C1 top.CPU.control_unit.instruction\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_152_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10881__B _06471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11469__S net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07967__A1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13131_ _06887_ _07428_ vssd1 vssd1 vccd1 vccd1 _02734_ sky130_fd_sc_hd__nor2_1
XFILLER_174_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10343_ _03859_ _05973_ vssd1 vssd1 vccd1 vccd1 _05974_ sky130_fd_sc_hd__xnor2_1
XFILLER_152_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08351__B net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09708__A2 net1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13062_ net2790 top.CPU.data_out\[9\] net557 vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__mux2_1
X_10274_ net530 _05907_ vssd1 vssd1 vccd1 vccd1 _05908_ sky130_fd_sc_hd__nor2_1
XANTENNA__11515__A2 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12013_ net363 _06719_ _06783_ _06782_ vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__a31o_1
Xfanout1401 net1402 vssd1 vssd1 vccd1 vccd1 net1401 sky130_fd_sc_hd__buf_4
XANTENNA__10723__B1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout480 net481 vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_161_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout491 net497 vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_161_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12476__B1 _04155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08144__A1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15703_ net2037 _01913_ net1180 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[503\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09341__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12915_ top.CPU.alu.program_counter\[27\] _05429_ vssd1 vssd1 vccd1 vccd1 _07358_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08695__A2 net1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15634_ net1968 _01844_ net1100 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[434\]
+ sky130_fd_sc_hd__dfrtp_1
X_12846_ top.CPU.alu.program_counter\[19\] _03986_ _07280_ _07294_ _07292_ vssd1 vssd1
+ vccd1 vccd1 _07296_ sky130_fd_sc_hd__o221a_1
XFILLER_73_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15565_ net1899 _01775_ net1059 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[365\]
+ sky130_fd_sc_hd__dfrtp_1
X_12777_ top.CPU.alu.program_counter\[14\] _04325_ vssd1 vssd1 vccd1 vccd1 _07233_
+ sky130_fd_sc_hd__or2_1
XANTENNA__08447__A2 net1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11728_ net1401 net534 net233 vssd1 vssd1 vccd1 vccd1 _06759_ sky130_fd_sc_hd__nand3_1
X_15496_ net1830 _01706_ net1088 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[296\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_80_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_104_Right_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11659_ _06430_ net205 net426 net3134 vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__a22o_1
XFILLER_128_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11203__B2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08542__A net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold906 top.CPU.registers.data\[791\] vssd1 vssd1 vccd1 vccd1 net3463 sky130_fd_sc_hd__dlygate4sd3_1
Xhold917 _03055_ vssd1 vssd1 vccd1 vccd1 net3474 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16117_ net2451 _02327_ net1216 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[917\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11754__A2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13329_ top.I2C.data_out\[6\] net553 _02865_ net596 vssd1 vssd1 vccd1 vccd1 _02866_
+ sky130_fd_sc_hd__a22o_1
XFILLER_116_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold928 top.CPU.registers.data\[118\] vssd1 vssd1 vccd1 vccd1 net3485 sky130_fd_sc_hd__dlygate4sd3_1
Xhold939 net84 vssd1 vssd1 vccd1 vccd1 net3496 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_50_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16048_ net2382 _02258_ net1106 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[848\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12164__C1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11506__A2 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08907__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14151__321 clknet_leaf_183_clk vssd1 vssd1 vccd1 vccd1 net1790 sky130_fd_sc_hd__inv_2
X_08870_ net784 _04508_ vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__or2_1
XFILLER_97_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10714__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14448__618 clknet_leaf_197_clk vssd1 vssd1 vccd1 vccd1 net2087 sky130_fd_sc_hd__inv_2
X_07821_ top.CPU.registers.data\[349\] net1318 net849 top.CPU.registers.data\[381\]
+ net768 vssd1 vssd1 vccd1 vccd1 _03460_ sky130_fd_sc_hd__a221o_1
XANTENNA__13607__B _05988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09007__S0 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12511__B _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07591__C1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07605__B net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07752_ top.CPU.registers.data\[190\] top.CPU.registers.data\[158\] net834 vssd1
+ vssd1 vccd1 vccd1 _03391_ sky130_fd_sc_hd__mux2_1
XANTENNA__12467__B1 _03887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07683_ _03270_ _03284_ vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__nor2_4
XFILLER_64_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09422_ net677 _05059_ _05060_ vssd1 vssd1 vccd1 vccd1 _05061_ sky130_fd_sc_hd__and3_1
XANTENNA__10493__A2 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11690__A1 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07894__B1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08276__X _03915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07621__A net1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09353_ top.CPU.registers.data\[291\] top.CPU.registers.data\[259\] net990 vssd1
+ vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__mux2_1
XANTENNA__08438__A2 net1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09096__C1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout242_A net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08304_ net695 _03941_ _03942_ vssd1 vssd1 vccd1 vccd1 _03943_ sky130_fd_sc_hd__and3_1
XANTENNA__11143__A net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11442__A1 _05960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09284_ _04891_ _04920_ vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_43_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11993__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08235_ top.CPU.registers.data\[758\] net1392 net835 top.CPU.registers.data\[726\]
+ net731 vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__a221o_1
XFILLER_20_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10982__A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1151_A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout128_X net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1249_A net1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08166_ top.CPU.registers.data\[599\] net1325 net856 top.CPU.registers.data\[631\]
+ net748 vssd1 vssd1 vccd1 vccd1 _03805_ sky130_fd_sc_hd__a221o_1
XFILLER_134_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08452__A _04090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11745__A2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10402__C1 _06028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08097_ top.CPU.registers.data\[85\] net1330 net861 top.CPU.registers.data\[117\]
+ net776 vssd1 vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__a221o_1
XANTENNA__08071__B1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08610__A2 net1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1037_X net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload90 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 clkload90/Y sky130_fd_sc_hd__inv_12
XFILLER_134_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13498__A2 _02967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout497_X net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout876_A net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09571__B1 net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12170__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout664_X net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08999_ _04636_ _04637_ net672 vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__o21a_1
XFILLER_130_895 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07582__C1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09323__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12140__C net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11037__B net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10961_ net3720 net218 _06531_ net317 vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout831_X net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08677__A2 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout929_X net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13533__A _05361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12700_ top.CPU.alu.program_counter\[6\] _03118_ _07161_ _07163_ vssd1 vssd1 vccd1
+ vccd1 _01169_ sky130_fd_sc_hd__a22o_1
X_13680_ net2640 net337 vssd1 vssd1 vccd1 vccd1 _02608_ sky130_fd_sc_hd__and2_1
X_10892_ net3555 net223 _06489_ net467 vssd1 vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__a22o_1
XANTENNA__10876__B _05906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07531__A top.CPU.control_unit.instruction\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12631_ net2608 net35 vssd1 vssd1 vccd1 vccd1 top.I2C.inter_received_n sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_100_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10368__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09626__A1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08429__A2 net1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13422__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11053__A _06056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11433__A1 _06577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15350_ net1684 _01560_ net1229 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[150\]
+ sky130_fd_sc_hd__dfrtp_1
X_12562_ _06087_ _06102_ _06124_ _07066_ vssd1 vssd1 vccd1 vccd1 _07067_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_80_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08834__C1 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11984__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11513_ net492 net137 net356 net253 net2855 vssd1 vssd1 vccd1 vccd1 _02016_ sky130_fd_sc_hd__a32o_1
X_15281_ net1615 _01491_ net1191 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[81\]
+ sky130_fd_sc_hd__dfrtp_1
X_12493_ _04890_ _04918_ _04952_ _04986_ vssd1 vssd1 vccd1 vccd1 _07002_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_11_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14592__762 clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 net2231 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_22_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11444_ net567 net530 _05694_ _06487_ vssd1 vssd1 vccd1 vccd1 _06722_ sky130_fd_sc_hd__and4_1
XFILLER_153_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11736__A2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11375_ net474 _06490_ net273 net3277 vssd1 vssd1 vccd1 vccd1 _02135_ sky130_fd_sc_hd__a22o_1
XFILLER_153_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13114_ top.SPI.command\[3\] net1410 top.SPI.paroutput\[27\] net1358 vssd1 vssd1
+ vccd1 vccd1 _02722_ sky130_fd_sc_hd__a22o_1
XFILLER_4_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10326_ _05595_ _05951_ _05957_ vssd1 vssd1 vccd1 vccd1 _05958_ sky130_fd_sc_hd__a21oi_4
X_14135__305 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 net1774 sky130_fd_sc_hd__inv_2
XFILLER_152_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13045_ top.SPI.parameters\[24\] top.SPI.paroutput\[16\] net1357 vssd1 vssd1 vccd1
+ vccd1 _07448_ sky130_fd_sc_hd__mux2_1
XFILLER_124_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10257_ _05890_ vssd1 vssd1 vccd1 vccd1 _05891_ sky130_fd_sc_hd__inv_2
XANTENNA__09011__C1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1220 net1226 vssd1 vssd1 vccd1 vccd1 net1220 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08365__A1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12161__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1231 net1232 vssd1 vssd1 vccd1 vccd1 net1231 sky130_fd_sc_hd__clkbuf_4
Xfanout1242 net1276 vssd1 vssd1 vccd1 vccd1 net1242 sky130_fd_sc_hd__clkbuf_4
X_10188_ _05817_ _05823_ net400 vssd1 vssd1 vccd1 vccd1 _05824_ sky130_fd_sc_hd__mux2_2
Xfanout1253 net1254 vssd1 vssd1 vccd1 vccd1 net1253 sky130_fd_sc_hd__clkbuf_4
XFILLER_67_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1264 net1266 vssd1 vssd1 vccd1 vccd1 net1264 sky130_fd_sc_hd__clkbuf_4
XFILLER_38_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1275 net1276 vssd1 vssd1 vccd1 vccd1 net1275 sky130_fd_sc_hd__buf_2
XFILLER_15_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1286 net1293 vssd1 vssd1 vccd1 vccd1 net1286 sky130_fd_sc_hd__clkbuf_4
XFILLER_93_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13146__C top.CPU.alu.program_counter\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14996_ clknet_leaf_92_clk _01241_ net1269 vssd1 vssd1 vccd1 vccd1 top.SPI.counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1297 net1301 vssd1 vssd1 vccd1 vccd1 net1297 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08117__A1 net1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09921__A _04829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11672__A1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15617_ net1951 _01827_ net1232 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[417\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10278__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12829_ _07278_ _07279_ vssd1 vssd1 vccd1 vccd1 _07281_ sky130_fd_sc_hd__nor2_1
XFILLER_43_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15548_ net1882 _01758_ net1195 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[348\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_139_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07723__S0 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11975__A2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_150_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_150_clk
+ sky130_fd_sc_hd__clkbuf_8
X_15479_ net1813 _01689_ net1181 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[279\]
+ sky130_fd_sc_hd__dfrtp_1
X_08020_ top.CPU.registers.data\[468\] net1318 net849 top.CPU.registers.data\[500\]
+ net768 vssd1 vssd1 vccd1 vccd1 _03659_ sky130_fd_sc_hd__a221o_1
XANTENNA__09368__A net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold703 top.mmio.mem_data_i\[16\] vssd1 vssd1 vccd1 vccd1 net3260 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11727__A2 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold714 top.CPU.registers.data\[375\] vssd1 vssd1 vccd1 vccd1 net3271 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08053__B1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold725 top.CPU.registers.data\[146\] vssd1 vssd1 vccd1 vccd1 net3282 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold736 top.CPU.registers.data\[357\] vssd1 vssd1 vccd1 vccd1 net3293 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10935__B1 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold747 top.CPU.registers.data\[266\] vssd1 vssd1 vccd1 vccd1 net3304 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16017__RESET_B net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14901__1071 clknet_leaf_172_clk vssd1 vssd1 vccd1 vccd1 net2540 sky130_fd_sc_hd__inv_2
XFILLER_157_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold758 top.CPU.registers.data\[322\] vssd1 vssd1 vccd1 vccd1 net3315 sky130_fd_sc_hd__dlygate4sd3_1
X_09971_ _03375_ _05609_ vssd1 vssd1 vccd1 vccd1 _05610_ sky130_fd_sc_hd__nor2_1
Xhold769 top.CPU.registers.data\[947\] vssd1 vssd1 vccd1 vccd1 net3326 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08922_ net787 _04559_ _04560_ net715 vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__o211a_1
XANTENNA__08356__A1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12152__A2 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07616__A net1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13337__B net1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08853_ top.CPU.registers.data\[331\] net1370 net967 top.CPU.registers.data\[363\]
+ net1280 vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__o221a_1
Xhold1403 top.CPU.registers.data\[102\] vssd1 vssd1 vccd1 vccd1 net3960 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11360__B1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout192_A net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1414 top.CPU.registers.data\[90\] vssd1 vssd1 vccd1 vccd1 net3971 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1425 top.I2C.I2C_state\[3\] vssd1 vssd1 vccd1 vccd1 net3982 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07804_ _03407_ _03440_ vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__or2_1
XANTENNA__11138__A net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1436 top.CPU.registers.data\[110\] vssd1 vssd1 vccd1 vccd1 net3993 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1447 top.SPI.timem\[20\] vssd1 vssd1 vccd1 vccd1 net4004 sky130_fd_sc_hd__dlygate4sd3_1
X_08784_ net789 _04418_ _04419_ net718 vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__o211a_1
Xhold1458 top.mmio.mem_data_i\[17\] vssd1 vssd1 vccd1 vccd1 net4015 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1469 top.CPU.addressnew\[10\] vssd1 vssd1 vccd1 vccd1 net4026 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09305__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07735_ _03372_ _03373_ vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__or2_2
XFILLER_77_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08659__A2 net1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09856__A1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout457_A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11663__A1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07666_ _03262_ _03299_ _03300_ _03303_ vssd1 vssd1 vccd1 vccd1 _03305_ sky130_fd_sc_hd__a31o_1
XANTENNA__12860__B1 _03756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10696__B _06311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09405_ top.CPU.registers.data\[963\] net1328 net859 top.CPU.registers.data\[995\]
+ net727 vssd1 vssd1 vccd1 vccd1 _05044_ sky130_fd_sc_hd__a221o_1
XFILLER_164_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10188__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09608__A1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09069__C1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout245_X net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout624_A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07597_ top.CPU.registers.data\[127\] net1334 net865 top.CPU.registers.data\[95\]
+ net731 vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__o221a_1
XANTENNA__12207__A3 _06678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1366_A net1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09336_ top.CPU.registers.data\[580\] net1329 net860 top.CPU.registers.data\[612\]
+ net752 vssd1 vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__a221o_1
XANTENNA__08881__S net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14576__746 clknet_leaf_196_clk vssd1 vssd1 vccd1 vccd1 net2215 sky130_fd_sc_hd__inv_2
XANTENNA__08816__C1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11966__A2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout412_X net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09267_ top.CPU.registers.data\[741\] net1374 net971 top.CPU.registers.data\[709\]
+ net902 vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_141_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_141_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_166_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08218_ _03822_ _03855_ vssd1 vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__nand2_1
X_14320__490 clknet_leaf_197_clk vssd1 vssd1 vccd1 vccd1 net1959 sky130_fd_sc_hd__inv_2
XFILLER_5_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08182__A top.CPU.alu.program_counter\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09198_ _04835_ _04836_ net930 vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout993_A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14617__787 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 net2256 sky130_fd_sc_hd__inv_2
XANTENNA__11718__A2 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08149_ _03787_ vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__inv_2
XFILLER_107_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1321_X net1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload190 clknet_leaf_91_clk vssd1 vssd1 vccd1 vccd1 clkload190/X sky130_fd_sc_hd__clkbuf_4
X_11160_ net3729 net304 _06640_ net319 vssd1 vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout781_X net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout879_X net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10111_ _03407_ net379 _05748_ net309 vssd1 vssd1 vccd1 vccd1 _05749_ sky130_fd_sc_hd__o211a_1
XFILLER_121_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11091_ net652 net502 vssd1 vssd1 vccd1 vccd1 _06602_ sky130_fd_sc_hd__and2_2
XFILLER_0_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08347__A1 top.CPU.control_unit.instruction\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_49_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10042_ top.CPU.alu.immediate\[31\] net507 _05680_ _03372_ _05675_ vssd1 vssd1 vccd1
+ vccd1 _05681_ sky130_fd_sc_hd__a221o_1
XANTENNA__12143__A2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11351__B1 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold30 top.CPU.registers.data_out_r1_prev\[6\] vssd1 vssd1 vccd1 vccd1 net2587 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold41 top.CPU.registers.data_out_r2_prev\[2\] vssd1 vssd1 vccd1 vccd1 net2598 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 top.CPU.registers.data_out_r1_prev\[26\] vssd1 vssd1 vccd1 vccd1 net2609 sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 top.I2C.I2C_state\[20\] vssd1 vssd1 vccd1 vccd1 net2620 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold74 top.CPU.registers.data_out_r2_prev\[0\] vssd1 vssd1 vccd1 vccd1 net2631 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 top.CPU.registers.data\[831\] vssd1 vssd1 vccd1 vccd1 net2642 sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 top.SPI.percount\[0\] vssd1 vssd1 vccd1 vccd1 net2653 sky130_fd_sc_hd__dlygate4sd3_1
X_13801_ net2802 net335 net328 top.CPU.data_out\[3\] vssd1 vssd1 vccd1 vccd1 _02681_
+ sky130_fd_sc_hd__a22o_1
XFILLER_63_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input18_A DAT_I[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11993_ _06558_ net341 net180 net2787 vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__a22o_1
XANTENNA__11103__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16520_ clknet_leaf_100_clk _02682_ net1255 vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__dfrtp_1
X_13732_ net4014 _03073_ _03075_ _07113_ vssd1 vssd1 vccd1 vccd1 _02633_ sky130_fd_sc_hd__o211a_1
XFILLER_56_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12851__A0 _07300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10944_ net521 _05693_ _06519_ vssd1 vssd1 vccd1 vccd1 _06521_ sky130_fd_sc_hd__and3_1
XFILLER_43_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08357__A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16451_ clknet_leaf_81_clk _02614_ net1263 vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_27_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13663_ top.wm.curr_state\[2\] top.wm.curr_state\[1\] top.wm.curr_state\[0\] _07091_
+ vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__and4bb_2
XTAP_TAPCELL_ROW_27_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10875_ net3659 net222 _06477_ net466 vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__a22o_1
X_15402_ net1736 _01612_ net1085 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[202\]
+ sky130_fd_sc_hd__dfrtp_1
X_12614_ _07097_ _07103_ _07113_ vssd1 vssd1 vccd1 vccd1 _07114_ sky130_fd_sc_hd__a21bo_1
X_16382_ clknet_leaf_63_clk _02591_ net1144 vssd1 vssd1 vccd1 vccd1 top.CPU.fetch.current_ra\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_156_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13594_ top.CPU.alu.program_counter\[18\] net1349 net583 vssd1 vssd1 vccd1 vccd1
+ _03023_ sky130_fd_sc_hd__o21a_1
XANTENNA__09075__A2 net1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08807__C1 net1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15333_ net1667 _01543_ net1063 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[133\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11957__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12545_ _03133_ top.mmio.m2 top.mmio.m1 top.mmio.s2 _03134_ vssd1 vssd1 vccd1 vccd1
+ _07054_ sky130_fd_sc_hd__a32oi_4
XANTENNA__09480__C1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_132_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_132_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08822__A2 _04459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13202__S _02780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15264_ net1598 _01474_ net1096 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[64\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_145_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08092__A net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12476_ _04090_ _04122_ _04155_ _04188_ vssd1 vssd1 vccd1 vccd1 _06985_ sky130_fd_sc_hd__a22o_1
XANTENNA__11709__A2 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11427_ _06569_ net280 net267 net3096 vssd1 vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__a22o_1
XANTENNA__08035__B1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_5 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15195_ net1532 _01405_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r1_prev\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08586__A1 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11358_ net3567 net287 net284 _06393_ vssd1 vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__a22o_1
XFILLER_140_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07794__C1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10309_ _03613_ _05332_ net380 vssd1 vssd1 vccd1 vccd1 _05941_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11289_ net3510 net291 _06703_ net496 vssd1 vssd1 vccd1 vccd1 _02209_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_5_Left_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08338__A1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12134__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09535__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13028_ net2746 _07439_ net894 vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__mux2_1
XFILLER_140_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_199_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_199_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_67_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11342__B1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1050 _03093_ vssd1 vssd1 vccd1 vccd1 net1050 sky130_fd_sc_hd__buf_2
Xfanout1061 net1068 vssd1 vssd1 vccd1 vccd1 net1061 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1072 net1074 vssd1 vssd1 vccd1 vccd1 net1072 sky130_fd_sc_hd__clkbuf_4
Xfanout1083 net1086 vssd1 vssd1 vccd1 vccd1 net1083 sky130_fd_sc_hd__clkbuf_4
XFILLER_13_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07870__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1094 net1097 vssd1 vssd1 vccd1 vccd1 net1094 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13095__A0 top.CPU.data_out\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09299__C1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14979_ clknet_leaf_95_clk _01224_ net1260 vssd1 vssd1 vccd1 vccd1 top.SPI.paroutput\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_07520_ top.CPU.control_unit.instruction\[0\] top.CPU.control_unit.instruction\[1\]
+ top.CPU.control_unit.instruction\[3\] _03157_ vssd1 vssd1 vccd1 vccd1 _03159_ sky130_fd_sc_hd__nand4_4
XFILLER_81_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10448__A2 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14263__433 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 net1902 sky130_fd_sc_hd__inv_2
XANTENNA__16257__Q top.CPU.handler.toreg\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14304__474 clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 net1943 sky130_fd_sc_hd__inv_2
XANTENNA__11948__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09121_ net754 _04758_ _04759_ net712 vssd1 vssd1 vccd1 vccd1 _04760_ sky130_fd_sc_hd__o211a_1
XANTENNA__12070__A1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_123_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_123_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09471__C1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08813__A2 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10081__A0 _04430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09052_ top.CPU.registers.data\[232\] net1388 net808 top.CPU.registers.data\[200\]
+ net763 vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__a221o_1
X_08003_ net675 _03640_ _03641_ net604 vssd1 vssd1 vccd1 vccd1 _03642_ sky130_fd_sc_hd__a31o_1
XFILLER_163_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold500 top.CPU.registers.data\[872\] vssd1 vssd1 vccd1 vccd1 net3057 sky130_fd_sc_hd__dlygate4sd3_1
Xhold511 top.CPU.registers.data\[377\] vssd1 vssd1 vccd1 vccd1 net3068 sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 top.CPU.registers.data\[10\] vssd1 vssd1 vccd1 vccd1 net3079 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout205_A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_976 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold533 top.CPU.registers.data\[971\] vssd1 vssd1 vccd1 vccd1 net3090 sky130_fd_sc_hd__dlygate4sd3_1
Xhold544 top.CPU.fetch.current_ra\[24\] vssd1 vssd1 vccd1 vccd1 net3101 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold555 top.CPU.fetch.current_ra\[27\] vssd1 vssd1 vccd1 vccd1 net3112 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08730__A net1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold566 top.CPU.registers.data\[437\] vssd1 vssd1 vccd1 vccd1 net3123 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold577 top.CPU.registers.data\[482\] vssd1 vssd1 vccd1 vccd1 net3134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold588 top.CPU.registers.data\[191\] vssd1 vssd1 vccd1 vccd1 net3145 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09954_ _03822_ _03856_ _05590_ vssd1 vssd1 vccd1 vccd1 _05593_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_38_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold599 top.CPU.registers.data\[28\] vssd1 vssd1 vccd1 vccd1 net3156 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1114_A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09526__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12125__A2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08905_ top.CPU.registers.data\[170\] top.CPU.registers.data\[138\] net809 vssd1
+ vssd1 vccd1 vccd1 _04544_ sky130_fd_sc_hd__mux2_1
XFILLER_170_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09885_ _03476_ _03510_ _05523_ vssd1 vssd1 vccd1 vccd1 _05524_ sky130_fd_sc_hd__a21oi_2
Xhold1200 top.CPU.registers.data\[755\] vssd1 vssd1 vccd1 vccd1 net3757 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout574_A net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11333__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout195_X net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1211 top.CPU.registers.data\[79\] vssd1 vssd1 vccd1 vccd1 net3768 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1222 top.I2C.I2C_state\[4\] vssd1 vssd1 vccd1 vccd1 net3779 sky130_fd_sc_hd__dlygate4sd3_1
X_08836_ top.CPU.registers.data\[715\] net1369 net964 top.CPU.registers.data\[747\]
+ net926 vssd1 vssd1 vccd1 vccd1 _04475_ sky130_fd_sc_hd__o221a_1
Xhold1233 top.I2C.data_out\[16\] vssd1 vssd1 vccd1 vccd1 net3790 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10687__A2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1244 top.CPU.registers.data_out_r1_prev\[12\] vssd1 vssd1 vccd1 vccd1 net3801
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1255 top.CPU.registers.data\[933\] vssd1 vssd1 vccd1 vccd1 net3812 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1266 top.I2C.data_out\[23\] vssd1 vssd1 vccd1 vccd1 net3823 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1277 net95 vssd1 vssd1 vccd1 vccd1 net3834 sky130_fd_sc_hd__dlygate4sd3_1
X_08767_ top.CPU.registers.data\[908\] net1317 net848 top.CPU.registers.data\[940\]
+ net718 vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__a221o_1
Xhold1288 top.CPU.registers.data\[1015\] vssd1 vssd1 vccd1 vccd1 net3845 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout741_A net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout362_X net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1299 top.CPU.registers.data\[660\] vssd1 vssd1 vccd1 vccd1 net3856 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout839_A _03204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07718_ net681 _03355_ _03354_ net923 vssd1 vssd1 vccd1 vccd1 _03357_ sky130_fd_sc_hd__a211o_1
XANTENNA__10500__A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08698_ top.CPU.registers.data\[589\] net1311 net842 top.CPU.registers.data\[621\]
+ net738 vssd1 vssd1 vccd1 vccd1 _04337_ sky130_fd_sc_hd__a221o_1
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07649_ _03152_ _03249_ _03263_ _03287_ vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__a31o_1
XFILLER_26_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout627_X net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10660_ _05642_ _05920_ _06276_ vssd1 vssd1 vccd1 vccd1 _06277_ sky130_fd_sc_hd__a21o_1
XANTENNA__09057__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09319_ _04952_ _04956_ net455 vssd1 vssd1 vccd1 vccd1 _04958_ sky130_fd_sc_hd__mux2_1
XANTENNA__12061__A1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10591_ net603 _06210_ _06211_ vssd1 vssd1 vccd1 vccd1 _06212_ sky130_fd_sc_hd__a21o_2
Xclkbuf_leaf_114_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_114_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08183__Y _03822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13022__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08624__B net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12330_ net2563 _04594_ net1236 vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__mux2_1
XFILLER_127_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12574__A_N _06008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12146__B net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout996_X net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12261_ net3079 net145 net432 vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__mux2_1
XANTENNA__13010__B1 _07431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08568__A1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12364__A2 top.I2C.output_state\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11212_ net3622 net299 _06661_ _03190_ vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__a22o_1
XFILLER_134_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09736__A net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12192_ top.CPU.registers.data\[55\] net651 net362 vssd1 vssd1 vccd1 vccd1 _06863_
+ sky130_fd_sc_hd__o21a_1
XFILLER_150_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput42 net42 vssd1 vssd1 vccd1 vccd1 ADR_O[12] sky130_fd_sc_hd__buf_2
Xoutput53 net53 vssd1 vssd1 vccd1 vccd1 ADR_O[22] sky130_fd_sc_hd__buf_2
XANTENNA__13258__A top.I2C.output_state\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11143_ net572 net524 _06312_ vssd1 vssd1 vccd1 vccd1 _06631_ sky130_fd_sc_hd__and3_1
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 ADR_O[7] sky130_fd_sc_hd__buf_2
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 DAT_O[16] sky130_fd_sc_hd__buf_2
Xoutput86 net86 vssd1 vssd1 vccd1 vccd1 DAT_O[26] sky130_fd_sc_hd__buf_2
XANTENNA__07791__A2 net1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12116__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput97 net97 vssd1 vssd1 vccd1 vccd1 DAT_O[7] sky130_fd_sc_hd__buf_2
XFILLER_122_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15951_ net2285 _02161_ net1096 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[751\]
+ sky130_fd_sc_hd__dfrtp_1
X_11074_ net3611 net369 _06592_ net321 vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__a22o_1
XANTENNA__11324__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10025_ _03286_ _03292_ _03321_ vssd1 vssd1 vccd1 vccd1 _05664_ sky130_fd_sc_hd__o21a_4
X_15882_ net2216 _02092_ net1090 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[682\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_91_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14247__417 clknet_leaf_183_clk vssd1 vssd1 vccd1 vccd1 net1886 sky130_fd_sc_hd__inv_2
XFILLER_17_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07703__B net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10410__A net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11976_ _06533_ net352 net183 net3734 vssd1 vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__a22o_1
XANTENNA__09296__A2 net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13715_ top.SPI.timem\[9\] _03062_ vssd1 vssd1 vccd1 vccd1 _03064_ sky130_fd_sc_hd__and2_1
X_16503_ clknet_leaf_48_clk _02665_ net1128 vssd1 vssd1 vccd1 vccd1 top.mmio.mem_data_i\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_14900__1070 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 net2539 sky130_fd_sc_hd__inv_2
XFILLER_60_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10927_ _05694_ _06508_ vssd1 vssd1 vccd1 vccd1 _06510_ sky130_fd_sc_hd__nor2_2
X_16434_ clknet_leaf_67_clk _02597_ net1168 vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__dfrtp_1
X_13646_ net2740 _07274_ net663 vssd1 vssd1 vccd1 vccd1 _02580_ sky130_fd_sc_hd__mux2_1
XFILLER_72_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10858_ net3636 net226 net312 _06465_ vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__a22o_1
XANTENNA__09048__A2 net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09410__S net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_832 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16365_ clknet_leaf_58_clk _02574_ net1144 vssd1 vssd1 vccd1 vccd1 top.CPU.fetch.current_ra\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08256__B1 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13577_ top.CPU.alu.program_counter\[11\] net1350 net582 vssd1 vssd1 vccd1 vccd1
+ _03013_ sky130_fd_sc_hd__o21a_1
XANTENNA__09453__C1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_105_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_105_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10789_ net407 _05861_ _06072_ _05664_ vssd1 vssd1 vccd1 vccd1 _06400_ sky130_fd_sc_hd__a211o_1
X_15316_ net1650 _01526_ net1074 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[116\]
+ sky130_fd_sc_hd__dfrtp_1
X_12528_ _06996_ _07022_ _07035_ _07036_ vssd1 vssd1 vccd1 vccd1 _07037_ sky130_fd_sc_hd__and4_1
XFILLER_172_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16296_ clknet_leaf_108_clk _02505_ net1246 vssd1 vssd1 vccd1 vccd1 top.CPU.data_out\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_157_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_132_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08008__A0 _03645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15247_ net1581 _01457_ net1099 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_172_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12459_ _06967_ _06966_ _06965_ vssd1 vssd1 vccd1 vccd1 _06968_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_10_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09205__C1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09756__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15178_ net1515 _01388_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r1_prev\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_141_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11579__A2_N _06726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout309 net310 vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__clkbuf_2
XFILLER_99_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12107__A2 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09508__B1 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11315__B1 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09670_ top.CPU.registers.data\[185\] net1394 net837 top.CPU.registers.data\[153\]
+ net732 vssd1 vssd1 vccd1 vccd1 _05309_ sky130_fd_sc_hd__a221o_1
XFILLER_55_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08549__X _04188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08731__A1 net1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08621_ _04258_ _04259_ vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__nand2b_1
XANTENNA__13068__A0 top.CPU.data_out\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09381__A top.CPU.control_unit.instruction\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_82_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08552_ _04158_ _04190_ vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__nor2_1
XFILLER_70_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09287__A2 net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07503_ top.SPI.percount\[0\] vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_59_Left_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08483_ _04113_ _04116_ _04121_ net627 vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__a22o_2
XFILLER_50_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10841__A2 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09320__S net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08247__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_8_0_clk_X clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout322_A _03195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11151__A net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08798__A1 net1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09104_ net800 _04738_ _04739_ net754 vssd1 vssd1 vccd1 vccd1 _04743_ sky130_fd_sc_hd__o211a_1
XFILLER_164_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09035_ top.CPU.registers.data\[840\] net1314 net845 top.CPU.registers.data\[872\]
+ net740 vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout208_X net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1329_A net1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14391__561 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 net2030 sky130_fd_sc_hd__inv_2
XANTENNA__07775__S net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13543__A1 _03439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_68_Left_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold330 top.CPU.registers.data\[988\] vssd1 vssd1 vccd1 vccd1 net2887 sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 top.SPI.parameters\[16\] vssd1 vssd1 vccd1 vccd1 net2898 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10357__A1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10357__B2 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold352 top.CPU.addressnew\[22\] vssd1 vssd1 vccd1 vccd1 net2909 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11554__B1 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout691_A net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09211__A2 net1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14688__858 clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 net2327 sky130_fd_sc_hd__inv_2
XANTENNA__07758__C1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold363 top.CPU.registers.data\[571\] vssd1 vssd1 vccd1 vccd1 net2920 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout789_A net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold374 top.CPU.registers.data\[885\] vssd1 vssd1 vccd1 vccd1 net2931 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10054__X _05693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold385 top.CPU.registers.data\[984\] vssd1 vssd1 vccd1 vccd1 net2942 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold396 top.CPU.registers.data\[833\] vssd1 vssd1 vccd1 vccd1 net2953 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout810 net812 vssd1 vssd1 vccd1 vccd1 net810 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07773__A2 net1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout821 net822 vssd1 vssd1 vccd1 vccd1 net821 sky130_fd_sc_hd__clkbuf_2
X_09937_ _05293_ _05295_ _05297_ vssd1 vssd1 vccd1 vccd1 _05576_ sky130_fd_sc_hd__or3b_1
Xfanout832 net834 vssd1 vssd1 vccd1 vccd1 net832 sky130_fd_sc_hd__clkbuf_4
Xfanout843 net854 vssd1 vssd1 vccd1 vccd1 net843 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11306__B1 _06704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout956_A net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14729__899 clknet_leaf_158_clk vssd1 vssd1 vccd1 vccd1 net2368 sky130_fd_sc_hd__inv_2
XANTENNA_fanout577_X net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout854 _03203_ vssd1 vssd1 vccd1 vccd1 net854 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout865 net870 vssd1 vssd1 vccd1 vccd1 net865 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11857__A1 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout876 net877 vssd1 vssd1 vccd1 vccd1 net876 sky130_fd_sc_hd__clkbuf_8
Xfanout887 _03094_ vssd1 vssd1 vccd1 vccd1 net887 sky130_fd_sc_hd__clkbuf_2
X_09868_ _03649_ _05365_ _05366_ vssd1 vssd1 vccd1 vccd1 _05507_ sky130_fd_sc_hd__o21a_1
Xfanout898 _06894_ vssd1 vssd1 vccd1 vccd1 net898 sky130_fd_sc_hd__buf_2
Xhold1030 top.CPU.registers.data\[586\] vssd1 vssd1 vccd1 vccd1 net3587 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1041 top.CPU.registers.data\[754\] vssd1 vssd1 vccd1 vccd1 net3598 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_93_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07804__A _03407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08819_ _03116_ _04453_ _04456_ _04457_ net610 vssd1 vssd1 vccd1 vccd1 _04458_ sky130_fd_sc_hd__a311o_1
Xhold1052 top.CPU.registers.data\[182\] vssd1 vssd1 vccd1 vccd1 net3609 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1063 top.CPU.registers.data\[466\] vssd1 vssd1 vccd1 vccd1 net3620 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1074 top.CPU.registers.data\[246\] vssd1 vssd1 vccd1 vccd1 net3631 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout744_X net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09799_ top.CPU.registers.data\[570\] net838 vssd1 vssd1 vccd1 vccd1 _05438_ sky130_fd_sc_hd__or2_1
Xhold1085 top.CPU.registers.data\[1014\] vssd1 vssd1 vccd1 vccd1 net3642 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13017__S net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11326__A net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11830_ net131 net3604 net156 vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_77_Left_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1096 top.CPU.registers.data\[924\] vssd1 vssd1 vccd1 vccd1 net3653 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_165_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout911_X net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11761_ net1404 net551 _06754_ vssd1 vssd1 vccd1 vccd1 _06760_ sky130_fd_sc_hd__or3_4
XFILLER_14_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13500_ _04656_ _02967_ vssd1 vssd1 vccd1 vccd1 _02970_ sky130_fd_sc_hd__and2_1
XANTENNA__13541__A _03508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10712_ net412 _06317_ _06320_ _06326_ vssd1 vssd1 vccd1 vccd1 _06327_ sky130_fd_sc_hd__o211a_1
XFILLER_14_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11692_ _06428_ net3954 net166 vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__mux2_1
XANTENNA__08635__A net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13431_ net3894 _02864_ net120 vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__mux2_1
X_10643_ _04532_ _04567_ net376 vssd1 vssd1 vccd1 vccd1 _06261_ sky130_fd_sc_hd__mux2_1
XFILLER_139_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16150_ net2484 _02360_ net1228 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[950\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_167_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13362_ top.mmio.mem_data_i\[15\] net592 net1344 vssd1 vssd1 vccd1 vccd1 _02890_
+ sky130_fd_sc_hd__a21o_1
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10574_ _04397_ _04465_ _06152_ _06194_ net370 vssd1 vssd1 vccd1 vccd1 _06195_ sky130_fd_sc_hd__a311o_1
X_14632__802 clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 net2271 sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_5_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11793__B1 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15101_ net1483 _01314_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r2_prev\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_158_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12313_ net2576 _05428_ net1213 vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__mux2_1
X_16081_ net2415 _02291_ net1176 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[881\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_86_Left_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13293_ top.mmio.mem_data_i\[8\] _02835_ top.mmio.mem_data_i\[10\] _02834_ vssd1
+ vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__or4b_1
X_13928__98 clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 net1567 sky130_fd_sc_hd__inv_2
XFILLER_170_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15032_ clknet_leaf_89_clk _01277_ net1273 vssd1 vssd1 vccd1 vccd1 top.SPI.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_12244_ net3244 _06478_ net434 vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__mux2_1
XANTENNA__10348__A1 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11545__B1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12175_ net3935 net175 _06855_ _06520_ vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__a22o_1
XANTENNA__10405__A net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11126_ net1405 net576 net525 net143 vssd1 vssd1 vccd1 vccd1 _06621_ sky130_fd_sc_hd__and4_1
XFILLER_111_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09913__B _05123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11057_ net324 net141 net536 net367 net2643 vssd1 vssd1 vccd1 vccd1 _02324_ sky130_fd_sc_hd__a32o_1
X_15934_ net2268 _02144_ net1204 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[734\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08174__C1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09061__S1 net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10008_ _03822_ _03889_ net379 vssd1 vssd1 vccd1 vccd1 _05647_ sky130_fd_sc_hd__mux2_1
XFILLER_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_95_Left_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10520__A1 _03315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15865_ net2199 _02075_ net1245 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[665\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_64_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10520__B2 _04189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07921__C1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11236__A net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15796_ net2130 _02006_ net1074 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[596\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_92_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10808__C1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13470__A0 top.CPU.handler.toreg\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11076__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11959_ _06506_ net341 net229 net3727 vssd1 vssd1 vccd1 vccd1 _01611_ sky130_fd_sc_hd__a22o_1
XANTENNA__08477__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10284__B1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09140__S net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16417_ clknet_leaf_56_clk net2566 net1141 vssd1 vssd1 vccd1 vccd1 top.I2C.I2C_state\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13629_ net3137 top.CPU.alu.program_counter\[1\] net663 vssd1 vssd1 vccd1 vccd1 _02563_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09426__C1 net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16348_ clknet_leaf_80_clk _02557_ net1241 vssd1 vssd1 vccd1 vccd1 top.CPU.addressnew\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10587__A1 _05643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11784__B1 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14375__545 clknet_leaf_185_clk vssd1 vssd1 vccd1 vccd1 net2014 sky130_fd_sc_hd__inv_2
X_16279_ clknet_leaf_43_clk _02489_ net1123 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.toreg\[23\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_8_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08280__A _03889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11536__B1 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10960__D net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14416__586 clknet_leaf_196_clk vssd1 vssd1 vccd1 vccd1 net2055 sky130_fd_sc_hd__inv_2
XANTENNA__11000__A2 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08401__B1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout128 net129 vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__buf_4
XFILLER_113_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout139 _06126_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__buf_2
X_07983_ top.CPU.registers.data\[600\] net1289 net1009 top.CPU.registers.data\[632\]
+ net932 vssd1 vssd1 vccd1 vccd1 _03622_ sky130_fd_sc_hd__a221o_1
XANTENNA__10034__B _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09722_ _05352_ _05355_ _05360_ net629 vssd1 vssd1 vccd1 vccd1 _05361_ sky130_fd_sc_hd__a22o_4
XANTENNA__15130__SET_B net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10969__B net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08704__A1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09653_ _04192_ _05291_ vssd1 vssd1 vccd1 vccd1 _05292_ sky130_fd_sc_hd__and2_1
XFILLER_41_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout272_A _06714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08180__A2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08604_ net1284 _04241_ _04242_ vssd1 vssd1 vccd1 vccd1 _04243_ sky130_fd_sc_hd__or3_1
XFILLER_103_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09584_ top.CPU.registers.data\[416\] top.CPU.registers.data\[384\] net973 vssd1
+ vssd1 vccd1 vccd1 _05223_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_118_Right_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08535_ net610 _04172_ _04173_ vssd1 vssd1 vccd1 vccd1 _04174_ sky130_fd_sc_hd__or3_1
XANTENNA__11067__A2 _06253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08468__B1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13461__B1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1181_A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout158_X net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10275__B1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08466_ top.CPU.registers.data\[241\] top.CPU.registers.data\[209\] net988 vssd1
+ vssd1 vccd1 vccd1 _04105_ sky130_fd_sc_hd__mux2_1
X_13983__153 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 net1622 sky130_fd_sc_hd__inv_2
XANTENNA__09680__A2 net1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08397_ top.CPU.registers.data\[978\] net1287 net1006 top.CPU.registers.data\[1010\]
+ net904 vssd1 vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout704_A net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout325_X net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09432__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11775__B1 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07979__C1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12705__A top.CPU.alu.program_counter\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07994__A2 net1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09018_ _03331_ _04656_ vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__or2_1
XFILLER_163_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10290_ _05666_ _05922_ vssd1 vssd1 vccd1 vccd1 _05923_ sky130_fd_sc_hd__nand2_1
XFILLER_145_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11527__B1 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout694_X net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12424__B _06948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold160 top.CPU.registers.data\[767\] vssd1 vssd1 vccd1 vccd1 net2717 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_72_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold171 top.CPU.registers.data\[174\] vssd1 vssd1 vccd1 vccd1 net2728 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1401_X net1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold182 top.CPU.registers.data\[679\] vssd1 vssd1 vccd1 vccd1 net2739 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 top.CPU.fetch.current_ra\[17\] vssd1 vssd1 vccd1 vccd1 net2750 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08943__A1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout861_X net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout640 net641 vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__buf_4
XANTENNA_fanout959_X net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout651 net652 vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__clkbuf_4
Xfanout662 _03168_ vssd1 vssd1 vccd1 vccd1 net662 sky130_fd_sc_hd__buf_6
XFILLER_120_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout673 net676 vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__buf_4
XANTENNA__08156__C1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout684 _03336_ vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10879__B _05693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout695 net697 vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12931_ _07371_ _07372_ vssd1 vssd1 vccd1 vccd1 _07373_ sky130_fd_sc_hd__nor2_1
XANTENNA__07534__A net1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12862_ top.CPU.alu.program_counter\[21\] _03756_ _07296_ _07308_ _07307_ vssd1 vssd1
+ vccd1 vccd1 _07310_ sky130_fd_sc_hd__o221a_1
X_15650_ net1984 _01860_ net1171 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[450\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11813_ top.CPU.registers.data\[336\] net159 vssd1 vssd1 vccd1 vccd1 _06765_ sky130_fd_sc_hd__and2_1
XANTENNA__08459__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12255__A1 _06149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15581_ net1915 _01791_ net1113 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[381\]
+ sky130_fd_sc_hd__dfrtp_1
X_12793_ _07246_ _07247_ vssd1 vssd1 vccd1 vccd1 _07248_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_1_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10895__A net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11744_ net146 net537 net499 net193 net2797 vssd1 vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_120_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14062__232 clknet_leaf_121_clk vssd1 vssd1 vccd1 vccd1 net1701 sky130_fd_sc_hd__inv_2
XANTENNA__09408__C1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11675_ net465 _06492_ net238 net166 net3060 vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__a32o_1
XANTENNA__10018__A0 _05399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14359__529 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 net1998 sky130_fd_sc_hd__inv_2
X_13414_ top.I2C.data_out\[29\] net555 _02859_ top.mmio.mem_data_i\[29\] vssd1 vssd1
+ vccd1 vccd1 _02928_ sky130_fd_sc_hd__a22o_1
XFILLER_128_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16202_ net2536 _02412_ net1084 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[1002\]
+ sky130_fd_sc_hd__dfrtp_1
X_10626_ net406 _06244_ vssd1 vssd1 vccd1 vccd1 _06245_ sky130_fd_sc_hd__nor2_1
XANTENNA__10119__B net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11766__B1 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16133_ net2467 _02343_ net1062 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[933\]
+ sky130_fd_sc_hd__dfrtp_1
X_13345_ _02830_ _02877_ vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__nor2_1
X_14103__273 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 net1742 sky130_fd_sc_hd__inv_2
X_10557_ _06089_ _06178_ net387 vssd1 vssd1 vccd1 vccd1 _06179_ sky130_fd_sc_hd__mux2_1
XANTENNA__09908__B _05266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08812__B net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13507__B2 _02973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16064_ net2398 _02274_ net1092 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[864\]
+ sky130_fd_sc_hd__dfrtp_1
X_13276_ top.CPU.handler.state\[5\] net1353 top.CPU.control_unit.instruction\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02823_ sky130_fd_sc_hd__o21a_1
X_10488_ net395 _06112_ _06110_ vssd1 vssd1 vccd1 vccd1 _06113_ sky130_fd_sc_hd__o21ai_1
XFILLER_142_326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11518__B1 _06734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15015_ clknet_leaf_95_clk _01260_ net1260 vssd1 vssd1 vccd1 vccd1 top.SPI.parameters\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_170_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12227_ _06374_ net542 _06796_ net168 top.CPU.registers.data\[37\] vssd1 vssd1 vccd1
+ vccd1 _06880_ sky130_fd_sc_hd__a32o_1
XFILLER_170_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_166_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09924__A _04765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11533__A3 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12158_ top.CPU.registers.data\[73\] net645 net144 net360 net354 vssd1 vssd1 vccd1
+ vccd1 _06847_ sky130_fd_sc_hd__o2111a_1
X_11109_ net3869 net302 _06612_ net313 vssd1 vssd1 vccd1 vccd1 _02298_ sky130_fd_sc_hd__a22o_1
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12089_ net562 net360 _06625_ net176 top.CPU.registers.data\[108\] vssd1 vssd1 vccd1
+ vccd1 _06813_ sky130_fd_sc_hd__a32o_1
XANTENNA__09135__S net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14760__930 clknet_leaf_126_clk vssd1 vssd1 vccd1 vccd1 net2399 sky130_fd_sc_hd__inv_2
XFILLER_110_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15917_ net2251 _02127_ net1069 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[717\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12494__A1 _04952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08698__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11297__A2 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12494__B2 _05054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15848_ net2182 _02058_ net1100 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[648\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_94_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14801__971 clknet_leaf_188_clk vssd1 vssd1 vccd1 vccd1 net2440 sky130_fd_sc_hd__inv_2
XFILLER_92_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13967__137 clknet_leaf_192_clk vssd1 vssd1 vccd1 vccd1 net1606 sky130_fd_sc_hd__inv_2
X_15779_ net2113 _01989_ net1207 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[579\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08320_ net880 _03955_ _03957_ vssd1 vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__o21a_1
XFILLER_21_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08251_ top.CPU.registers.data\[310\] top.CPU.registers.data\[278\] net998 vssd1
+ vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__mux2_1
XANTENNA__10955__D net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10009__A0 _03683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12549__A2 _03152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08182_ top.CPU.alu.program_counter\[23\] net1035 vssd1 vssd1 vccd1 vccd1 _03821_
+ sky130_fd_sc_hd__nor2_1
Xteam_08_1440 vssd1 vssd1 vccd1 vccd1 team_08_1440/HI gpio_out[25] sky130_fd_sc_hd__conb_1
XANTENNA__11757__A0 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_08_1451 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] team_08_1451/LO sky130_fd_sc_hd__conb_1
XANTENNA__10029__B _05667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_08_1462 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] team_08_1462/LO sky130_fd_sc_hd__conb_1
XFILLER_146_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11221__A2 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10971__C _06523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07976__A2 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10980__B2 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08925__A1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12182__B1 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10732__A1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout487_A net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07966_ net719 _03602_ _03603_ _03604_ vssd1 vssd1 vccd1 vccd1 _03605_ sky130_fd_sc_hd__a31o_1
XFILLER_101_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08138__C1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09705_ top.CPU.registers.data\[217\] net1001 net960 _05343_ vssd1 vssd1 vccd1 vccd1
+ _05344_ sky130_fd_sc_hd__a211o_1
XFILLER_74_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07897_ net712 _03534_ _03535_ vssd1 vssd1 vccd1 vccd1 _03536_ sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_94_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_94_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout654_A net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout275_X net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1396_A net1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09636_ _04862_ _04923_ _05274_ vssd1 vssd1 vccd1 vccd1 _05275_ sky130_fd_sc_hd__or3_1
XFILLER_55_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08884__S net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09567_ net929 _05204_ _05205_ net951 vssd1 vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__o211a_1
XANTENNA__13434__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout442_X net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout821_A net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14046__216 clknet_leaf_150_clk vssd1 vssd1 vccd1 vccd1 net1685 sky130_fd_sc_hd__inv_2
XFILLER_24_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout919_A net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08518_ top.CPU.alu.program_counter\[16\] net878 vssd1 vssd1 vccd1 vccd1 _04157_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_65_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09498_ net945 _05134_ _05136_ net622 vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__o211a_1
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10799__A1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08310__C1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11996__B1 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08449_ _04084_ _04087_ net1308 vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__o21a_1
XFILLER_157_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout707_X net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11460_ _06230_ net3652 net263 vssd1 vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__mux2_1
XANTENNA__09405__A2 net1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11748__B1 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10411_ _03683_ _03755_ net378 vssd1 vssd1 vccd1 vccd1 _06039_ sky130_fd_sc_hd__mux2_1
XANTENNA__16552__D net4000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11212__A2 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11391_ net480 net472 _06513_ net271 net3160 vssd1 vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13130_ _07095_ _02728_ _02730_ _02732_ vssd1 vssd1 vccd1 vccd1 _02733_ sky130_fd_sc_hd__nor4_1
XFILLER_137_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10342_ _03923_ _05972_ _05591_ vssd1 vssd1 vccd1 vccd1 _05973_ sky130_fd_sc_hd__a21bo_1
XANTENNA__07529__A _03148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11763__A3 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09169__A1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13061_ net3097 top.CPU.data_out\[8\] net557 vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__mux2_1
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10273_ net575 _05906_ vssd1 vssd1 vccd1 vccd1 _05907_ sky130_fd_sc_hd__nand2_1
XANTENNA__08377__C1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12012_ top.CPU.registers.data\[155\] net653 vssd1 vssd1 vccd1 vccd1 _06783_ sky130_fd_sc_hd__or2_1
XFILLER_105_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11515__A3 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1402 top.CPU.control_unit.instruction\[10\] vssd1 vssd1 vccd1 vccd1 net1402
+ sky130_fd_sc_hd__buf_6
XFILLER_132_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14744__914 clknet_leaf_160_clk vssd1 vssd1 vccd1 vccd1 net2383 sky130_fd_sc_hd__inv_2
XFILLER_132_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11920__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_144_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_144_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout470 _03194_ vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout481 net482 vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout492 net493 vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12476__A1 _04090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12476__B2 _04188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13673__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_85_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_clk sky130_fd_sc_hd__clkbuf_8
X_15702_ net2036 _01912_ net1227 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[502\]
+ sky130_fd_sc_hd__dfrtp_1
X_12914_ top.CPU.alu.program_counter\[27\] _05429_ vssd1 vssd1 vccd1 vccd1 _07357_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_122_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12845_ top.CPU.alu.program_counter\[19\] _03986_ _07280_ _07294_ vssd1 vssd1 vccd1
+ vccd1 _07295_ sky130_fd_sc_hd__o22a_1
X_15633_ net1967 _01843_ net1189 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[433\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13205__S _02782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12776_ top.CPU.alu.program_counter\[14\] _04325_ vssd1 vssd1 vccd1 vccd1 _07232_
+ sky130_fd_sc_hd__nand2_1
X_15564_ net1898 _01774_ net1069 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[364\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_159_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11987__B1 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_14_Left_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11727_ _06573_ net198 net420 net3009 vssd1 vssd1 vccd1 vccd1 _01826_ sky130_fd_sc_hd__a22o_1
XFILLER_42_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15495_ net1829 _01705_ net1201 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[295\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11658_ _06413_ net204 net426 net3105 vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__a22o_1
XFILLER_174_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11739__B1 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10609_ top.CPU.fetch.current_ra\[12\] net1043 net882 top.CPU.handler.toreg\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06229_ sky130_fd_sc_hd__a22oi_2
XFILLER_127_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11203__A2 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11589_ net570 _06601_ vssd1 vssd1 vccd1 vccd1 _06748_ sky130_fd_sc_hd__nor2_2
XANTENNA__10411__A0 _03683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold907 top.CPU.registers.data\[229\] vssd1 vssd1 vccd1 vccd1 net3464 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07958__A2 net1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13328_ top.mmio.mem_data_i\[6\] net592 net1343 vssd1 vssd1 vccd1 vccd1 _02865_ sky130_fd_sc_hd__a21o_1
Xhold918 top.CPU.registers.data\[577\] vssd1 vssd1 vccd1 vccd1 net3475 sky130_fd_sc_hd__dlygate4sd3_1
X_16116_ net2450 _02326_ net1120 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[916\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08034__S net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold929 top.I2C.data_out\[27\] vssd1 vssd1 vccd1 vccd1 net3486 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13259_ net1053 _02813_ _02814_ net3928 vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__a22o_1
X_16047_ net2381 _02257_ net1095 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[847\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08368__C1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07873__S net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_23_Left_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14190__360 clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 net1829 sky130_fd_sc_hd__inv_2
XFILLER_151_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11911__B1 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07820_ top.CPU.registers.data\[317\] top.CPU.registers.data\[285\] net817 vssd1
+ vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__mux2_1
XFILLER_9_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13912__82 clknet_leaf_167_clk vssd1 vssd1 vccd1 vccd1 net1551 sky130_fd_sc_hd__inv_2
X_14487__657 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 net2126 sky130_fd_sc_hd__inv_2
XANTENNA__09007__S1 net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07591__B1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07751_ net778 _03378_ _03382_ _03389_ vssd1 vssd1 vccd1 vccd1 _03390_ sky130_fd_sc_hd__a31o_1
XANTENNA__15164__Q top.CPU.handler.readout vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_92_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12467__A1 _03819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12467__B2 _03915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_76_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__10478__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08135__A2 net1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09332__A1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14528__698 clknet_leaf_125_clk vssd1 vssd1 vccd1 vccd1 net2167 sky130_fd_sc_hd__inv_2
X_07682_ net632 _03320_ vssd1 vssd1 vccd1 vccd1 _03321_ sky130_fd_sc_hd__nand2_2
X_09421_ top.CPU.registers.data\[578\] net1294 net1015 top.CPU.registers.data\[610\]
+ net936 vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__a221o_1
XANTENNA__13416__A0 top.CPU.control_unit.instruction\[29\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_64_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09352_ _04988_ _04989_ vssd1 vssd1 vccd1 vccd1 _04991_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_47_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09096__B1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08303_ top.CPU.registers.data\[755\] net1393 net824 top.CPU.registers.data\[723\]
+ net724 vssd1 vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__a221o_1
XANTENNA__11978__B1 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_150_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11143__B net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09283_ _04921_ vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__inv_2
XANTENNA__11442__A2 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout235_A net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08234_ top.CPU.registers.data\[598\] net1334 net865 top.CPU.registers.data\[630\]
+ net756 vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_30_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08165_ _03800_ _03803_ net637 vssd1 vssd1 vccd1 vccd1 _03804_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_60_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout402_A net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1144_A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_165_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08096_ top.CPU.registers.data\[53\] top.CPU.registers.data\[21\] net830 vssd1 vssd1
+ vccd1 vccd1 _03735_ sky130_fd_sc_hd__mux2_1
XFILLER_173_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10046__Y _05685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14431__601 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 net2070 sky130_fd_sc_hd__inv_2
Xclkload80 clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 clkload80/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA_clkbuf_leaf_45_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload91 clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 clkload91/Y sky130_fd_sc_hd__inv_12
XFILLER_162_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1311_A net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08359__C1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout392_X net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10705__A1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout771_A net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11902__B1 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08374__A2 net1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout869_A net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08998_ top.CPU.registers.data\[713\] net1369 net965 top.CPU.registers.data\[745\]
+ net926 vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__o221a_1
XFILLER_85_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07582__B1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07949_ net1048 _03164_ net1039 net1390 top.CPU.registers.data\[440\] vssd1 vssd1
+ vccd1 vccd1 _03588_ sky130_fd_sc_hd__o311a_1
XFILLER_29_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_67_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_91_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout657_X net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1399_X net1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_170_Right_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_103_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10960_ net517 net441 net135 net546 vssd1 vssd1 vccd1 vccd1 _06531_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_67_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08531__C1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09619_ top.CPU.registers.data\[896\] net1315 net846 top.CPU.registers.data\[928\]
+ net715 vssd1 vssd1 vccd1 vccd1 _05258_ sky130_fd_sc_hd__a221o_1
XANTENNA__07885__A1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout824_X net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11681__A2 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10891_ net490 net517 _06488_ vssd1 vssd1 vccd1 vccd1 _06489_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_84_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13025__S net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12630_ _06891_ _07120_ vssd1 vssd1 vccd1 vccd1 _00044_ sky130_fd_sc_hd__and2_1
XANTENNA__07531__B net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08119__S net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11969__B1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_118_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12561_ _06147_ _06210_ _06228_ _06251_ vssd1 vssd1 vccd1 vccd1 _07066_ sky130_fd_sc_hd__and4bb_1
XFILLER_54_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11053__B net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11433__A2 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11512_ net3503 net253 _06734_ _06473_ vssd1 vssd1 vccd1 vccd1 _02017_ sky130_fd_sc_hd__a22o_1
XANTENNA__10641__B1 _05643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15280_ net1614 _01490_ net1156 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[80\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_141_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12492_ _04763_ _04792_ vssd1 vssd1 vccd1 vccd1 _07001_ sky130_fd_sc_hd__or2_1
XANTENNA__08643__A net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11443_ net133 net3635 net265 vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__mux2_1
XFILLER_137_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08598__C1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11374_ net474 _06489_ net273 net3584 vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__a22o_1
X_13113_ net2694 _02721_ net897 vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__mux2_1
X_10325_ _05300_ net447 _05936_ _05954_ _05956_ vssd1 vssd1 vccd1 vccd1 _05957_ sky130_fd_sc_hd__a311o_1
X_14174__344 clknet_leaf_154_clk vssd1 vssd1 vccd1 vccd1 net1813 sky130_fd_sc_hd__inv_2
XFILLER_112_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13044_ net2765 _07447_ net896 vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__mux2_1
XANTENNA__09474__A net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10256_ _05710_ _05717_ net388 vssd1 vssd1 vccd1 vccd1 _05890_ sky130_fd_sc_hd__mux2_1
XFILLER_61_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1210 net1212 vssd1 vssd1 vccd1 vccd1 net1210 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09562__A1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1221 net1226 vssd1 vssd1 vccd1 vccd1 net1221 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08996__S0 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1232 net1233 vssd1 vssd1 vccd1 vccd1 net1232 sky130_fd_sc_hd__buf_2
X_10187_ _05822_ vssd1 vssd1 vccd1 vccd1 _05823_ sky130_fd_sc_hd__inv_2
X_14215__385 clknet_leaf_183_clk vssd1 vssd1 vccd1 vccd1 net1854 sky130_fd_sc_hd__inv_2
Xfanout1243 net1259 vssd1 vssd1 vccd1 vccd1 net1243 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07573__B1 top.CPU.control_unit.instruction\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1254 net1258 vssd1 vssd1 vccd1 vccd1 net1254 sky130_fd_sc_hd__clkbuf_4
Xfanout1265 net1266 vssd1 vssd1 vccd1 vccd1 net1265 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08770__C1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1276 net1277 vssd1 vssd1 vccd1 vccd1 net1276 sky130_fd_sc_hd__buf_4
XFILLER_38_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11228__B net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1287 net1292 vssd1 vssd1 vccd1 vccd1 net1287 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_58_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_clk sky130_fd_sc_hd__clkbuf_8
X_14995_ clknet_leaf_92_clk _01240_ net1269 vssd1 vssd1 vccd1 vccd1 top.SPI.counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10132__B net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09314__A1 net1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1298 net1301 vssd1 vssd1 vccd1 vccd1 net1298 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13110__A2 net1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_11_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_11_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__11121__B2 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08522__C1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07876__A1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11244__A net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15616_ net1950 _01826_ net1090 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[416\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10880__B1 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12828_ _07251_ _07257_ _07266_ _07278_ _07265_ vssd1 vssd1 vccd1 vccd1 _07280_ sky130_fd_sc_hd__o311a_1
XFILLER_61_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09617__A2 net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12059__B net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12774__S net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15547_ net1881 _01757_ net1213 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[347\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11424__A2 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12759_ _07204_ _07206_ vssd1 vssd1 vccd1 vccd1 _07217_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_139_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10632__B1 _06250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07723__S1 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11898__B net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08553__A _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15478_ net1812 _01688_ net1229 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[278\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_163_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold704 top.CPU.registers.data\[677\] vssd1 vssd1 vccd1 vccd1 net3261 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08053__A1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold715 top.CPU.registers.data\[638\] vssd1 vssd1 vccd1 vccd1 net3272 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10396__C1 _05664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10935__A1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold726 top.CPU.registers.data\[353\] vssd1 vssd1 vccd1 vccd1 net3283 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_31_Left_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold737 top.CPU.registers.data\[481\] vssd1 vssd1 vccd1 vccd1 net3294 sky130_fd_sc_hd__dlygate4sd3_1
X_09970_ _05602_ _05603_ _05607_ _05608_ vssd1 vssd1 vccd1 vccd1 _05609_ sky130_fd_sc_hd__a31o_1
Xhold748 top.CPU.registers.data\[215\] vssd1 vssd1 vccd1 vccd1 net3305 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07800__A1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold759 top.CPU.registers.data\[595\] vssd1 vssd1 vccd1 vccd1 net3316 sky130_fd_sc_hd__dlygate4sd3_1
X_13889__59 clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 net1528 sky130_fd_sc_hd__inv_2
X_08921_ top.CPU.registers.data\[842\] net1313 net844 top.CPU.registers.data\[874\]
+ net765 vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__a221o_1
XANTENNA__10302__A_N _05933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09553__A1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08852_ top.CPU.registers.data\[427\] top.CPU.registers.data\[395\] top.CPU.registers.data\[299\]
+ top.CPU.registers.data\[267\] net967 net1280 vssd1 vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__mux4_1
XANTENNA__10699__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12152__A3 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07616__B _03148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1404 top.CPU.registers.data\[99\] vssd1 vssd1 vccd1 vccd1 net3961 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1415 top.CPU.registers.data\[244\] vssd1 vssd1 vccd1 vccd1 net3972 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07564__B1 net1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07803_ _03407_ _03440_ vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__nand2_1
Xhold1426 top.I2C.output_state\[10\] vssd1 vssd1 vccd1 vccd1 net3983 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1437 top.SPI.timem\[8\] vssd1 vssd1 vccd1 vccd1 net3994 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11138__B net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08783_ net704 _04420_ _04421_ vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__or3_1
Xhold1448 top.CPU.data_out\[25\] vssd1 vssd1 vccd1 vccd1 net4005 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1459 top.I2C.I2C_state\[1\] vssd1 vssd1 vccd1 vccd1 net4016 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_49_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_38_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout185_A net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07734_ net417 _03371_ vssd1 vssd1 vccd1 vccd1 _03373_ sky130_fd_sc_hd__nor2_1
XFILLER_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_40_Left_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08513__C1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07665_ _03262_ _03299_ _03300_ net631 vssd1 vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__a31oi_4
XANTENNA__07867__A1 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout352_A net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09404_ top.CPU.registers.data\[835\] net1328 net859 top.CPU.registers.data\[867\]
+ net751 vssd1 vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__a221o_1
XANTENNA__11154__A net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09069__B1 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10871__B1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07596_ top.CPU.registers.data\[159\] net1392 net836 top.CPU.registers.data\[191\]
+ net756 vssd1 vssd1 vccd1 vccd1 _03235_ sky130_fd_sc_hd__o221a_1
XFILLER_111_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09335_ top.CPU.registers.data\[836\] net1329 net860 top.CPU.registers.data\[868\]
+ net752 vssd1 vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__a221o_1
XANTENNA__11415__A2 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08816__B1 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout617_A net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout238_X net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1359_A net1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09266_ top.CPU.registers.data\[581\] net1286 net1005 top.CPU.registers.data\[613\]
+ net928 vssd1 vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__a221o_1
X_08217_ _03855_ vssd1 vssd1 vccd1 vccd1 _03856_ sky130_fd_sc_hd__inv_2
XFILLER_166_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09197_ top.CPU.registers.data\[166\] top.CPU.registers.data\[134\] net978 vssd1
+ vssd1 vccd1 vccd1 _04836_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout405_X net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1147_X net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09993__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14158__328 clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 net1797 sky130_fd_sc_hd__inv_2
X_08148_ _03755_ _03784_ vssd1 vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__nor2_1
XANTENNA__08044__A1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout986_A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08079_ _03716_ _03685_ net454 vssd1 vssd1 vccd1 vccd1 _03718_ sky130_fd_sc_hd__mux2_1
XFILLER_107_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload180 clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 clkload180/Y sky130_fd_sc_hd__inv_8
Xclkload191 clknet_leaf_92_clk vssd1 vssd1 vccd1 vccd1 clkload191/Y sky130_fd_sc_hd__bufinv_16
XANTENNA_fanout1314_X net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10110_ _03476_ net374 vssd1 vssd1 vccd1 vccd1 _05748_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_8_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11090_ _03186_ net501 vssd1 vssd1 vccd1 vccd1 _06601_ sky130_fd_sc_hd__or2_2
XFILLER_88_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout774_X net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10041_ net505 vssd1 vssd1 vccd1 vccd1 _05680_ sky130_fd_sc_hd__inv_2
XFILLER_102_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold20 top.CPU.registers.data_out_r2_prev\[28\] vssd1 vssd1 vccd1 vccd1 net2577 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 top.CPU.registers.data_out_r2_prev\[5\] vssd1 vssd1 vccd1 vccd1 net2588 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold42 top.CPU.registers.data_out_r1_prev\[24\] vssd1 vssd1 vccd1 vccd1 net2599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 top.SPI.register\[3\] vssd1 vssd1 vccd1 vccd1 net2610 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 _00034_ vssd1 vssd1 vccd1 vccd1 net2621 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout941_X net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold75 top.I2C.I2C_state\[7\] vssd1 vssd1 vccd1 vccd1 net2632 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13800_ net3014 net334 net327 top.CPU.data_out\[2\] vssd1 vssd1 vccd1 vccd1 _02680_
+ sky130_fd_sc_hd__a22o_1
XFILLER_57_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold86 top.CPU.registers.data\[914\] vssd1 vssd1 vccd1 vccd1 net2643 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07570__A3 net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold97 top.CPU.registers.data\[315\] vssd1 vssd1 vccd1 vccd1 net2654 sky130_fd_sc_hd__dlygate4sd3_1
X_11992_ _06556_ net342 net180 net2784 vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__a22o_1
XANTENNA__11103__A1 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10887__B net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08504__C1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09847__A2 net1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07542__A net1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13731_ top.SPI.timem\[13\] top.SPI.timem\[14\] _03071_ vssd1 vssd1 vccd1 vccd1 _03075_
+ sky130_fd_sc_hd__nand3_1
X_10943_ _05693_ _06519_ vssd1 vssd1 vccd1 vccd1 _06520_ sky130_fd_sc_hd__and2_1
XANTENNA__07858__A1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11654__A2 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15709__RESET_B net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11064__A _06212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16450_ clknet_leaf_81_clk _02613_ net1242 vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__dfrtp_1
X_13662_ net3951 _03044_ _03043_ vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_27_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10874_ net489 net135 net437 vssd1 vssd1 vccd1 vccd1 _06477_ sky130_fd_sc_hd__and3_1
X_15401_ net1735 _01611_ net1056 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[201\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12613_ _03127_ _03136_ _07112_ vssd1 vssd1 vccd1 vccd1 _07113_ sky130_fd_sc_hd__or3_4
X_16381_ clknet_leaf_66_clk _02590_ net1165 vssd1 vssd1 vccd1 vccd1 top.CPU.fetch.current_ra\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_13593_ net1352 _06103_ vssd1 vssd1 vccd1 vccd1 _03022_ sky130_fd_sc_hd__nand2_1
XANTENNA__11406__A2 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08807__B1 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14600__770 clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 net2239 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_156_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12544_ _07051_ _07052_ vssd1 vssd1 vccd1 vccd1 _07053_ sky130_fd_sc_hd__nand2_1
XANTENNA__09469__A net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15332_ net1666 _01542_ net1221 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[132\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10614__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10090__A1 _03755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11511__B _06726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15263_ net1597 _01473_ net1223 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[63\]
+ sky130_fd_sc_hd__dfrtp_1
X_12475_ _04090_ _04122_ vssd1 vssd1 vccd1 vccd1 _06984_ sky130_fd_sc_hd__or2_1
XFILLER_138_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11426_ _06568_ net281 net269 net2864 vssd1 vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__a22o_1
X_15194_ net1531 _01404_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r1_prev\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09232__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_6 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11230__C net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08586__A2 _04222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09783__A1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11357_ net3523 net285 net276 _06375_ vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__a22o_1
XFILLER_141_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07794__B1 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10308_ _05752_ _05939_ _05938_ vssd1 vssd1 vccd1 vccd1 _05940_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_130_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11288_ net475 net138 _06471_ net428 vssd1 vssd1 vccd1 vccd1 _06703_ sky130_fd_sc_hd__and4_1
X_13027_ top.SPI.parameters\[15\] top.SPI.paroutput\[7\] net1356 vssd1 vssd1 vccd1
+ vccd1 _07439_ sky130_fd_sc_hd__mux2_1
X_10239_ net414 _05873_ net224 vssd1 vssd1 vccd1 vccd1 _05874_ sky130_fd_sc_hd__o21ba_1
XFILLER_67_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1040 net1042 vssd1 vssd1 vccd1 vccd1 net1040 sky130_fd_sc_hd__clkbuf_4
Xfanout1051 net1052 vssd1 vssd1 vccd1 vccd1 net1051 sky130_fd_sc_hd__buf_2
Xfanout1062 net1063 vssd1 vssd1 vccd1 vccd1 net1062 sky130_fd_sc_hd__clkbuf_4
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1073 net1074 vssd1 vssd1 vccd1 vccd1 net1073 sky130_fd_sc_hd__clkbuf_2
Xfanout1084 net1086 vssd1 vssd1 vccd1 vccd1 net1084 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11673__S net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1095 net1097 vssd1 vssd1 vccd1 vccd1 net1095 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09299__B1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14978_ clknet_leaf_84_clk _01223_ net1264 vssd1 vssd1 vccd1 vccd1 top.SPI.paroutput\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09838__A2 net1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13173__B top.I2C.output_state\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11645__A2 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08510__A2 net1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14599__769 clknet_leaf_186_clk vssd1 vssd1 vccd1 vccd1 net2238 sky130_fd_sc_hd__inv_2
XFILLER_90_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09120_ top.CPU.registers.data\[903\] net1333 net864 top.CPU.registers.data\[935\]
+ net729 vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_106_Left_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10605__B1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08274__A1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12070__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09471__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16273__Q top.CPU.handler.toreg\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10081__A1 _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09051_ net785 _04686_ _04687_ net714 vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__o211a_1
XFILLER_163_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08002_ top.CPU.registers.data\[472\] net1290 net1010 top.CPU.registers.data\[504\]
+ net907 vssd1 vssd1 vccd1 vccd1 _03641_ sky130_fd_sc_hd__a221o_1
Xhold501 top.CPU.registers.data_out_r2_prev\[12\] vssd1 vssd1 vccd1 vccd1 net3058
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold512 top.CPU.registers.data\[664\] vssd1 vssd1 vccd1 vccd1 net3069 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08577__A2 net1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold523 top.CPU.registers.data\[478\] vssd1 vssd1 vccd1 vccd1 net3080 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13570__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold534 net83 vssd1 vssd1 vccd1 vccd1 net3091 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold545 top.CPU.registers.data\[412\] vssd1 vssd1 vccd1 vccd1 net3102 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold556 top.CPU.registers.data\[574\] vssd1 vssd1 vccd1 vccd1 net3113 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07785__B1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09318__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08982__C1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold567 top.CPU.registers.data_out_r2_prev\[9\] vssd1 vssd1 vccd1 vccd1 net3124 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07627__A net1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold578 top.CPU.registers.data\[732\] vssd1 vssd1 vccd1 vccd1 net3135 sky130_fd_sc_hd__dlygate4sd3_1
X_09953_ _03859_ _05591_ vssd1 vssd1 vccd1 vccd1 _05592_ sky130_fd_sc_hd__or2_1
Xhold589 top.CPU.registers.data\[635\] vssd1 vssd1 vccd1 vccd1 net3146 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_115_Left_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08329__A2 net1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09526__A1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11149__A net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08904_ net640 _04539_ _04542_ vssd1 vssd1 vccd1 vccd1 _04543_ sky130_fd_sc_hd__or3_1
XANTENNA__10373__A2_N _05733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09884_ _05512_ _05522_ vssd1 vssd1 vccd1 vccd1 _05523_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_55_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1107_A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_4_0_clk_X clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1201 top.CPU.registers.data_out_r1_prev\[30\] vssd1 vssd1 vccd1 vccd1 net3758
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1212 top.CPU.registers.data\[104\] vssd1 vssd1 vccd1 vccd1 net3769 sky130_fd_sc_hd__dlygate4sd3_1
X_08835_ top.CPU.registers.data\[587\] net1369 net964 top.CPU.registers.data\[619\]
+ net900 vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__o221a_1
Xhold1223 top.CPU.registers.data\[235\] vssd1 vssd1 vccd1 vccd1 net3780 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1234 top.CPU.registers.data\[442\] vssd1 vssd1 vccd1 vccd1 net3791 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout188_X net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout567_A net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1245 top.CPU.registers.data\[38\] vssd1 vssd1 vccd1 vccd1 net3802 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1256 top.CPU.registers.data\[1009\] vssd1 vssd1 vccd1 vccd1 net3813 sky130_fd_sc_hd__dlygate4sd3_1
X_14543__713 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 net2182 sky130_fd_sc_hd__inv_2
Xhold1267 top.I2C.data_out\[19\] vssd1 vssd1 vccd1 vccd1 net3824 sky130_fd_sc_hd__dlygate4sd3_1
X_08766_ top.CPU.registers.data\[812\] top.CPU.registers.data\[780\] net814 vssd1
+ vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__mux2_1
Xhold1278 top.CPU.registers.data\[56\] vssd1 vssd1 vccd1 vccd1 net3835 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1289 top.mmio.mem_data_i\[11\] vssd1 vssd1 vccd1 vccd1 net3846 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07717_ net959 _03350_ _03351_ net947 vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__a211o_1
XANTENNA__11097__B1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08697_ top.CPU.registers.data\[557\] top.CPU.registers.data\[525\] net808 vssd1
+ vssd1 vccd1 vccd1 _04336_ sky130_fd_sc_hd__mux2_1
XFILLER_72_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11636__A2 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15802__RESET_B net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10500__B _06124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout355_X net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout734_A net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07648_ top.CPU.control_unit.instruction\[6\] net1399 _03146_ _03149_ vssd1 vssd1
+ vccd1 vccd1 _03287_ sky130_fd_sc_hd__a211o_1
XFILLER_54_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout901_A net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout522_X net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07579_ top.CPU.registers.data\[799\] net865 net779 _03217_ vssd1 vssd1 vccd1 vccd1
+ _03218_ sky130_fd_sc_hd__o211a_1
X_09318_ _04951_ _04955_ net455 vssd1 vssd1 vccd1 vccd1 _04957_ sky130_fd_sc_hd__mux2_1
XFILLER_15_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08265__A1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10590_ top.CPU.fetch.current_ra\[13\] net1043 net882 top.CPU.handler.toreg\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06211_ sky130_fd_sc_hd__a22o_1
XANTENNA__12061__A2 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09249_ _04880_ _04881_ net786 vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__o21a_1
XANTENNA__11331__B net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_151_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12260_ net3012 net142 net431 vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__mux2_1
XFILLER_110_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09214__B1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11211_ _06428_ net430 vssd1 vssd1 vccd1 vccd1 _06661_ sky130_fd_sc_hd__and2_1
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout989_X net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13539__A _03575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12191_ net3835 net649 _06862_ vssd1 vssd1 vccd1 vccd1 _01466_ sky130_fd_sc_hd__o21a_1
XFILLER_162_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07776__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput43 net43 vssd1 vssd1 vccd1 vccd1 ADR_O[13] sky130_fd_sc_hd__buf_2
XFILLER_123_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11142_ net3595 net301 _06630_ net456 vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__a22o_1
XANTENNA__07537__A net1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13258__B net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput54 net54 vssd1 vssd1 vccd1 vccd1 ADR_O[23] sky130_fd_sc_hd__buf_2
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 ADR_O[8] sky130_fd_sc_hd__buf_2
XFILLER_150_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12162__B net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 DAT_O[17] sky130_fd_sc_hd__buf_2
XANTENNA__09517__A1 net1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput87 net87 vssd1 vssd1 vccd1 vccd1 DAT_O[27] sky130_fd_sc_hd__buf_2
XANTENNA__12116__A3 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11073_ _06333_ _06575_ vssd1 vssd1 vccd1 vccd1 _06592_ sky130_fd_sc_hd__nor2_1
X_15950_ net2284 _02160_ net1108 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[750\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput98 net98 vssd1 vssd1 vccd1 vccd1 DAT_O[8] sky130_fd_sc_hd__buf_2
XFILLER_0_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10127__A2 _05722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11324__B2 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10024_ net396 net385 _05655_ vssd1 vssd1 vccd1 vccd1 _05663_ sky130_fd_sc_hd__or3_1
XANTENNA_input30_A DAT_I[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15881_ net2215 _02091_ net1060 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[681\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11875__A2 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14286__456 clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 net1925 sky130_fd_sc_hd__inv_2
XFILLER_29_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11975_ _06531_ net348 net182 net3535 vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__a22o_1
X_16502_ clknet_leaf_48_clk _02664_ net1128 vssd1 vssd1 vccd1 vccd1 top.mmio.mem_data_i\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_13714_ _03062_ _03063_ vssd1 vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__nor2_1
XFILLER_147_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10926_ _06508_ vssd1 vssd1 vccd1 vccd1 _06509_ sky130_fd_sc_hd__inv_2
XFILLER_71_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14327__497 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 net1966 sky130_fd_sc_hd__inv_2
XFILLER_44_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16433_ clknet_leaf_66_clk _02596_ net1166 vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__dfrtp_1
XFILLER_31_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13645_ net2750 _07272_ net663 vssd1 vssd1 vccd1 vccd1 _02579_ sky130_fd_sc_hd__mux2_1
X_10857_ net1405 net576 net513 net130 vssd1 vssd1 vccd1 vccd1 _06465_ sky130_fd_sc_hd__and4_1
XFILLER_108_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16364_ clknet_leaf_45_clk _02573_ net1138 vssd1 vssd1 vccd1 vccd1 top.CPU.fetch.current_ra\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_171_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10788_ _05672_ _06079_ vssd1 vssd1 vccd1 vccd1 _06399_ sky130_fd_sc_hd__nand2_1
X_13576_ net1349 _06251_ vssd1 vssd1 vccd1 vccd1 _03012_ sky130_fd_sc_hd__nand2_1
XANTENNA__09453__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15315_ net1649 _01525_ net1176 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[115\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_145_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_719 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12527_ _07003_ _07006_ vssd1 vssd1 vccd1 vccd1 _07036_ sky130_fd_sc_hd__nor2_1
XFILLER_158_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16295_ clknet_leaf_108_clk _02504_ net1246 vssd1 vssd1 vccd1 vccd1 top.CPU.data_out\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_145_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15246_ net1580 _01456_ net1105 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09205__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12458_ _03541_ _03575_ vssd1 vssd1 vccd1 vccd1 _06967_ sky130_fd_sc_hd__nor2_1
XFILLER_172_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09756__A1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11409_ _06540_ net278 net268 net3362 vssd1 vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__a22o_1
X_12389_ top.CPU.addressnew\[1\] top.CPU.addressnew\[8\] top.CPU.addressnew\[11\]
+ _06926_ vssd1 vssd1 vccd1 vccd1 _06927_ sky130_fd_sc_hd__or4b_1
X_15177_ net1514 _01387_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r1_prev\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_141_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11563__B2 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_169_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13859__29 clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 net1498 sky130_fd_sc_hd__inv_2
X_14230__400 clknet_leaf_182_clk vssd1 vssd1 vccd1 vccd1 net1869 sky130_fd_sc_hd__inv_2
XANTENNA__10118__A2 _05742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11315__B2 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09662__A top.CPU.alu.program_counter\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08716__C1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08620_ _04225_ _04257_ vssd1 vssd1 vccd1 vccd1 _04259_ sky130_fd_sc_hd__nand2_1
XFILLER_55_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08551_ _04188_ _04189_ net455 vssd1 vssd1 vccd1 vccd1 _04190_ sky130_fd_sc_hd__mux2_1
XANTENNA__11079__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10958__D net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15284__RESET_B net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07502_ top.SPI.percount\[1\] vssd1 vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__inv_2
XANTENNA__09141__C1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08482_ net606 _04117_ _04118_ _04119_ _04120_ vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__o32a_1
XANTENNA__08495__A1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09601__S net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12579__B1 _03137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout148_A _06412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10419__A1_N _03685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09444__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12043__A2 net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09103_ net800 _04736_ _04737_ net729 vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__o211a_1
XFILLER_164_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13791__A2 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout315_A _03195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09034_ top.CPU.registers.data\[744\] net1388 net808 top.CPU.registers.data\[712\]
+ net714 vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_96_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold320 top.CPU.registers.data\[417\] vssd1 vssd1 vccd1 vccd1 net2877 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold331 top.CPU.registers.data\[851\] vssd1 vssd1 vccd1 vccd1 net2888 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold342 net92 vssd1 vssd1 vccd1 vccd1 net2899 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07758__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold353 top.CPU.registers.data\[458\] vssd1 vssd1 vccd1 vccd1 net2910 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold364 top.CPU.registers.data\[25\] vssd1 vssd1 vccd1 vccd1 net2921 sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 top.CPU.registers.data\[802\] vssd1 vssd1 vccd1 vccd1 net2932 sky130_fd_sc_hd__dlygate4sd3_1
Xhold386 top.CPU.registers.data\[51\] vssd1 vssd1 vccd1 vccd1 net2943 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout684_A _03336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout800 net804 vssd1 vssd1 vccd1 vccd1 net800 sky130_fd_sc_hd__clkbuf_4
Xhold397 top.CPU.registers.data\[19\] vssd1 vssd1 vccd1 vccd1 net2954 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout811 net812 vssd1 vssd1 vccd1 vccd1 net811 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09936_ _05564_ _05573_ _05574_ vssd1 vssd1 vccd1 vccd1 _05575_ sky130_fd_sc_hd__a21oi_2
Xfanout822 _03204_ vssd1 vssd1 vccd1 vccd1 net822 sky130_fd_sc_hd__clkbuf_4
Xfanout833 net834 vssd1 vssd1 vccd1 vccd1 net833 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1012_X net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout844 net846 vssd1 vssd1 vccd1 vccd1 net844 sky130_fd_sc_hd__clkbuf_4
Xfanout855 net858 vssd1 vssd1 vccd1 vccd1 net855 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11306__B2 _06084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout866 net870 vssd1 vssd1 vccd1 vccd1 net866 sky130_fd_sc_hd__clkbuf_2
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09867_ _04060_ _05299_ _05505_ _03650_ vssd1 vssd1 vccd1 vccd1 _05506_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout472_X net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout851_A net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout877 _03201_ vssd1 vssd1 vccd1 vccd1 net877 sky130_fd_sc_hd__buf_4
Xfanout888 net889 vssd1 vssd1 vccd1 vccd1 net888 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11029__D net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1020 top.CPU.registers.data\[855\] vssd1 vssd1 vccd1 vccd1 net3577 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout899 _03408_ vssd1 vssd1 vccd1 vccd1 net899 sky130_fd_sc_hd__buf_2
Xhold1031 top.CPU.registers.data\[793\] vssd1 vssd1 vccd1 vccd1 net3588 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11166__X _06645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08722__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1042 top.CPU.registers.data\[840\] vssd1 vssd1 vccd1 vccd1 net3599 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1053 top.CPU.registers.data\[361\] vssd1 vssd1 vccd1 vccd1 net3610 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09291__B net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08818_ net1366 _04449_ _04448_ top.CPU.control_unit.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 _04457_ sky130_fd_sc_hd__o211a_1
XFILLER_85_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1064 top.CPU.registers.data\[935\] vssd1 vssd1 vccd1 vccd1 net3621 sky130_fd_sc_hd__dlygate4sd3_1
X_09798_ top.CPU.registers.data\[826\] net1335 net867 top.CPU.registers.data\[794\]
+ net710 vssd1 vssd1 vccd1 vccd1 _05437_ sky130_fd_sc_hd__o221a_1
X_14014__184 clknet_leaf_150_clk vssd1 vssd1 vccd1 vccd1 net1653 sky130_fd_sc_hd__inv_2
X_13873__43 clknet_leaf_183_clk vssd1 vssd1 vccd1 vccd1 net1512 sky130_fd_sc_hd__inv_2
Xhold1075 top.CPU.registers.data\[592\] vssd1 vssd1 vccd1 vccd1 net3632 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1086 top.CPU.registers.data\[853\] vssd1 vssd1 vccd1 vccd1 net3643 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1097 top.CPU.registers.data\[657\] vssd1 vssd1 vccd1 vccd1 net3654 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11326__B _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15082__Q top.I2C.output_state\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08749_ net1366 _04381_ _04387_ vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__o21a_1
XFILLER_73_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout737_X net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1381_X net1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09132__C1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11760_ _06597_ net498 net193 net3062 vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__a22o_1
XFILLER_42_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10711_ _06141_ _06325_ vssd1 vssd1 vccd1 vccd1 _06326_ sky130_fd_sc_hd__nand2_1
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11490__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07694__C1 net1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11691_ _06515_ net204 net166 net3557 vssd1 vssd1 vccd1 vccd1 _01861_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout904_X net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12438__A net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13033__S net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10642_ _06258_ _06259_ vssd1 vssd1 vccd1 vccd1 _06260_ sky130_fd_sc_hd__nand2_1
X_13430_ net3568 _02861_ net120 vssd1 vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__mux2_1
XFILLER_167_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12034__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13361_ net670 net890 _02888_ _02889_ vssd1 vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__a31o_1
X_10573_ _04465_ _06152_ _04397_ vssd1 vssd1 vccd1 vccd1 _06194_ sky130_fd_sc_hd__a21oi_1
XFILLER_167_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14671__841 clknet_leaf_179_clk vssd1 vssd1 vccd1 vccd1 net2310 sky130_fd_sc_hd__inv_2
X_15100_ net1482 _01313_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r2_prev\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_77_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07997__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12312_ net2577 _03575_ net1196 vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__mux2_1
XFILLER_154_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13292_ top.mmio.mem_data_i\[9\] top.mmio.mem_data_i\[11\] vssd1 vssd1 vccd1 vccd1
+ _02835_ sky130_fd_sc_hd__nand2_1
X_16080_ net2414 _02290_ net1106 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[880\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09199__C1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15031_ clknet_leaf_91_clk _01276_ net1270 vssd1 vssd1 vccd1 vccd1 top.SPI.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_142_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12243_ net2871 net136 net433 vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__mux2_1
XANTENNA__13534__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10392__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12742__A0 net1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14712__882 clknet_leaf_169_clk vssd1 vssd1 vccd1 vccd1 net2351 sky130_fd_sc_hd__inv_2
XANTENNA__07749__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08410__A1 top.CPU.control_unit.instruction\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12174_ top.CPU.registers.data\[65\] net655 _06749_ vssd1 vssd1 vccd1 vccd1 _06855_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__10405__B _06033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13556__X _03000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11125_ net486 net462 _06620_ net302 net2849 vssd1 vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__a32o_1
XFILLER_110_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12901__A top.CPU.alu.program_counter\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07554__X _03193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09482__A _05120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15933_ net2267 _02143_ net1113 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[733\]
+ sky130_fd_sc_hd__dfrtp_1
X_11056_ net3218 net368 _06586_ net487 vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__a22o_1
XFILLER_114_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11848__A2 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10007_ _05644_ _05645_ net383 vssd1 vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__mux2_1
XANTENNA__09371__C1 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15864_ net2198 _02074_ net1150 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[664\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_18_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07921__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15795_ net2129 _02005_ net1177 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[595\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09123__C1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11958_ _06505_ net342 net229 net3269 vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__a22o_1
X_10909_ _06498_ vssd1 vssd1 vccd1 vccd1 _06499_ sky130_fd_sc_hd__inv_2
XANTENNA__11481__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11889_ _06311_ net3188 net188 vssd1 vssd1 vccd1 vccd1 _01674_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1000 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16416_ clknet_leaf_56_clk net2603 net1141 vssd1 vssd1 vccd1 vccd1 top.I2C.I2C_state\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08229__A1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13628_ net3118 top.CPU.alu.program_counter\[0\] net663 vssd1 vssd1 vccd1 vccd1 _02562_
+ sky130_fd_sc_hd__mux2_1
XFILLER_158_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09426__B1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12025__A2 net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08037__S net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10036__A1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16347_ clknet_leaf_67_clk _02556_ net1168 vssd1 vssd1 vccd1 vccd1 top.CPU.addressnew\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13559_ _03137_ _06389_ net583 _03001_ vssd1 vssd1 vccd1 vccd1 _03002_ sky130_fd_sc_hd__o211a_1
XFILLER_121_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07988__B1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09657__A _04020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16278_ clknet_leaf_43_clk _02488_ net1123 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.toreg\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15229_ net1563 _01439_ net1119 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_172_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11536__A1 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08937__C1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08401__A1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15167__Q top.CPU.registers.data_out_r1_prev\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10315__B net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout129 _07121_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__buf_2
X_07982_ net952 _03615_ _03617_ _03620_ vssd1 vssd1 vccd1 vccd1 _03621_ sky130_fd_sc_hd__a31o_1
XFILLER_99_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09721_ net609 _05356_ _05357_ _05358_ _05359_ vssd1 vssd1 vccd1 vccd1 _05360_ sky130_fd_sc_hd__o32a_1
XFILLER_86_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11839__A2 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08165__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09362__C1 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09652_ _04093_ _04124_ vssd1 vssd1 vccd1 vccd1 _05291_ sky130_fd_sc_hd__nand2_1
XANTENNA__07624__B net1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10331__A net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07912__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08603_ top.CPU.registers.data\[847\] net1375 net974 top.CPU.registers.data\[879\]
+ net1281 vssd1 vssd1 vccd1 vccd1 _04242_ sky130_fd_sc_hd__o221a_1
XANTENNA__12564__A_N _06410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09583_ net951 _05221_ vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__or2_1
XFILLER_94_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09114__C1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout265_A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08534_ net675 _04164_ _04165_ vssd1 vssd1 vccd1 vccd1 _04173_ sky130_fd_sc_hd__and3_1
XFILLER_42_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13461__A1 net1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11067__A3 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09665__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08465_ top.CPU.registers.data\[177\] net1383 net988 top.CPU.registers.data\[145\]
+ net678 vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout432_A _06602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1174_A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14655__825 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 net2294 sky130_fd_sc_hd__inv_2
XANTENNA__12016__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08396_ top.CPU.registers.data_out_r2_prev\[18\] net685 net953 _04034_ vssd1 vssd1
+ vccd1 vccd1 _04035_ sky130_fd_sc_hd__o211a_1
XFILLER_137_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout220_X net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout318_X net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11775__A1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07979__B1 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12705__B _04793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout899_A _03408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09017_ net611 _04650_ _04655_ _04645_ vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__a31o_4
XANTENNA__13516__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold150 top.CPU.registers.data\[181\] vssd1 vssd1 vccd1 vccd1 net2707 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_72_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold161 top.SPI.parameters\[0\] vssd1 vssd1 vccd1 vccd1 net2718 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_72_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold172 net116 vssd1 vssd1 vccd1 vccd1 net2729 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 top.CPU.fetch.current_ra\[18\] vssd1 vssd1 vccd1 vccd1 net2740 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout687_X net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold194 top.SPI.parameters\[18\] vssd1 vssd1 vccd1 vccd1 net2751 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07600__C1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout630 _03339_ vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__buf_4
XFILLER_77_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07815__A net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout641 net644 vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__buf_6
X_09919_ _04892_ _04920_ vssd1 vssd1 vccd1 vccd1 _05558_ sky130_fd_sc_hd__nor2_1
Xfanout652 net658 vssd1 vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__buf_2
Xfanout663 net664 vssd1 vssd1 vccd1 vccd1 net663 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08156__B1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout854_X net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout674 net675 vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout685 net686 vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__buf_4
XANTENNA__13028__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12930_ _07369_ _07370_ vssd1 vssd1 vccd1 vccd1 _07372_ sky130_fd_sc_hd__nor2_1
XANTENNA__07534__B net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout696 net697 vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__clkbuf_4
XFILLER_18_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12861_ top.CPU.alu.program_counter\[21\] _03756_ _07296_ _07308_ vssd1 vssd1 vccd1
+ vccd1 _07309_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_107_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11812_ net3440 net139 _06762_ vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15580_ net1914 _01790_ net1194 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[380\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_87_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ top.CPU.alu.program_counter\[14\] _04325_ _07237_ vssd1 vssd1 vccd1 vccd1
+ _07247_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11058__A3 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10895__B _06056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11463__A0 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07550__A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09120__A2 net1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11743_ net139 net535 net498 net192 net3420 vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__a32o_1
XFILLER_30_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09408__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12007__A2 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14398__568 clknet_leaf_152_clk vssd1 vssd1 vccd1 vccd1 net2037 sky130_fd_sc_hd__inv_2
X_11674_ net460 _06491_ net235 net165 net2946 vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__a32o_1
X_16201_ net2535 _02411_ net1055 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[1001\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09959__A1 _03650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13413_ top.CPU.control_unit.instruction\[28\] _02927_ net670 vssd1 vssd1 vccd1 vccd1
+ _02462_ sky130_fd_sc_hd__mux2_1
X_10625_ _06163_ _06243_ net389 vssd1 vssd1 vccd1 vccd1 _06244_ sky130_fd_sc_hd__mux2_1
XFILLER_139_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11766__A1 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08652__Y _04291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11222__D net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16132_ net2466 _02342_ net1198 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[932\]
+ sky130_fd_sc_hd__dfrtp_1
X_10556_ _06134_ _06177_ net306 vssd1 vssd1 vccd1 vccd1 _06178_ sky130_fd_sc_hd__mux2_1
X_13344_ top.I2C.data_out\[10\] net553 _02876_ vssd1 vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__a21oi_1
XFILLER_128_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16063_ net2397 _02273_ net1222 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[863\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_170_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13275_ net3077 net594 _02734_ _02822_ vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__a31o_1
X_10487_ _06069_ _06111_ net310 vssd1 vssd1 vccd1 vccd1 _06112_ sky130_fd_sc_hd__mux2_1
X_15014_ clknet_leaf_84_clk _01259_ net1264 vssd1 vssd1 vccd1 vccd1 top.SPI.parameters\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_142_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_12_0_clk_X clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12226_ net3802 net169 _06879_ _06747_ vssd1 vssd1 vccd1 vccd1 _01448_ sky130_fd_sc_hd__a22o_1
XFILLER_135_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_166_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11946__S net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_166_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12157_ net3973 net172 _06846_ _06657_ vssd1 vssd1 vccd1 vccd1 _01484_ sky130_fd_sc_hd__a22o_1
XFILLER_78_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11108_ net573 net526 _05962_ vssd1 vssd1 vccd1 vccd1 _06612_ sky130_fd_sc_hd__and3_1
XFILLER_150_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12088_ net3948 net176 _06812_ _06623_ vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_127_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15916_ net2250 _02126_ net1075 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[716\]
+ sky130_fd_sc_hd__dfrtp_1
X_11039_ _05847_ net537 vssd1 vssd1 vccd1 vccd1 _06579_ sky130_fd_sc_hd__and2_1
XANTENNA__12494__A2 _04986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15847_ net2181 _02057_ net1201 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[647\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_94_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07731__Y _03370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15778_ net2112 _01988_ net1174 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[578\]
+ sky130_fd_sc_hd__dfrtp_1
X_14342__512 clknet_leaf_122_clk vssd1 vssd1 vccd1 vccd1 net1981 sky130_fd_sc_hd__inv_2
XANTENNA__09111__A2 net1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14639__809 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 net2278 sky130_fd_sc_hd__inv_2
XFILLER_33_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08250_ net1035 _03887_ _03860_ vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__a21oi_4
XFILLER_21_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08990__S net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10009__A1 _03755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08181_ _03819_ vssd1 vssd1 vccd1 vccd1 _03820_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xteam_08_1430 vssd1 vssd1 vccd1 vccd1 team_08_1430/HI gpio_out[15] sky130_fd_sc_hd__conb_1
XFILLER_158_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xteam_08_1441 vssd1 vssd1 vccd1 vccd1 team_08_1441/HI gpio_out[26] sky130_fd_sc_hd__conb_1
XANTENNA__13401__S net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xteam_08_1452 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] team_08_1452/LO sky130_fd_sc_hd__conb_1
Xteam_08_1463 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] team_08_1463/LO sky130_fd_sc_hd__conb_1
XFILLER_174_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07619__B top.CPU.control_unit.instruction\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_133_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10980__A2 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12182__A1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_151_Right_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07965_ net743 _03598_ _03599_ net1308 vssd1 vssd1 vccd1 vccd1 _03604_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout382_A net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09335__C1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11157__A net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09704_ top.CPU.registers.data\[249\] net1384 vssd1 vssd1 vccd1 vccd1 _05343_ sky130_fd_sc_hd__and2_1
X_13950__120 clknet_leaf_150_clk vssd1 vssd1 vccd1 vccd1 net1589 sky130_fd_sc_hd__inv_2
XFILLER_114_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07896_ net801 _03526_ _03527_ net755 vssd1 vssd1 vccd1 vccd1 _03535_ sky130_fd_sc_hd__o211a_1
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09635_ _04990_ _05057_ _05271_ _04988_ _04922_ vssd1 vssd1 vccd1 vccd1 _05274_ sky130_fd_sc_hd__a311oi_2
XANTENNA_clkbuf_leaf_4_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11693__B1 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout170_X net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13843__13 clknet_leaf_76_clk vssd1 vssd1 vccd1 vccd1 net1482 sky130_fd_sc_hd__inv_2
XANTENNA__10996__A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1291_A net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout647_A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout268_X net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1389_A net1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09566_ top.CPU.registers.data\[896\] net1293 net1005 top.CPU.registers.data\[928\]
+ net902 vssd1 vssd1 vccd1 vccd1 _05205_ sky130_fd_sc_hd__a221o_1
X_14085__255 clknet_leaf_112_clk vssd1 vssd1 vccd1 vccd1 net1724 sky130_fd_sc_hd__inv_2
XANTENNA__11163__Y _06642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09102__A2 net1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08517_ _04155_ vssd1 vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout435_X net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout814_A net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09497_ net921 _05135_ vssd1 vssd1 vccd1 vccd1 _05136_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_102_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10000__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08861__A1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08448_ net754 _04085_ _04086_ net712 vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__o211a_1
XANTENNA__08753__X _04392_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_82_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14126__296 clknet_leaf_121_clk vssd1 vssd1 vccd1 vccd1 net1765 sky130_fd_sc_hd__inv_2
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout602_X net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08379_ net701 _04016_ _04017_ _04014_ _04015_ vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__o32a_1
XFILLER_139_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11748__A1 _06230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10410_ net446 _05965_ _06037_ vssd1 vssd1 vccd1 vccd1 _06038_ sky130_fd_sc_hd__nand3_1
XFILLER_99_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08613__A1 net1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11390_ _06512_ net277 net272 net3202 vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__a22o_1
XANTENNA__08074__C1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09810__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10341_ _03789_ _05971_ _05581_ vssd1 vssd1 vccd1 vccd1 _05972_ sky130_fd_sc_hd__a21o_1
XANTENNA__10420__A1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07529__B net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07821__C1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12158__D1 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13060_ net3660 _07455_ net896 vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__mux2_1
X_10272_ net601 _05904_ _05905_ vssd1 vssd1 vccd1 vccd1 _05906_ sky130_fd_sc_hd__a21o_4
XTAP_TAPCELL_ROW_148_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12011_ top.CPU.registers.data\[155\] _06781_ vssd1 vssd1 vccd1 vccd1 _06782_ sky130_fd_sc_hd__and2_1
XANTENNA__10523__X _06147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15316__RESET_B net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1403 net1404 vssd1 vssd1 vccd1 vccd1 net1403 sky130_fd_sc_hd__buf_2
X_14783__953 clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 net2422 sky130_fd_sc_hd__inv_2
XFILLER_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07545__A net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout460 net463 vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__buf_2
XFILLER_171_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout471 net473 vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__buf_4
XFILLER_93_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout482 net497 vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_161_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout493 net497 vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__buf_2
XFILLER_65_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12476__A2 _04122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15701_ net2035 _01911_ net1215 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[501\]
+ sky130_fd_sc_hd__dfrtp_1
X_14824__994 clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 net2463 sky130_fd_sc_hd__inv_2
X_12913_ top.CPU.alu.program_counter\[27\] _05429_ vssd1 vssd1 vccd1 vccd1 _07356_
+ sky130_fd_sc_hd__or2_1
XANTENNA__09341__A2 net1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11684__B1 net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07888__C1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07551__Y _03190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15632_ net1966 _01842_ net1107 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[432\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_104_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12844_ _07293_ vssd1 vssd1 vccd1 vccd1 _07294_ sky130_fd_sc_hd__inv_2
XANTENNA__12228__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15563_ net1897 _01773_ net1058 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[363\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11514__B net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12775_ top.CPU.alu.program_counter\[13\] _07231_ net1361 vssd1 vssd1 vccd1 vccd1
+ _01176_ sky130_fd_sc_hd__mux2_1
XANTENNA__08301__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11726_ _06571_ net208 net423 net2877 vssd1 vssd1 vccd1 vccd1 _01827_ sky130_fd_sc_hd__a22o_1
X_15494_ net1828 _01704_ net1080 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[294\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11657_ _06393_ net203 net426 net3408 vssd1 vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__a22o_1
XFILLER_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10608_ net444 _06227_ _06226_ _06216_ vssd1 vssd1 vccd1 vccd1 _06228_ sky130_fd_sc_hd__o211a_2
XANTENNA__08065__C1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11588_ _06699_ _06726_ net246 net3830 vssd1 vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_127_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10411__A1 _03755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16115_ net2449 _02325_ net1197 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[915\]
+ sky130_fd_sc_hd__dfrtp_1
X_13327_ top.CPU.control_unit.instruction\[5\] _02864_ net667 vssd1 vssd1 vccd1 vccd1
+ _02439_ sky130_fd_sc_hd__mux2_1
Xhold908 top.CPU.registers.data\[240\] vssd1 vssd1 vccd1 vccd1 net3465 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07812__C1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10539_ _04159_ _04226_ net376 vssd1 vssd1 vccd1 vccd1 _06162_ sky130_fd_sc_hd__mux2_1
XFILLER_128_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold919 top.CPU.registers.data\[590\] vssd1 vssd1 vccd1 vccd1 net3476 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_170_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16046_ net2380 _02256_ net1106 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[846\]
+ sky130_fd_sc_hd__dfrtp_1
X_13258_ top.I2C.output_state\[28\] net1053 vssd1 vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__nand2_2
XFILLER_124_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08368__B1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08907__A2 net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12209_ _06743_ net233 net169 net2722 vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__a22o_1
XFILLER_111_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13189_ top.I2C.output_state\[13\] top.I2C.output_state\[22\] vssd1 vssd1 vccd1 vccd1
+ _02770_ sky130_fd_sc_hd__nor2_1
XANTENNA__10175__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13934__104 clknet_leaf_170_clk vssd1 vssd1 vccd1 vccd1 net1573 sky130_fd_sc_hd__inv_2
XFILLER_96_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire448_A _05397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07750_ net801 _03385_ _03388_ net642 vssd1 vssd1 vccd1 vccd1 _03389_ sky130_fd_sc_hd__a31o_1
XANTENNA__12467__A2 _03854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07681_ _03313_ net547 vssd1 vssd1 vccd1 vccd1 _03320_ sky130_fd_sc_hd__and2_1
XANTENNA__11675__B1 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14069__239 clknet_leaf_174_clk vssd1 vssd1 vccd1 vccd1 net1708 sky130_fd_sc_hd__inv_2
X_09420_ top.CPU.registers.data\[738\] net1383 net986 top.CPU.registers.data\[706\]
+ net911 vssd1 vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__a221o_1
XFILLER_65_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12219__A2 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07894__A2 net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11690__A3 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09351_ _04988_ _04989_ vssd1 vssd1 vccd1 vccd1 _04990_ sky130_fd_sc_hd__nor2_1
XANTENNA__11427__B1 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08302_ top.CPU.registers.data\[595\] net1324 net855 top.CPU.registers.data\[627\]
+ net748 vssd1 vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__a221o_1
X_09282_ _04891_ _04920_ vssd1 vssd1 vccd1 vccd1 _04921_ sky130_fd_sc_hd__nand2_1
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08233_ net711 _03868_ _03869_ _03870_ _03871_ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__o32a_1
XANTENNA__10608__X _06228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout130_A _06464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08164_ net695 _03801_ _03802_ vssd1 vssd1 vccd1 vccd1 _03803_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_60_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08056__C1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08225__S net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08095_ top.CPU.registers.data\[245\] net1392 net830 top.CPU.registers.data\[213\]
+ net776 vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__a221o_1
XANTENNA__10056__A net1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload70 clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 clkload70/Y sky130_fd_sc_hd__inv_16
XFILLER_109_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14470__640 clknet_leaf_125_clk vssd1 vssd1 vccd1 vccd1 net2109 sky130_fd_sc_hd__inv_2
XFILLER_173_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload81 clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 clkload81/Y sky130_fd_sc_hd__clkinv_8
Xclkload92 clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 clkload92/Y sky130_fd_sc_hd__inv_16
X_14767__937 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 net2406 sky130_fd_sc_hd__inv_2
XFILLER_133_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08359__B1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout597_A net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1304_A _03113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14511__681 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 net2150 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_89_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09571__A2 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout385_X net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08997_ top.CPU.registers.data\[585\] net1369 net965 top.CPU.registers.data\[617\]
+ net900 vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout764_A net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14808__978 clknet_leaf_168_clk vssd1 vssd1 vccd1 vccd1 net2447 sky130_fd_sc_hd__inv_2
XFILLER_75_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07948_ top.CPU.registers.data\[248\] net1390 net820 top.CPU.registers.data\[216\]
+ net771 vssd1 vssd1 vccd1 vccd1 _03587_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_3_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10469__A1 _04049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09580__A net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09323__A2 net1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11666__B1 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout931_A net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout552_X net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07879_ _03515_ _03517_ net1308 vssd1 vssd1 vccd1 vccd1 _03518_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_104_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1294_X net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08531__B1 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09618_ top.CPU.registers.data\[800\] top.CPU.registers.data\[768\] net810 vssd1
+ vssd1 vccd1 vccd1 _05257_ sky130_fd_sc_hd__mux2_1
XANTENNA__13407__B2 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10890_ net662 _05693_ _06010_ _06471_ vssd1 vssd1 vccd1 vccd1 _06488_ sky130_fd_sc_hd__and4_2
XTAP_TAPCELL_ROW_84_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11418__B1 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09087__A1 _03342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09549_ net759 _05182_ _05184_ net699 vssd1 vssd1 vccd1 vccd1 _05188_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_100_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout817_X net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12560_ _05688_ _05767_ _07064_ vssd1 vssd1 vccd1 vccd1 _07065_ sky130_fd_sc_hd__or3_1
XANTENNA__08834__A1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12091__B1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08295__C1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08483__X _04122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10641__A1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11511_ _03181_ _06726_ vssd1 vssd1 vccd1 vccd1 _06734_ sky130_fd_sc_hd__nor2_4
XANTENNA__10641__B2 _05892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12491_ _04763_ _04792_ vssd1 vssd1 vccd1 vccd1 _07000_ sky130_fd_sc_hd__nand2_1
XANTENNA__13041__S net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11442_ _05960_ net263 _06721_ vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13591__B1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11373_ _06486_ net280 net273 net3331 vssd1 vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__a22o_1
X_10324_ net413 _05940_ _05955_ vssd1 vssd1 vccd1 vccd1 _05956_ sky130_fd_sc_hd__a21o_1
X_13112_ top.SPI.command\[2\] net1410 top.SPI.paroutput\[26\] net1358 vssd1 vssd1
+ vccd1 vccd1 _02721_ sky130_fd_sc_hd__a22o_1
XFILLER_124_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09547__C1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13043_ top.SPI.parameters\[23\] top.SPI.paroutput\[15\] net1356 vssd1 vssd1 vccd1
+ vccd1 _07447_ sky130_fd_sc_hd__mux2_1
X_10255_ net386 _05704_ vssd1 vssd1 vccd1 vccd1 _05889_ sky130_fd_sc_hd__nand2_1
XANTENNA__07546__Y _03185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10157__B1 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09011__A1 net1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1200 net1205 vssd1 vssd1 vccd1 vccd1 net1200 sky130_fd_sc_hd__clkbuf_2
Xfanout1211 net1212 vssd1 vssd1 vccd1 vccd1 net1211 sky130_fd_sc_hd__buf_2
XFILLER_78_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10186_ _05820_ _05821_ net388 vssd1 vssd1 vccd1 vccd1 _05822_ sky130_fd_sc_hd__mux2_1
XANTENNA__08996__S1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11509__B _06731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1222 net1226 vssd1 vssd1 vccd1 vccd1 net1222 sky130_fd_sc_hd__buf_2
Xfanout1233 net1277 vssd1 vssd1 vccd1 vccd1 net1233 sky130_fd_sc_hd__buf_2
Xfanout1244 net1259 vssd1 vssd1 vccd1 vccd1 net1244 sky130_fd_sc_hd__buf_2
XFILLER_67_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1255 net1257 vssd1 vssd1 vccd1 vccd1 net1255 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13564__X _03005_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08770__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1266 net1276 vssd1 vssd1 vccd1 vccd1 net1266 sky130_fd_sc_hd__clkbuf_2
Xfanout1277 top.CPU.fetch.nrst vssd1 vssd1 vccd1 vccd1 net1277 sky130_fd_sc_hd__clkbuf_8
X_14994_ clknet_leaf_91_clk _01239_ net1270 vssd1 vssd1 vccd1 vccd1 top.SPI.counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11228__C net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout290 net292 vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__buf_4
Xfanout1288 net1289 vssd1 vssd1 vccd1 vccd1 net1288 sky130_fd_sc_hd__buf_2
Xfanout1299 net1301 vssd1 vssd1 vccd1 vccd1 net1299 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11657__B1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11121__A2 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload6_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11672__A3 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15615_ net1949 _01825_ net1203 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[415\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11409__B1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12827_ _07251_ _07257_ _07266_ _07265_ vssd1 vssd1 vccd1 vccd1 _07279_ sky130_fd_sc_hd__o31a_1
XANTENNA__10880__A1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11244__B net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15546_ net1880 _01756_ net1252 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[346\]
+ sky130_fd_sc_hd__dfrtp_1
X_12758_ _07185_ _07196_ _07197_ _07203_ _07194_ vssd1 vssd1 vccd1 vccd1 _07216_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_139_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11709_ _06544_ net200 net421 net2731 vssd1 vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_174_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10428__X _06056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15477_ net1811 _01687_ net1216 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[277\]
+ sky130_fd_sc_hd__dfrtp_1
X_12689_ _07152_ _07153_ vssd1 vssd1 vccd1 vccd1 _07154_ sky130_fd_sc_hd__nor2_1
XFILLER_129_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08038__C1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14454__624 clknet_leaf_176_clk vssd1 vssd1 vccd1 vccd1 net2093 sky130_fd_sc_hd__inv_2
XANTENNA__13582__A0 top.CPU.alu.program_counter\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12075__B net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09786__C1 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold705 top.CPU.fetch.current_ra\[6\] vssd1 vssd1 vccd1 vccd1 net3262 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09250__A1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold716 top.CPU.registers.data\[808\] vssd1 vssd1 vccd1 vccd1 net3273 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10935__A2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold727 top.CPU.registers.data\[238\] vssd1 vssd1 vccd1 vccd1 net3284 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold738 top.CPU.registers.data\[678\] vssd1 vssd1 vccd1 vccd1 net3295 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_170_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold749 top.CPU.registers.data\[443\] vssd1 vssd1 vccd1 vccd1 net3306 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16029_ net2363 _02239_ net1122 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[829\]
+ sky130_fd_sc_hd__dfrtp_1
X_08920_ top.CPU.registers.data\[810\] top.CPU.registers.data\[778\] net809 vssd1
+ vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__mux2_1
XFILLER_69_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09553__A2 _05190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08851_ net950 _04486_ _04489_ net624 vssd1 vssd1 vccd1 vccd1 _04490_ sky130_fd_sc_hd__a211o_1
XANTENNA__11896__B1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1405 top.CPU.handler.toreg\[26\] vssd1 vssd1 vccd1 vccd1 net3962 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11360__A2 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08761__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07802_ _03440_ vssd1 vssd1 vccd1 vccd1 _03441_ sky130_fd_sc_hd__inv_2
Xhold1416 top.CPU.registers.data\[74\] vssd1 vssd1 vccd1 vccd1 net3973 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1427 top.CPU.data_out\[24\] vssd1 vssd1 vccd1 vccd1 net3984 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1438 top.mmio.mem_data_i\[3\] vssd1 vssd1 vccd1 vccd1 net3995 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11138__C net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08782_ net789 _04412_ _04413_ net738 vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__o211a_1
XFILLER_85_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1449 top.CPU.addressnew\[3\] vssd1 vssd1 vccd1 vccd1 net4006 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09305__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07733_ net417 _03371_ vssd1 vssd1 vccd1 vccd1 _03372_ sky130_fd_sc_hd__and2_1
XANTENNA__11648__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10610__Y _06230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout178_A _06795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12030__S net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07664_ _03262_ _03278_ _03302_ vssd1 vssd1 vccd1 vccd1 _03303_ sky130_fd_sc_hd__nor3_1
XFILLER_52_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12860__A2 _03685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11663__A3 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09403_ net696 _05040_ _05041_ vssd1 vssd1 vccd1 vccd1 _05042_ sky130_fd_sc_hd__and3_1
XANTENNA__10871__A1 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07595_ top.CPU.registers.data\[31\] net865 net731 _03233_ vssd1 vssd1 vccd1 vccd1
+ _03234_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout345_A net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09334_ top.CPU.registers.data\[964\] net1329 net860 top.CPU.registers.data\[996\]
+ net726 vssd1 vssd1 vccd1 vccd1 _04973_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_62_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_892 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12073__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_531 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09265_ top.CPU.registers.data\[197\] net971 net950 _04903_ vssd1 vssd1 vccd1 vccd1
+ _04904_ sky130_fd_sc_hd__a211o_1
XANTENNA__11820__B1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_0_0_clk_X clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08292__A2 net1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08216_ _03854_ _03823_ net454 vssd1 vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__mux2_1
XANTENNA__08029__C1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09196_ top.CPU.registers.data\[38\] top.CPU.registers.data\[6\] net978 vssd1 vssd1
+ vccd1 vccd1 _04835_ sky130_fd_sc_hd__mux2_1
XFILLER_14_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14197__367 clknet_leaf_173_clk vssd1 vssd1 vccd1 vccd1 net1836 sky130_fd_sc_hd__inv_2
X_08147_ _03755_ _03784_ vssd1 vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout300_X net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1042_X net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08044__A2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload170 clknet_leaf_109_clk vssd1 vssd1 vccd1 vccd1 clkload170/Y sky130_fd_sc_hd__clkinv_8
X_08078_ _03716_ vssd1 vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__inv_2
Xclkload181 clknet_leaf_129_clk vssd1 vssd1 vccd1 vccd1 clkload181/Y sky130_fd_sc_hd__inv_12
XANTENNA_fanout881_A net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12272__Y _06887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload192 clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 clkload192/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_8_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout979_A net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1307_X net1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10040_ net632 net547 _03322_ _03311_ _03313_ vssd1 vssd1 vccd1 vccd1 _05679_ sky130_fd_sc_hd__a32oi_4
XANTENNA__11887__A0 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08201__C1 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11329__B net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold10 top.CPU.registers.data_out_r2_prev\[18\] vssd1 vssd1 vccd1 vccd1 net2567 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11351__A2 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold21 top.CPU.registers.data_out_r2_prev\[19\] vssd1 vssd1 vccd1 vccd1 net2578 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout767_X net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold32 top.CPU.registers.data_out_r1_prev\[22\] vssd1 vssd1 vccd1 vccd1 net2589 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13628__A1 top.CPU.alu.program_counter\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10801__X _06412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold43 top.CPU.registers.data_out_r2_prev\[17\] vssd1 vssd1 vccd1 vccd1 net2600 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 _00070_ vssd1 vssd1 vccd1 vccd1 net2611 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08919__A net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold65 top.CPU.registers.data_out_r1_prev\[8\] vssd1 vssd1 vccd1 vccd1 net2622 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 top.CPU.registers.data\[551\] vssd1 vssd1 vccd1 vccd1 net2633 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 net51 vssd1 vssd1 vccd1 vccd1 net2644 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11639__B1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold98 net46 vssd1 vssd1 vccd1 vccd1 net2655 sky130_fd_sc_hd__dlygate4sd3_1
X_11991_ _06554_ net341 net180 net2923 vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout934_X net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11103__A2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08504__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13036__S net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13730_ top.SPI.timem\[13\] top.SPI.timem\[14\] _03071_ vssd1 vssd1 vccd1 vccd1 _03074_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07542__B net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09701__C1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10942_ _06472_ _06517_ vssd1 vssd1 vccd1 vccd1 _06519_ sky130_fd_sc_hd__nor2_2
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_954 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11064__B net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13661_ net1353 _03152_ vssd1 vssd1 vccd1 vccd1 _03044_ sky130_fd_sc_hd__nand2_1
X_10873_ net492 net468 _06476_ net223 net2887 vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_27_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15400_ net1734 _01610_ net1077 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[200\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12612_ _07102_ _07111_ vssd1 vssd1 vccd1 vccd1 _07112_ sky130_fd_sc_hd__nand2_1
X_16380_ clknet_leaf_65_clk _02589_ net1163 vssd1 vssd1 vccd1 vccd1 top.CPU.fetch.current_ra\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12064__B1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13592_ top.CPU.addressnew\[17\] net578 _03020_ _03021_ vssd1 vssd1 vccd1 vccd1 _02547_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08654__A top.CPU.alu.program_counter\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13800__B2 top.CPU.data_out\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14141__311 clknet_leaf_133_clk vssd1 vssd1 vccd1 vccd1 net1780 sky130_fd_sc_hd__inv_2
X_15331_ net1665 _01541_ net1185 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[131\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_101_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12543_ net1397 _03251_ _03286_ _06450_ vssd1 vssd1 vccd1 vccd1 _07052_ sky130_fd_sc_hd__or4_1
XANTENNA__11811__B1 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09480__A1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14438__608 clknet_leaf_126_clk vssd1 vssd1 vccd1 vccd1 net2077 sky130_fd_sc_hd__inv_2
XANTENNA__09480__B2 _03110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10090__A2 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15262_ net1596 _01472_ net1237 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_145_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12474_ _06981_ _06982_ vssd1 vssd1 vccd1 vccd1 _06983_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_117_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_91_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13564__A0 top.CPU.alu.program_counter\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13559__X _03002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09768__C1 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11425_ _06566_ net281 net269 net2851 vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__a22o_1
XANTENNA__08035__A2 net1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15193_ net1530 _01403_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r1_prev\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12904__A top.CPU.alu.program_counter\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10378__B1 _06007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11356_ net3820 net286 net277 _06357_ vssd1 vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__a22o_1
XFILLER_113_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08991__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10307_ _05816_ _05819_ net386 vssd1 vssd1 vccd1 vccd1 _05939_ sky130_fd_sc_hd__mux2_1
XFILLER_141_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11287_ net138 _06471_ net428 vssd1 vssd1 vccd1 vccd1 _06702_ sky130_fd_sc_hd__and3_1
X_13026_ net3085 _07438_ net894 vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__mux2_1
XFILLER_117_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11878__A0 _06084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10238_ net404 net391 _05859_ _05758_ vssd1 vssd1 vccd1 vccd1 _05873_ sky130_fd_sc_hd__a31o_1
XFILLER_121_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1030 net1031 vssd1 vssd1 vccd1 vccd1 net1030 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11342__A2 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1041 net1042 vssd1 vssd1 vccd1 vccd1 net1041 sky130_fd_sc_hd__buf_4
XFILLER_67_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10169_ _05523_ _05612_ _05804_ _05805_ vssd1 vssd1 vccd1 vccd1 _05806_ sky130_fd_sc_hd__o31ai_4
Xfanout1052 _03092_ vssd1 vssd1 vccd1 vccd1 net1052 sky130_fd_sc_hd__buf_2
Xfanout1063 net1068 vssd1 vssd1 vccd1 vccd1 net1063 sky130_fd_sc_hd__buf_2
XFILLER_120_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1074 net1075 vssd1 vssd1 vccd1 vccd1 net1074 sky130_fd_sc_hd__clkbuf_4
XFILLER_94_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07733__A net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1085 net1086 vssd1 vssd1 vccd1 vccd1 net1085 sky130_fd_sc_hd__clkbuf_2
Xfanout1096 net1097 vssd1 vssd1 vccd1 vccd1 net1096 sky130_fd_sc_hd__clkbuf_4
X_14977_ clknet_leaf_94_clk _01222_ net1261 vssd1 vssd1 vccd1 vccd1 top.SPI.paroutput\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11255__A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_164_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10853__A1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_44_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08259__C1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12055__B1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10605__A1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15529_ net1863 _01739_ net1055 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[329\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_179_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09050_ top.CPU.registers.data\[328\] net1314 net845 top.CPU.registers.data\[360\]
+ net772 vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_59_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08001_ top.CPU.registers.data\[344\] net1290 net1010 top.CPU.registers.data\[376\]
+ net933 vssd1 vssd1 vccd1 vccd1 _03640_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_102_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold502 top.CPU.registers.data\[973\] vssd1 vssd1 vccd1 vccd1 net3059 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold513 top.CPU.registers.data\[113\] vssd1 vssd1 vccd1 vccd1 net3070 sky130_fd_sc_hd__dlygate4sd3_1
Xhold524 top.CPU.registers.data\[805\] vssd1 vssd1 vccd1 vccd1 net3081 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09774__A2 net1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11030__B2 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold535 top.CPU.registers.data\[721\] vssd1 vssd1 vccd1 vccd1 net3092 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12533__B _05601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07785__A1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold546 top.CPU.registers.data\[980\] vssd1 vssd1 vccd1 vccd1 net3103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 top.CPU.registers.data\[683\] vssd1 vssd1 vccd1 vccd1 net3114 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold568 top.CPU.registers.data\[311\] vssd1 vssd1 vccd1 vccd1 net3125 sky130_fd_sc_hd__dlygate4sd3_1
X_09952_ _03889_ _03918_ vssd1 vssd1 vccd1 vccd1 _05591_ sky130_fd_sc_hd__nand2_1
Xhold579 top.CPU.registers.data\[334\] vssd1 vssd1 vccd1 vccd1 net3136 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08903_ net787 _04540_ _04541_ net741 vssd1 vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__o211a_1
XANTENNA__11149__B net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_117_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09883_ _03577_ _03544_ vssd1 vssd1 vccd1 vccd1 _05522_ sky130_fd_sc_hd__nand2b_1
XFILLER_44_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_672 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout295_A _06662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11333__A2 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1202 top.CPU.registers.data\[756\] vssd1 vssd1 vccd1 vccd1 net3759 sky130_fd_sc_hd__dlygate4sd3_1
X_08834_ net926 _04471_ _04472_ net950 vssd1 vssd1 vccd1 vccd1 _04473_ sky130_fd_sc_hd__o211a_1
Xhold1213 net69 vssd1 vssd1 vccd1 vccd1 net3770 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1002_A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1224 top.CPU.registers.data\[270\] vssd1 vssd1 vccd1 vccd1 net3781 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1235 top.CPU.registers.data\[863\] vssd1 vssd1 vccd1 vccd1 net3792 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07643__A _03262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1246 top.I2C.data_out\[12\] vssd1 vssd1 vccd1 vccd1 net3803 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14582__752 clknet_leaf_179_clk vssd1 vssd1 vccd1 vccd1 net2221 sky130_fd_sc_hd__inv_2
Xhold1257 top.CPU.registers.data\[967\] vssd1 vssd1 vccd1 vccd1 net3814 sky130_fd_sc_hd__dlygate4sd3_1
X_08765_ net789 _04403_ _04402_ net718 vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__o211a_1
Xhold1268 top.CPU.registers.data_out_r1_prev\[1\] vssd1 vssd1 vccd1 vccd1 net3825
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout462_A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1279 top.CPU.registers.data\[669\] vssd1 vssd1 vccd1 vccd1 net3836 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11165__A net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07716_ top.CPU.registers.data\[255\] top.CPU.registers.data\[223\] net999 vssd1
+ vssd1 vccd1 vccd1 _03355_ sky130_fd_sc_hd__mux2_1
XANTENNA__11097__A1 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08498__C1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08696_ top.CPU.registers.data\[653\] net1312 net843 top.CPU.registers.data\[685\]
+ net714 vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__a221o_1
XFILLER_82_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07647_ _03270_ _03284_ vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__nand2_2
XFILLER_26_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout250_X net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14623__793 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 net2262 sky130_fd_sc_hd__inv_2
XFILLER_80_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout727_A net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout348_X net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1371_A net1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12046__A0 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07578_ top.CPU.registers.data\[831\] net836 vssd1 vssd1 vccd1 vccd1 _03217_ sky130_fd_sc_hd__or2_1
XANTENNA__13794__B1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09317_ _04955_ vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__inv_2
XFILLER_51_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout515_X net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1028 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09248_ net702 _04884_ _04885_ _04886_ vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__a31o_1
XFILLER_108_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09214__A1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_10_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_10_0_clk sky130_fd_sc_hd__clkbuf_8
X_09179_ top.CPU.registers.data\[582\] net1316 net848 top.CPU.registers.data\[614\]
+ net742 vssd1 vssd1 vccd1 vccd1 _04818_ sky130_fd_sc_hd__a221o_1
XFILLER_147_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13010__A2 _07429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11210_ net148 net3685 net299 vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__mux2_1
X_12190_ net564 net361 _06670_ net169 top.CPU.registers.data\[56\] vssd1 vssd1 vccd1
+ vccd1 _06862_ sky130_fd_sc_hd__a32o_1
XANTENNA__10515__Y _06139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_112_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07776__A1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11141_ net478 _06629_ vssd1 vssd1 vccd1 vccd1 _06630_ sky130_fd_sc_hd__and2_1
Xoutput44 net44 vssd1 vssd1 vccd1 vccd1 ADR_O[14] sky130_fd_sc_hd__buf_2
XANTENNA__07537__B net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10244__A _03167_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput55 net55 vssd1 vssd1 vccd1 vccd1 ADR_O[24] sky130_fd_sc_hd__buf_2
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 ADR_O[9] sky130_fd_sc_hd__buf_2
XFILLER_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 DAT_O[18] sky130_fd_sc_hd__buf_2
XFILLER_122_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11072_ net3366 net366 _06591_ net312 vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__a22o_1
Xoutput88 net88 vssd1 vssd1 vccd1 vccd1 DAT_O[28] sky130_fd_sc_hd__buf_2
Xoutput99 net99 vssd1 vssd1 vccd1 vccd1 DAT_O[9] sky130_fd_sc_hd__buf_2
XANTENNA__11324__A2 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10023_ net408 _05650_ _05661_ vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15880_ net2214 _02090_ net1099 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[680\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07553__A net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input23_A DAT_I[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11075__A _06354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11974_ _06530_ net353 net183 net3119 vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__a22o_1
XFILLER_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16501_ clknet_leaf_49_clk _02663_ net1128 vssd1 vssd1 vccd1 vccd1 top.mmio.mem_data_i\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09150__B1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13713_ net3994 _03060_ _07113_ vssd1 vssd1 vccd1 vccd1 _03063_ sky130_fd_sc_hd__o21ai_1
X_10925_ _06333_ _06472_ vssd1 vssd1 vccd1 vccd1 _06508_ sky130_fd_sc_hd__or2_1
XANTENNA__08655__Y _04294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16432_ clknet_leaf_66_clk net2796 net1166 vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12037__A0 _06230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13644_ net2737 _07262_ net665 vssd1 vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__mux2_1
X_10856_ net601 _06462_ _06463_ vssd1 vssd1 vccd1 vccd1 _06464_ sky130_fd_sc_hd__a21o_2
XANTENNA__12588__A1 top.CPU.handler.readout vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13785__B1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16363_ clknet_leaf_45_clk _02572_ net1125 vssd1 vssd1 vccd1 vccd1 top.CPU.fetch.current_ra\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13575_ net3999 net578 _03011_ vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_136_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08256__A2 net1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10787_ _06244_ _06397_ net403 vssd1 vssd1 vccd1 vccd1 _06398_ sky130_fd_sc_hd__mux2_1
XFILLER_158_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15314_ net1648 _01524_ net1101 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[114\]
+ sky130_fd_sc_hd__dfrtp_1
X_12526_ _05227_ _05265_ _07000_ _07005_ _07034_ vssd1 vssd1 vccd1 vccd1 _07035_ sky130_fd_sc_hd__o2111a_1
X_16294_ clknet_leaf_107_clk _02503_ net1248 vssd1 vssd1 vccd1 vccd1 top.CPU.data_out\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__11260__B2 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12557__C_N net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15245_ net1579 _01455_ net1066 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_157_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_132_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12457_ _03475_ _03508_ _03541_ _03575_ vssd1 vssd1 vccd1 vccd1 _06966_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_10_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11408_ _06538_ net284 net269 net2711 vssd1 vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__a22o_1
XFILLER_114_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15176_ net1513 _01386_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r1_prev\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_12388_ top.CPU.addressnew\[19\] top.CPU.addressnew\[10\] top.CPU.addressnew\[9\]
+ top.CPU.addressnew\[2\] vssd1 vssd1 vccd1 vccd1 _06926_ sky130_fd_sc_hd__and4b_1
XANTENNA__11563__A2 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11339_ net3887 net287 net280 _05991_ vssd1 vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_169_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10771__B1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09943__A _03684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09508__A2 net1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16371__RESET_B net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12512__A1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11315__A2 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08716__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14566__736 clknet_leaf_122_clk vssd1 vssd1 vccd1 vccd1 net2205 sky130_fd_sc_hd__inv_2
X_13009_ top.SPI.paroutput\[4\] _07429_ _07431_ net3438 vssd1 vssd1 vccd1 vccd1 _01210_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09662__B net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08192__A1 net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14310__480 clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 net1949 sky130_fd_sc_hd__inv_2
XFILLER_54_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11079__A1 _03190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14607__777 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 net2246 sky130_fd_sc_hd__inv_2
X_08550_ top.CPU.control_unit.instruction\[16\] _03160_ _03985_ vssd1 vssd1 vccd1
+ vccd1 _04189_ sky130_fd_sc_hd__o21a_1
X_07501_ top.SPI.percount\[2\] vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__inv_2
X_08481_ net678 _04099_ _04100_ net612 vssd1 vssd1 vccd1 vccd1 _04120_ sky130_fd_sc_hd__a31o_1
XFILLER_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08247__A2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09444__A1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10329__A _03167_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09102_ top.CPU.registers.data\[455\] net1332 net863 top.CPU.registers.data\[487\]
+ net778 vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__a221o_1
XANTENNA__13528__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09033_ top.CPU.registers.data\[584\] net1317 net848 top.CPU.registers.data\[616\]
+ net739 vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_96_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout210_A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout308_A net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold310 top.CPU.registers.data\[128\] vssd1 vssd1 vccd1 vccd1 net2867 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11003__B2 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08404__C1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold321 top.CPU.registers.data\[421\] vssd1 vssd1 vccd1 vccd1 net2878 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold332 top.CPU.fetch.current_ra\[14\] vssd1 vssd1 vccd1 vccd1 net2889 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11554__A2 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold343 top.CPU.registers.data\[60\] vssd1 vssd1 vccd1 vccd1 net2900 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold354 top.CPU.registers.data\[798\] vssd1 vssd1 vccd1 vccd1 net2911 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10064__A net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold365 top.CPU.registers.data\[579\] vssd1 vssd1 vccd1 vccd1 net2922 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold376 top.CPU.registers.data\[576\] vssd1 vssd1 vccd1 vccd1 net2933 sky130_fd_sc_hd__dlygate4sd3_1
Xhold387 top.I2C.output_state\[1\] vssd1 vssd1 vccd1 vccd1 net2944 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1217_A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold398 top.mmio.mem_data_i\[25\] vssd1 vssd1 vccd1 vccd1 net2955 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout801 net804 vssd1 vssd1 vccd1 vccd1 net801 sky130_fd_sc_hd__clkbuf_2
X_09935_ _05530_ _05540_ _05570_ _04260_ _05572_ vssd1 vssd1 vccd1 vccd1 _05574_ sky130_fd_sc_hd__a221o_1
Xfanout812 net813 vssd1 vssd1 vccd1 vccd1 net812 sky130_fd_sc_hd__buf_2
Xfanout823 net831 vssd1 vssd1 vccd1 vccd1 net823 sky130_fd_sc_hd__buf_4
XANTENNA__10999__A net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout834 net839 vssd1 vssd1 vccd1 vccd1 net834 sky130_fd_sc_hd__clkbuf_4
XFILLER_131_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout677_A net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08707__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11306__A2 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13375__A _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout845 net846 vssd1 vssd1 vccd1 vccd1 net845 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout298_X net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout856 net858 vssd1 vssd1 vccd1 vccd1 net856 sky130_fd_sc_hd__clkbuf_4
X_09866_ _05367_ _05504_ vssd1 vssd1 vccd1 vccd1 _05505_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_70_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout867 net868 vssd1 vssd1 vccd1 vccd1 net867 sky130_fd_sc_hd__buf_2
Xfanout878 net879 vssd1 vssd1 vccd1 vccd1 net878 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1005_X net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1010 top.CPU.registers.data\[740\] vssd1 vssd1 vccd1 vccd1 net3567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1021 top.CPU.registers.data\[1023\] vssd1 vssd1 vccd1 vccd1 net3578 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11857__A3 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout889 net890 vssd1 vssd1 vccd1 vccd1 net889 sky130_fd_sc_hd__clkbuf_2
XFILLER_133_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08817_ net1283 _04454_ _04455_ vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__or3_1
Xhold1032 top.CPU.registers.data\[892\] vssd1 vssd1 vccd1 vccd1 net3589 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1043 top.CPU.registers.data\[957\] vssd1 vssd1 vccd1 vccd1 net3600 sky130_fd_sc_hd__dlygate4sd3_1
X_09797_ _05432_ _05433_ vssd1 vssd1 vccd1 vccd1 _05436_ sky130_fd_sc_hd__or2_2
XANTENNA_fanout844_A net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1054 top.CPU.registers.data\[903\] vssd1 vssd1 vccd1 vccd1 net3611 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1065 top.CPU.registers.data\[834\] vssd1 vssd1 vccd1 vccd1 net3622 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout465_X net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1076 top.mmio.mem_data_i\[18\] vssd1 vssd1 vccd1 vccd1 net3633 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08748_ net1283 _04379_ _04380_ top.CPU.control_unit.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 _04387_ sky130_fd_sc_hd__o31a_1
Xhold1087 top.CPU.registers.data\[999\] vssd1 vssd1 vccd1 vccd1 net3644 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1098 top.CPU.registers.data\[659\] vssd1 vssd1 vccd1 vccd1 net3655 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11326__C net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09132__B1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08679_ top.CPU.registers.data\[718\] net1378 net981 top.CPU.registers.data\[750\]
+ net934 vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__o221a_1
XANTENNA__09683__A1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1374_X net1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10710_ net409 _06164_ _06321_ _06324_ vssd1 vssd1 vccd1 vccd1 _06325_ sky130_fd_sc_hd__a22o_1
XFILLER_42_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11690_ net466 _06514_ net239 net166 net3189 vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__a32o_1
XFILLER_13_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10641_ net548 _04603_ _05643_ _05892_ vssd1 vssd1 vccd1 vccd1 _06259_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_153_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09587__X _05226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13360_ _03107_ net670 vssd1 vssd1 vccd1 vccd1 _02889_ sky130_fd_sc_hd__nor2_1
XFILLER_166_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10572_ net3668 net228 net315 _06193_ vssd1 vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_165_Right_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12311_ net2604 _03508_ net1123 vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__mux2_1
XANTENNA__11793__A2 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13291_ top.mmio.mem_data_i\[14\] top.mmio.mem_data_i\[15\] top.mmio.mem_data_i\[13\]
+ top.mmio.mem_data_i\[12\] vssd1 vssd1 vccd1 vccd1 _02834_ sky130_fd_sc_hd__and4b_1
XANTENNA__12454__A _03241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15030_ clknet_leaf_90_clk _01275_ net1267 vssd1 vssd1 vccd1 vccd1 top.SPI.count\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_6_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12242_ net3156 _05847_ net434 vssd1 vssd1 vccd1 vccd1 _01438_ sky130_fd_sc_hd__mux2_1
XFILLER_5_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12742__A1 net1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11545__A2 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08946__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14253__423 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 net1892 sky130_fd_sc_hd__inv_2
XFILLER_174_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12173_ net3979 net174 _06854_ _06661_ vssd1 vssd1 vccd1 vccd1 _01476_ sky130_fd_sc_hd__a22o_1
XFILLER_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07835__X _03474_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11124_ net516 _06150_ vssd1 vssd1 vccd1 vccd1 _06620_ sky130_fd_sc_hd__nor2_1
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11055_ net571 net441 net132 net538 vssd1 vssd1 vccd1 vccd1 _06586_ sky130_fd_sc_hd__and4_1
XFILLER_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15932_ net2266 _02142_ net1196 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[732\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08174__A1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10006_ _04093_ _04158_ net378 vssd1 vssd1 vccd1 vccd1 _05645_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15863_ net2197 _02073_ net1180 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[663\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_92_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11236__C net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15794_ net2128 _02004_ net1098 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[594\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10808__A1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09702__S net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11957_ _06504_ net343 net229 net3356 vssd1 vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__a22o_1
XFILLER_91_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08477__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10284__A2 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10908_ _06190_ _06472_ vssd1 vssd1 vccd1 vccd1 _06498_ sky130_fd_sc_hd__or2_1
X_11888_ net144 net3274 net188 vssd1 vssd1 vccd1 vccd1 _01675_ sky130_fd_sc_hd__mux2_1
XFILLER_149_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16415_ clknet_leaf_54_clk net2616 net1141 vssd1 vssd1 vccd1 vccd1 top.I2C.I2C_state\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13627_ net1360 net1040 vssd1 vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__and2_1
XFILLER_34_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10839_ net552 _06447_ vssd1 vssd1 vccd1 vccd1 _06448_ sky130_fd_sc_hd__or2_1
XFILLER_13_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16346_ clknet_leaf_80_clk _02555_ net1241 vssd1 vssd1 vccd1 vccd1 top.CPU.addressnew\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13558_ top.CPU.alu.program_counter\[4\] net1348 vssd1 vssd1 vccd1 vccd1 _03001_
+ sky130_fd_sc_hd__or2_1
XANTENNA__11233__B2 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08634__C1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_132_Right_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07988__A1 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11784__A2 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12509_ _04362_ _04391_ net450 _04461_ _07017_ vssd1 vssd1 vccd1 vccd1 _07018_ sky130_fd_sc_hd__a221oi_1
X_16277_ clknet_leaf_33_clk _02487_ net1123 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.toreg\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13489_ top.CPU.data_out\[3\] _05018_ net587 vssd1 vssd1 vccd1 vccd1 _02501_ sky130_fd_sc_hd__mux2_1
X_13919__89 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 net1558 sky130_fd_sc_hd__inv_2
XFILLER_66_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15228_ net1562 _01438_ net1201 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11536__A2 _06290_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15159_ clknet_leaf_40_clk _01369_ net1117 vssd1 vssd1 vccd1 vccd1 top.I2C.data_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12651__X _00000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10744__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07981_ net675 _03618_ _03619_ net604 vssd1 vssd1 vccd1 vccd1 _03620_ sky130_fd_sc_hd__a31o_1
XANTENNA__12811__B _04123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09720_ net682 _05337_ _05338_ net614 vssd1 vssd1 vccd1 vccd1 _05359_ sky130_fd_sc_hd__a31o_1
XANTENNA__10171__X _05808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10612__A net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09362__B1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09651_ _05280_ _05287_ _05288_ _04194_ vssd1 vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__a211o_1
XANTENNA__16279__Q top.CPU.handler.toreg\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10969__D net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10331__B net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07912__A1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08602_ top.CPU.registers.data\[975\] net1375 net974 top.CPU.registers.data\[1007\]
+ net1364 vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__o221a_1
XFILLER_103_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09582_ top.CPU.registers.data\[480\] top.CPU.registers.data\[448\] net973 vssd1
+ vssd1 vccd1 vccd1 _05221_ sky130_fd_sc_hd__mux2_1
XANTENNA__09114__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08533_ net933 _04162_ _04163_ net953 vssd1 vssd1 vccd1 vccd1 _04172_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout160_A _06760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08468__A2 net1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13461__A2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout258_A net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10275__A2 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08464_ top.CPU.registers.data\[113\] top.CPU.registers.data\[81\] top.CPU.registers.data\[49\]
+ top.CPU.registers.data\[17\] net988 net955 vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__mux4_1
XANTENNA__08873__C1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07771__S0 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14694__864 clknet_leaf_125_clk vssd1 vssd1 vccd1 vccd1 net2333 sky130_fd_sc_hd__inv_2
X_08395_ net619 _04029_ _04031_ _04033_ vssd1 vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout425_A _06756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08625__C1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout213_X net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1334_A net1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14237__407 clknet_leaf_133_clk vssd1 vssd1 vccd1 vccd1 net1876 sky130_fd_sc_hd__inv_2
X_09016_ net950 _04651_ _04654_ net624 vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__a211o_1
XFILLER_164_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11527__A2 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout794_A _03205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold140 top.CPU.registers.data\[874\] vssd1 vssd1 vccd1 vccd1 net2697 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09050__C1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold151 top.CPU.registers.data\[310\] vssd1 vssd1 vccd1 vccd1 net2708 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_72_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold162 _01206_ vssd1 vssd1 vccd1 vccd1 net2719 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10735__B1 _06347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08898__S net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold173 top.CPU.registers.data\[398\] vssd1 vssd1 vccd1 vccd1 net2730 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09583__A net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold184 top.I2C.output_state\[25\] vssd1 vssd1 vccd1 vccd1 net2741 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 top.CPU.registers.data\[455\] vssd1 vssd1 vccd1 vccd1 net2752 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout961_A net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout620 net623 vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__buf_4
XFILLER_59_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09918_ _05543_ _05556_ vssd1 vssd1 vccd1 vccd1 _05557_ sky130_fd_sc_hd__and2_1
Xfanout642 net643 vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__buf_6
XANTENNA__12488__B1 _04633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout653 net654 vssd1 vssd1 vccd1 vccd1 net653 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout664 net666 vssd1 vssd1 vccd1 vccd1 net664 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout675 net676 vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__buf_4
XFILLER_101_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout686 _03332_ vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__buf_4
Xfanout697 net701 vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__buf_2
XFILLER_86_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09849_ net682 _05483_ _05484_ _05487_ net615 vssd1 vssd1 vccd1 vccd1 _05488_ sky130_fd_sc_hd__a311o_1
XFILLER_160_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout847_X net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12860_ top.CPU.alu.program_counter\[20\] _03685_ _03756_ top.CPU.alu.program_counter\[21\]
+ vssd1 vssd1 vccd1 vccd1 _07308_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_107_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11811_ net1401 _06652_ net236 net159 net3338 vssd1 vssd1 vccd1 vccd1 _01748_ sky130_fd_sc_hd__a32o_1
X_12791_ _07244_ _07245_ vssd1 vssd1 vccd1 vccd1 _07246_ sky130_fd_sc_hd__and2b_1
XANTENNA__08459__A2 net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13044__S net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10895__C net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11742_ net141 net536 net499 net193 net2748 vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__a32o_1
XFILLER_18_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _06035_ net3650 net166 vssd1 vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16200_ net2534 _02410_ net1098 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[1000\]
+ sky130_fd_sc_hd__dfrtp_1
X_13412_ net890 _02926_ vssd1 vssd1 vccd1 vccd1 _02927_ sky130_fd_sc_hd__and2_1
XANTENNA__09959__A2 _05367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10624_ net385 _06197_ _06242_ vssd1 vssd1 vccd1 vccd1 _06243_ sky130_fd_sc_hd__a21o_1
XFILLER_139_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_133_Left_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10423__C1 _05664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16131_ net2465 _02341_ net1206 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[931\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_154_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13343_ net1343 top.mmio.mem_data_i\[10\] net596 vssd1 vssd1 vccd1 vccd1 _02876_
+ sky130_fd_sc_hd__o21a_1
X_10555_ _04225_ _04294_ net373 vssd1 vssd1 vccd1 vccd1 _06177_ sky130_fd_sc_hd__mux2_1
XFILLER_154_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16062_ net2396 _02272_ net1202 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[862\]
+ sky130_fd_sc_hd__dfrtp_1
X_13274_ _03139_ _02734_ vssd1 vssd1 vccd1 vccd1 _02822_ sky130_fd_sc_hd__nor2_1
X_14849__1019 clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 net2488 sky130_fd_sc_hd__inv_2
X_10486_ _04021_ _04094_ net376 vssd1 vssd1 vccd1 vccd1 _06111_ sky130_fd_sc_hd__mux2_1
X_15013_ clknet_leaf_94_clk _01258_ net1261 vssd1 vssd1 vccd1 vccd1 top.SPI.parameters\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_108_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11518__A2 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12225_ top.CPU.registers.data\[38\] net649 net361 vssd1 vssd1 vccd1 vccd1 _06879_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__07565__X _03204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08395__A1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12191__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12156_ top.CPU.registers.data\[74\] net647 net244 vssd1 vssd1 vccd1 vccd1 _06846_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_166_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11107_ net494 net469 _06611_ net304 net2977 vssd1 vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__a32o_1
X_12087_ top.CPU.registers.data\[109\] net471 net360 net343 vssd1 vssd1 vccd1 vccd1
+ _06812_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_127_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_142_Left_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13140__A1 top.CPU.data_out\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09344__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15915_ net2249 _02125_ net1057 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[715\]
+ sky130_fd_sc_hd__dfrtp_1
X_11038_ net3913 net367 _06578_ net324 vssd1 vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__a22o_1
XFILLER_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08698__A2 net1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15846_ net2180 _02056_ net1081 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[646\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14381__551 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 net2020 sky130_fd_sc_hd__inv_2
X_12989_ top.SPI.busy _03135_ _07418_ vssd1 vssd1 vccd1 vccd1 _07419_ sky130_fd_sc_hd__a21oi_1
X_15777_ net2111 _01987_ net1252 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[577\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11263__A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14678__848 clknet_leaf_175_clk vssd1 vssd1 vccd1 vccd1 net2317 sky130_fd_sc_hd__inv_2
XANTENNA__12078__B net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_180_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_180_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_21_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14422__592 clknet_leaf_176_clk vssd1 vssd1 vccd1 vccd1 net2061 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_151_Left_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07887__S net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_08_1420 vssd1 vssd1 vccd1 vccd1 team_08_1420/HI gpio_oeb[6] sky130_fd_sc_hd__conb_1
X_08180_ top.CPU.registers.data_out_r1_prev\[23\] net875 _03804_ _03818_ vssd1 vssd1
+ vccd1 vccd1 _03819_ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_31_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14719__889 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 net2358 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xteam_08_1431 vssd1 vssd1 vccd1 vccd1 team_08_1431/HI gpio_out[16] sky130_fd_sc_hd__conb_1
XANTENNA__12954__A1 top.CPU.alu.program_counter\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xteam_08_1442 vssd1 vssd1 vccd1 vccd1 team_08_1442/HI gpio_out[27] sky130_fd_sc_hd__conb_1
XFILLER_9_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xteam_08_1453 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] team_08_1453/LO sky130_fd_sc_hd__conb_1
Xteam_08_1464 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] team_08_1464/LO sky130_fd_sc_hd__conb_1
X_16329_ clknet_leaf_68_clk _02538_ net1167 vssd1 vssd1 vccd1 vccd1 top.CPU.addressnew\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_145_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10717__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11390__B1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_160_Left_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07964_ top.CPU.registers.data\[856\] net1319 net850 top.CPU.registers.data\[888\]
+ net693 vssd1 vssd1 vccd1 vccd1 _03603_ sky130_fd_sc_hd__a221o_1
XFILLER_68_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09335__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09703_ top.CPU.registers.data\[89\] net1306 net1029 top.CPU.registers.data\[121\]
+ net960 vssd1 vssd1 vccd1 vccd1 _05342_ sky130_fd_sc_hd__a221o_1
XFILLER_114_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10061__B net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07895_ net801 _03530_ _03531_ net730 vssd1 vssd1 vccd1 vccd1 _03534_ sky130_fd_sc_hd__o211a_1
XFILLER_96_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout375_A net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09634_ _04988_ _05272_ vssd1 vssd1 vccd1 vccd1 _05273_ sky130_fd_sc_hd__nor2_1
XFILLER_83_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10996__B net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09565_ top.CPU.registers.data\[800\] top.CPU.registers.data\[768\] net973 vssd1
+ vssd1 vccd1 vccd1 _05204_ sky130_fd_sc_hd__mux2_1
XFILLER_83_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout542_A net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout163_X net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13434__A2 net1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1284_A net1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08516_ top.CPU.registers.data_out_r1_prev\[16\] net874 _04140_ _04154_ vssd1 vssd1
+ vccd1 vccd1 _04155_ sky130_fd_sc_hd__o211ai_4
XANTENNA__11445__B2 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09496_ top.CPU.registers.data\[673\] top.CPU.registers.data\[641\] net1000 vssd1
+ vssd1 vccd1 vccd1 _05135_ sky130_fd_sc_hd__mux2_1
XANTENNA__08310__A1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11996__A2 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08447_ top.CPU.registers.data\[913\] net1332 net863 top.CPU.registers.data\[945\]
+ net729 vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_65_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout330_X net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_171_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_171_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08861__A2 _04497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout807_A net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout428_X net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11901__A net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13833__3 clknet_leaf_157_clk vssd1 vssd1 vccd1 vccd1 net1472 sky130_fd_sc_hd__inv_2
X_08378_ net792 _04008_ _04009_ net744 vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__o211a_1
XANTENNA__11748__A2 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09271__C1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10517__A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1337_X net1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10340_ _03723_ _05970_ _05582_ vssd1 vssd1 vccd1 vccd1 _05971_ sky130_fd_sc_hd__a21o_1
XFILLER_118_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout797_X net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12158__C1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10271_ top.CPU.fetch.current_ra\[26\] net1044 net883 top.CPU.handler.toreg\[26\]
+ vssd1 vssd1 vccd1 vccd1 _05905_ sky130_fd_sc_hd__a22o_1
XFILLER_117_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08377__A1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12173__A2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12010_ _05847_ net3384 net151 vssd1 vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__mux2_1
XFILLER_133_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout964_X net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11381__B1 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1404 top.CPU.control_unit.instruction\[9\] vssd1 vssd1 vccd1 vccd1 net1404
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA__11920__A2 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout461 net462 vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__clkbuf_4
Xfanout472 net473 vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12878__S net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout483 net485 vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__clkbuf_4
XFILLER_101_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout494 net496 vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__clkbuf_4
XANTENNA__15356__RESET_B net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13673__A2 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08928__Y _04567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12912_ _07348_ _07351_ vssd1 vssd1 vccd1 vccd1 _07355_ sky130_fd_sc_hd__or2_1
X_15700_ net2034 _01910_ net1112 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[500\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11684__A1 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14365__535 clknet_leaf_133_clk vssd1 vssd1 vccd1 vccd1 net2004 sky130_fd_sc_hd__inv_2
XANTENNA__07888__B1 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09252__S net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12843_ top.CPU.alu.program_counter\[19\] _03986_ _07275_ vssd1 vssd1 vccd1 vccd1
+ _07293_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_122_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15631_ net1965 _01841_ net1095 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[431\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11083__A net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15562_ net1896 _01772_ net1088 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[362\]
+ sky130_fd_sc_hd__dfrtp_1
X_12774_ _07230_ _07227_ net128 vssd1 vssd1 vccd1 vccd1 _07231_ sky130_fd_sc_hd__mux2_1
X_14406__576 clknet_leaf_123_clk vssd1 vssd1 vccd1 vccd1 net2045 sky130_fd_sc_hd__inv_2
XANTENNA__11987__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11725_ _06569_ net205 net420 net2766 vssd1 vssd1 vccd1 vccd1 _01828_ sky130_fd_sc_hd__a22o_1
X_15493_ net1827 _01703_ net1063 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[293\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_162_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_162_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11656_ _06375_ net198 net424 net3341 vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__a22o_1
XFILLER_128_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08392__A net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11739__A2 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10607_ _04468_ _05567_ vssd1 vssd1 vccd1 vccd1 _06227_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08065__B1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10427__A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09262__C1 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11587_ net495 net476 _06698_ net249 net2648 vssd1 vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__a32o_1
X_16114_ net2448 _02324_ net1108 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[914\]
+ sky130_fd_sc_hd__dfrtp_1
X_13326_ _02830_ _02863_ vssd1 vssd1 vccd1 vccd1 _02864_ sky130_fd_sc_hd__nor2_1
XFILLER_155_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10538_ net397 _06070_ vssd1 vssd1 vccd1 vccd1 _06161_ sky130_fd_sc_hd__nand2_1
Xhold909 top.CPU.registers.data\[691\] vssd1 vssd1 vccd1 vccd1 net3466 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07812__B1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16045_ net2379 _02255_ net1071 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[845\]
+ sky130_fd_sc_hd__dfrtp_1
X_13257_ net891 top.I2C.data_out\[7\] _02789_ vssd1 vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__mux2_1
XANTENNA__09014__C1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10469_ _04049_ _05677_ _05889_ _05982_ vssd1 vssd1 vccd1 vccd1 _06095_ sky130_fd_sc_hd__o22a_1
XANTENNA__13361__A1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12164__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12208_ net3849 net650 _06871_ vssd1 vssd1 vccd1 vccd1 _01458_ sky130_fd_sc_hd__o21a_1
XFILLER_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13188_ _06901_ _07119_ _02768_ vssd1 vssd1 vccd1 vccd1 _02769_ sky130_fd_sc_hd__or3_1
XANTENNA__11372__B1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_1038 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07576__C1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11258__A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11911__A2 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13973__143 clknet_leaf_174_clk vssd1 vssd1 vccd1 vccd1 net1612 sky130_fd_sc_hd__inv_2
X_12139_ net3947 net174 _06837_ _06651_ vssd1 vssd1 vccd1 vccd1 _01493_ sky130_fd_sc_hd__a22o_1
XFILLER_29_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07591__A2 net1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12788__S net1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11692__S net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11675__A1 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07680_ _03285_ net632 net547 vssd1 vssd1 vccd1 vccd1 _03319_ sky130_fd_sc_hd__and3_2
XANTENNA__07879__B1 net1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07471__A top.CPU.control_unit.instruction\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_25_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15829_ net2163 _02039_ net1211 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[629\]
+ sky130_fd_sc_hd__dfrtp_1
X_09350_ net416 _04987_ vssd1 vssd1 vccd1 vccd1 _04989_ sky130_fd_sc_hd__nor2_1
XFILLER_18_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09096__A2 net1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08301_ _03936_ _03939_ net637 vssd1 vssd1 vccd1 vccd1 _03940_ sky130_fd_sc_hd__a21o_1
XANTENNA__11978__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09281_ _04918_ _04919_ net452 vssd1 vssd1 vccd1 vccd1 _04920_ sky130_fd_sc_hd__mux2_1
XFILLER_33_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_153_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_153_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_166_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08232_ net731 _03861_ net699 vssd1 vssd1 vccd1 vccd1 _03871_ sky130_fd_sc_hd__a21o_1
XANTENNA__08506__S net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16292__Q top.CPU.data_out\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08163_ net795 _03796_ _03797_ net749 vssd1 vssd1 vccd1 vccd1 _03802_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_60_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout123_A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08094_ net798 _03732_ vssd1 vssd1 vccd1 vccd1 _03733_ sky130_fd_sc_hd__or2_1
XANTENNA__10056__B net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload60 clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 clkload60/Y sky130_fd_sc_hd__clkinv_16
XANTENNA__11867__S net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload71 clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 clkload71/Y sky130_fd_sc_hd__inv_12
Xclkload82 clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 clkload82/X sky130_fd_sc_hd__clkbuf_8
XFILLER_162_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload93 clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 clkload93/Y sky130_fd_sc_hd__inv_16
XANTENNA__12155__A2 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09020__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout492_A net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11902__A2 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13903__73 clknet_leaf_192_clk vssd1 vssd1 vccd1 vccd1 net1542 sky130_fd_sc_hd__inv_2
X_14052__222 clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 net1691 sky130_fd_sc_hd__inv_2
X_08996_ top.CPU.registers.data\[681\] top.CPU.registers.data\[649\] top.CPU.registers.data\[553\]
+ top.CPU.registers.data\[521\] net965 net901 vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__mux4_1
XFILLER_130_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07582__A2 net1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14349__519 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 net1988 sky130_fd_sc_hd__inv_2
X_07947_ top.CPU.registers.data\[184\] top.CPU.registers.data\[152\] net820 vssd1
+ vssd1 vccd1 vccd1 _03586_ sky130_fd_sc_hd__mux2_1
XFILLER_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout280_X net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11115__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout757_A net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07652__Y _03291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11666__A1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07878_ net755 _03512_ _03516_ net700 vssd1 vssd1 vccd1 vccd1 _03517_ sky130_fd_sc_hd__o211a_1
XFILLER_141_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09617_ top.CPU.registers.data\[640\] net1313 net844 top.CPU.registers.data\[672\]
+ net715 vssd1 vssd1 vccd1 vccd1 _05256_ sky130_fd_sc_hd__a221o_1
XANTENNA__11174__Y _06648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout545_X net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout924_A net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14848__1018 clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 net2487 sky130_fd_sc_hd__inv_2
XANTENNA_fanout1287_X net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09548_ net803 _05185_ _05186_ net731 vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__o211a_1
XANTENNA__08819__C1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11969__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09479_ net695 _05113_ _05114_ _05117_ vssd1 vssd1 vccd1 vccd1 _05118_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_144_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_144_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout712_X net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09492__C1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11510_ _06466_ _06603_ _06731_ vssd1 vssd1 vccd1 vccd1 _06733_ sky130_fd_sc_hd__or3_4
XFILLER_156_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12490_ net449 _04727_ vssd1 vssd1 vccd1 vccd1 _06999_ sky130_fd_sc_hd__nor2_1
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08047__B1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11441_ net3069 net263 vssd1 vssd1 vccd1 vccd1 _06721_ sky130_fd_sc_hd__nand2_1
XFILLER_137_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09244__C1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14750__920 clknet_leaf_152_clk vssd1 vssd1 vccd1 vccd1 net2389 sky130_fd_sc_hd__inv_2
XFILLER_50_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11372_ _06485_ net279 net272 net3498 vssd1 vssd1 vccd1 vccd1 _02138_ sky130_fd_sc_hd__a22o_1
X_13111_ net3877 _02720_ _07422_ vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__mux2_1
X_10323_ _05793_ _05945_ _05684_ _05761_ vssd1 vssd1 vccd1 vccd1 _05955_ sky130_fd_sc_hd__a211oi_1
XANTENNA__13558__A top.CPU.alu.program_counter\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12462__A net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09547__B1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13957__127 clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 net1596 sky130_fd_sc_hd__inv_2
XFILLER_140_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13042_ net3672 _07446_ net894 vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__mux2_1
X_10254_ _05666_ _05887_ vssd1 vssd1 vccd1 vccd1 _05888_ sky130_fd_sc_hd__nand2_1
XANTENNA__08151__S net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15537__RESET_B net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11354__B1 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1201 net1204 vssd1 vssd1 vccd1 vccd1 net1201 sky130_fd_sc_hd__clkbuf_4
Xfanout1212 net1218 vssd1 vssd1 vccd1 vccd1 net1212 sky130_fd_sc_hd__clkbuf_4
X_10185_ _05713_ _05719_ net307 vssd1 vssd1 vccd1 vccd1 _05821_ sky130_fd_sc_hd__mux2_1
Xfanout1223 net1225 vssd1 vssd1 vccd1 vccd1 net1223 sky130_fd_sc_hd__clkbuf_4
Xfanout1234 net1235 vssd1 vssd1 vccd1 vccd1 net1234 sky130_fd_sc_hd__clkbuf_4
Xfanout1245 net1259 vssd1 vssd1 vccd1 vccd1 net1245 sky130_fd_sc_hd__clkbuf_4
XFILLER_94_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1256 net1257 vssd1 vssd1 vccd1 vccd1 net1256 sky130_fd_sc_hd__clkbuf_4
Xfanout1267 net1275 vssd1 vssd1 vccd1 vccd1 net1267 sky130_fd_sc_hd__clkbuf_4
X_14993_ clknet_leaf_92_clk _01238_ net1269 vssd1 vssd1 vccd1 vccd1 top.SPI.counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1278 _03146_ vssd1 vssd1 vccd1 vccd1 net1278 sky130_fd_sc_hd__buf_2
Xfanout280 net281 vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__clkbuf_4
Xfanout291 net292 vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__buf_6
Xfanout1289 net1292 vssd1 vssd1 vccd1 vccd1 net1289 sky130_fd_sc_hd__clkbuf_4
XFILLER_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12826_ _07277_ vssd1 vssd1 vccd1 vccd1 _07278_ sky130_fd_sc_hd__inv_2
X_15614_ net1948 _01824_ net1239 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[414\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10880__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09710__S net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12757_ _07213_ _07214_ vssd1 vssd1 vccd1 vccd1 _07215_ sky130_fd_sc_hd__or2_1
X_15545_ net1879 _01755_ net1223 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[345\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12637__A top.I2C.output_state\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_135_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_135_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_139_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11541__A _06373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11708_ _06542_ net205 net422 net2783 vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_139_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15476_ net1810 _01686_ net1119 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[276\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_174_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12688_ top.CPU.alu.program_counter\[5\] _07142_ vssd1 vssd1 vccd1 vccd1 _07153_
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_42_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08038__B1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11639_ _06011_ net203 net426 net3416 vssd1 vssd1 vccd1 vccd1 _01912_ sky130_fd_sc_hd__a22o_1
X_14493__663 clknet_leaf_133_clk vssd1 vssd1 vccd1 vccd1 net2132 sky130_fd_sc_hd__inv_2
XANTENNA__13582__A1 _06210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10396__A1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold706 top.CPU.registers.data\[258\] vssd1 vssd1 vccd1 vccd1 net3263 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_3_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold717 top.CPU.registers.data\[265\] vssd1 vssd1 vccd1 vccd1 net3274 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07797__C1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13309_ top.I2C.data_out\[1\] net553 _02850_ vssd1 vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__a21oi_1
Xhold728 top.CPU.registers.data\[881\] vssd1 vssd1 vccd1 vccd1 net3285 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold739 top.CPU.registers.data\[117\] vssd1 vssd1 vccd1 vccd1 net3296 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12137__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07466__A top.CPU.alu.program_counter\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14036__206 clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 net1675 sky130_fd_sc_hd__inv_2
X_16028_ net2362 _02238_ net1234 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[828\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_112_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11345__B1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15278__RESET_B net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08210__B1 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08850_ _04487_ _04488_ net673 vssd1 vssd1 vccd1 vccd1 _04489_ sky130_fd_sc_hd__o21a_1
XANTENNA__10699__A2 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15207__RESET_B net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07801_ _03439_ _03409_ net453 vssd1 vssd1 vccd1 vccd1 _03440_ sky130_fd_sc_hd__mux2_1
Xhold1406 top.CPU.registers.data\[75\] vssd1 vssd1 vccd1 vccd1 net3963 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1417 top.CPU.addressnew\[13\] vssd1 vssd1 vccd1 vccd1 net3974 sky130_fd_sc_hd__dlygate4sd3_1
X_08781_ net789 _04416_ _04417_ net718 vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__o211a_1
XFILLER_85_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1428 top.SPI.timem\[12\] vssd1 vssd1 vccd1 vccd1 net3985 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1439 top.SPI.timem\[17\] vssd1 vssd1 vccd1 vccd1 net3996 sky130_fd_sc_hd__dlygate4sd3_1
X_07732_ _03370_ top.CPU.alu.immediate\[31\] net454 vssd1 vssd1 vccd1 vccd1 _03371_
+ sky130_fd_sc_hd__mux2_2
XFILLER_84_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08297__A net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08513__A1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07663_ _03264_ _03301_ vssd1 vssd1 vccd1 vccd1 _03302_ sky130_fd_sc_hd__nor2_1
XFILLER_1_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10320__A1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07721__C1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09402_ top.CPU.registers.data\[739\] net1391 net828 top.CPU.registers.data\[707\]
+ net727 vssd1 vssd1 vccd1 vccd1 _05041_ sky130_fd_sc_hd__a221o_1
XFILLER_164_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09069__A2 net1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07594_ top.CPU.registers.data\[63\] net836 vssd1 vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__or2_1
XANTENNA__10871__A2 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09333_ net643 _04968_ _04971_ net876 top.CPU.registers.data_out_r1_prev\[4\] vssd1
+ vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__o32a_1
XANTENNA__08277__B1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout240_A net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_126_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_126_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout338_A _03047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14734__904 clknet_leaf_121_clk vssd1 vssd1 vccd1 vccd1 net2373 sky130_fd_sc_hd__inv_2
XFILLER_166_504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09264_ top.CPU.registers.data\[229\] net1374 vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__and2_1
XANTENNA__11820__A1 net1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10249__A1_N _05499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08215_ _03838_ _03853_ vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__or2_4
XFILLER_21_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08029__B1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10067__A _04829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09195_ top.CPU.registers.data\[646\] net1287 net1013 top.CPU.registers.data\[678\]
+ net904 vssd1 vssd1 vccd1 vccd1 _04834_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout126_X net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08146_ _03784_ vssd1 vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__inv_2
XFILLER_112_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11584__B1 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07788__C1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11597__S net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08077_ _03700_ _03715_ vssd1 vssd1 vccd1 vccd1 _03716_ sky130_fd_sc_hd__or2_4
Xclkload160 clknet_leaf_112_clk vssd1 vssd1 vccd1 vccd1 clkload160/Y sky130_fd_sc_hd__inv_2
Xclkload171 clknet_leaf_110_clk vssd1 vssd1 vccd1 vccd1 clkload171/Y sky130_fd_sc_hd__inv_2
Xclkload182 clknet_leaf_83_clk vssd1 vssd1 vccd1 vccd1 clkload182/Y sky130_fd_sc_hd__clkinv_4
Xclkload193 clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 clkload193/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__09067__S net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12128__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11336__B1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15630__RESET_B net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout495_X net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout874_A net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08201__B1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold11 top.CPU.registers.data_out_r2_prev\[16\] vssd1 vssd1 vccd1 vccd1 net2568 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 top.CPU.registers.data_out_r1_prev\[3\] vssd1 vssd1 vccd1 vccd1 net2579 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold33 top.CPU.registers.data_out_r2_prev\[15\] vssd1 vssd1 vccd1 vccd1 net2590 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 top.CPU.registers.data_out_r1_prev\[25\] vssd1 vssd1 vccd1 vccd1 net2601 sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ top.CPU.registers.data_out_r1_prev\[9\] net871 net690 _04610_ _04617_ vssd1
+ vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__o2111a_1
XANTENNA_fanout662_X net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold55 top.CPU.registers.data_out_r2_prev\[31\] vssd1 vssd1 vccd1 vccd1 net2612 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07960__C1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold66 top.CPU.registers.data_out_r1_prev\[11\] vssd1 vssd1 vccd1 vccd1 net2623 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 net45 vssd1 vssd1 vccd1 vccd1 net2634 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 net44 vssd1 vssd1 vccd1 vccd1 net2645 sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ _06552_ net344 net180 net2825 vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__a22o_1
Xhold99 top.CPU.registers.data\[304\] vssd1 vssd1 vccd1 vccd1 net2656 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09701__B1 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10941_ _06517_ vssd1 vssd1 vccd1 vccd1 _06518_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout927_X net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07712__C1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13660_ _03152_ _07055_ _02823_ _03126_ vssd1 vssd1 vccd1 vccd1 _03043_ sky130_fd_sc_hd__a31o_1
XFILLER_72_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10872_ net661 _05847_ net437 vssd1 vssd1 vccd1 vccd1 _06476_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_27_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09530__S net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12611_ _07104_ _07105_ _07110_ vssd1 vssd1 vccd1 vccd1 _07111_ sky130_fd_sc_hd__nor3_1
XFILLER_45_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12064__A1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13591_ _03117_ _03137_ net578 vssd1 vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_117_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_117_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10075__A0 _04567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14180__350 clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 net1819 sky130_fd_sc_hd__inv_2
X_15330_ net1664 _01540_ net1171 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[130\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_156_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12542_ _03252_ _03313_ _06450_ _07050_ vssd1 vssd1 vccd1 vccd1 _07051_ sky130_fd_sc_hd__a31oi_2
XANTENNA__10614__A2 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11811__A1 net1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14477__647 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 net2116 sky130_fd_sc_hd__inv_2
XANTENNA__12176__B net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15261_ net1595 _01471_ net1120 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[61\]
+ sky130_fd_sc_hd__dfrtp_1
X_12473_ _04019_ _04048_ vssd1 vssd1 vccd1 vccd1 _06982_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_117_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07985__S net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07838__X _03477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13564__A1 _06352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11424_ _06564_ net275 net267 net3261 vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__a22o_1
X_14221__391 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 net1860 sky130_fd_sc_hd__inv_2
X_15192_ net1529 _01402_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r1_prev\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14518__688 clknet_leaf_180_clk vssd1 vssd1 vccd1 vccd1 net2157 sky130_fd_sc_hd__inv_2
XFILLER_165_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12904__B _05499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09485__B _05123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08440__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11355_ net3524 net287 net281 _06336_ vssd1 vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__a22o_1
XFILLER_125_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12119__A2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10306_ net401 _05616_ _05937_ vssd1 vssd1 vccd1 vccd1 _05938_ sky130_fd_sc_hd__or3_1
XANTENNA__07794__A2 net1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11286_ net530 _05693_ vssd1 vssd1 vccd1 vccd1 _06701_ sky130_fd_sc_hd__nor2_1
X_13025_ top.SPI.parameters\[14\] top.SPI.paroutput\[6\] net1355 vssd1 vssd1 vccd1
+ vccd1 _07438_ sky130_fd_sc_hd__mux2_1
XFILLER_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10237_ _05870_ _05871_ net401 vssd1 vssd1 vccd1 vccd1 _05872_ sky130_fd_sc_hd__mux2_1
XFILLER_121_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1020 net1022 vssd1 vssd1 vccd1 vccd1 net1020 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07573__X _03212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1031 net1032 vssd1 vssd1 vccd1 vccd1 net1031 sky130_fd_sc_hd__clkbuf_4
Xfanout1042 _03165_ vssd1 vssd1 vccd1 vccd1 net1042 sky130_fd_sc_hd__clkbuf_2
Xfanout1053 _07118_ vssd1 vssd1 vccd1 vccd1 net1053 sky130_fd_sc_hd__clkbuf_4
X_10168_ _05773_ _05774_ _05799_ _05803_ vssd1 vssd1 vccd1 vccd1 _05805_ sky130_fd_sc_hd__o211a_1
XFILLER_121_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10550__A1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1064 net1067 vssd1 vssd1 vccd1 vccd1 net1064 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07951__C1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13894__64 clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 net1533 sky130_fd_sc_hd__inv_2
Xfanout1075 net1111 vssd1 vssd1 vccd1 vccd1 net1075 sky130_fd_sc_hd__buf_2
XANTENNA__07733__B _03371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1086 net1110 vssd1 vssd1 vccd1 vccd1 net1086 sky130_fd_sc_hd__clkbuf_2
Xfanout1097 net1110 vssd1 vssd1 vccd1 vccd1 net1097 sky130_fd_sc_hd__buf_2
X_10099_ net417 _03407_ net374 vssd1 vssd1 vccd1 vccd1 _05737_ sky130_fd_sc_hd__mux2_1
X_14976_ clknet_leaf_98_clk _01221_ net1256 vssd1 vssd1 vccd1 vccd1 top.SPI.paroutput\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09299__A2 net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12809_ _07262_ _07259_ net128 vssd1 vssd1 vccd1 vccd1 _07263_ sky130_fd_sc_hd__mux2_1
XFILLER_37_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08259__B1 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12055__A1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_108_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_108_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13789_ net18 net1052 net887 net3939 vssd1 vssd1 vccd1 vccd1 _02670_ sky130_fd_sc_hd__a22o_1
XFILLER_96_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11271__A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15528_ net1862 _01738_ net1099 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[328\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09471__A2 net1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15459_ net1793 _01669_ net1208 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[259\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08000_ top.CPU.registers.data\[280\] net983 _03638_ vssd1 vssd1 vccd1 vccd1 _03639_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__11566__B1 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold503 top.CPU.registers.data\[467\] vssd1 vssd1 vccd1 vccd1 net3060 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11030__A2 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold514 top.CPU.registers.data\[769\] vssd1 vssd1 vccd1 vccd1 net3071 sky130_fd_sc_hd__dlygate4sd3_1
Xhold525 top.CPU.registers.data\[768\] vssd1 vssd1 vccd1 vccd1 net3082 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold536 top.CPU.registers.data\[508\] vssd1 vssd1 vccd1 vccd1 net3093 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13307__A1 _02849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11210__S net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold547 top.CPU.registers.data\[616\] vssd1 vssd1 vccd1 vccd1 net3104 sky130_fd_sc_hd__dlygate4sd3_1
X_14847__1017 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 net2486 sky130_fd_sc_hd__inv_2
Xhold558 top.SPI.paroutput\[26\] vssd1 vssd1 vccd1 vccd1 net3115 sky130_fd_sc_hd__dlygate4sd3_1
X_09951_ _05581_ _05589_ _05578_ vssd1 vssd1 vccd1 vccd1 _05590_ sky130_fd_sc_hd__o21ba_1
Xhold569 top.CPU.registers.data\[783\] vssd1 vssd1 vccd1 vccd1 net3126 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11318__B1 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08902_ top.CPU.registers.data\[746\] net1387 net809 top.CPU.registers.data\[714\]
+ net765 vssd1 vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__a221o_1
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09882_ _03310_ _03320_ vssd1 vssd1 vccd1 vccd1 _05521_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_55_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08833_ top.CPU.registers.data\[683\] net1370 net966 top.CPU.registers.data\[651\]
+ net901 vssd1 vssd1 vccd1 vccd1 _04472_ sky130_fd_sc_hd__a221o_1
XFILLER_100_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1203 top.I2C.data_out\[20\] vssd1 vssd1 vccd1 vccd1 net3760 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1214 top.CPU.registers.data\[746\] vssd1 vssd1 vccd1 vccd1 net3771 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout190_A net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1225 top.CPU.registers.data\[234\] vssd1 vssd1 vccd1 vccd1 net3782 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout288_A _06712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11446__A _03193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1236 top.CPU.registers.data\[591\] vssd1 vssd1 vccd1 vccd1 net3793 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10350__A net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1247 top.CPU.registers.data\[765\] vssd1 vssd1 vccd1 vccd1 net3804 sky130_fd_sc_hd__dlygate4sd3_1
X_08764_ top.CPU.registers.data\[556\] top.CPU.registers.data\[524\] net815 vssd1
+ vssd1 vccd1 vccd1 _04403_ sky130_fd_sc_hd__mux2_1
Xhold1258 net94 vssd1 vssd1 vccd1 vccd1 net3815 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1269 top.CPU.registers.data\[749\] vssd1 vssd1 vccd1 vccd1 net3826 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07715_ top.CPU.registers.data\[159\] net1382 net999 top.CPU.registers.data\[191\]
+ net959 vssd1 vssd1 vccd1 vccd1 _03354_ sky130_fd_sc_hd__o221a_1
XANTENNA__11165__B net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12294__A1 _04361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11097__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08695_ top.CPU.registers.data\[909\] net1311 net842 top.CPU.registers.data\[941\]
+ net714 vssd1 vssd1 vccd1 vccd1 _04334_ sky130_fd_sc_hd__a221o_1
XANTENNA__09695__C1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11880__S net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07646_ _03271_ _03283_ vssd1 vssd1 vccd1 vccd1 _03285_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_146_Right_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08755__A _04363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14164__334 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 net1803 sky130_fd_sc_hd__inv_2
XFILLER_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07577_ net779 _03214_ _03215_ net756 vssd1 vssd1 vccd1 vccd1 _03216_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout243_X net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout622_A net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1364_A net1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09998__A0 _04225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09316_ top.CPU.control_unit.instruction\[11\] net1048 _04953_ _04954_ vssd1 vssd1
+ vccd1 vccd1 _04955_ sky130_fd_sc_hd__a22o_2
XANTENNA__10057__B1 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14205__375 clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 net1844 sky130_fd_sc_hd__inv_2
XFILLER_139_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09247_ net690 _04882_ _04883_ net635 vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout410_X net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1152_X net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout508_X net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13546__A1 top.CPU.done vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09178_ top.CPU.registers.data\[550\] top.CPU.registers.data\[518\] net815 vssd1
+ vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout991_A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15811__RESET_B net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11557__B1 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08129_ top.CPU.registers.data\[437\] top.CPU.registers.data\[405\] top.CPU.registers.data\[309\]
+ top.CPU.registers.data\[277\] net993 net917 vssd1 vssd1 vccd1 vccd1 _03768_ sky130_fd_sc_hd__mux4_1
XANTENNA__10084__X _05722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15129__RESET_B net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11140_ net514 _06292_ vssd1 vssd1 vccd1 vccd1 _06629_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_112_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput45 net45 vssd1 vssd1 vccd1 vccd1 ADR_O[15] sky130_fd_sc_hd__buf_2
XFILLER_162_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10244__B _05878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11309__B1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout877_X net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput56 net56 vssd1 vssd1 vccd1 vccd1 ADR_O[25] sky130_fd_sc_hd__buf_2
XFILLER_134_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput67 net1347 vssd1 vssd1 vccd1 vccd1 CYC_O sky130_fd_sc_hd__buf_2
XFILLER_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 DAT_O[19] sky130_fd_sc_hd__buf_2
X_11071_ _06311_ net534 vssd1 vssd1 vccd1 vccd1 _06591_ sky130_fd_sc_hd__and2_1
Xoutput89 net89 vssd1 vssd1 vccd1 vccd1 DAT_O[29] sky130_fd_sc_hd__buf_2
XFILLER_49_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10022_ _05652_ _05656_ _05660_ net395 net408 vssd1 vssd1 vccd1 vccd1 _05661_ sky130_fd_sc_hd__a221o_1
XFILLER_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input16_A DAT_I[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11075__B net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11973_ _06529_ net346 net181 net3229 vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__a22o_1
XANTENNA__09686__C1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16500_ clknet_leaf_49_clk _02662_ net1128 vssd1 vssd1 vccd1 vccd1 top.mmio.mem_data_i\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09150__A1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13712_ top.SPI.timem\[7\] top.SPI.timem\[8\] _03058_ vssd1 vssd1 vccd1 vccd1 _03062_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_158_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10924_ net482 net458 _06507_ net220 net3130 vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__a32o_1
XFILLER_45_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_113_Right_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16431_ clknet_leaf_55_clk _00013_ net1141 vssd1 vssd1 vccd1 vccd1 top.I2C.I2C_state\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13643_ net2884 _07249_ net665 vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__mux2_1
X_10855_ top.CPU.fetch.current_ra\[0\] net1041 net634 top.CPU.handler.toreg\[0\] vssd1
+ vssd1 vccd1 vccd1 _06463_ sky130_fd_sc_hd__a22o_1
XFILLER_72_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09438__C1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10048__B1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11091__A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13574_ _03137_ _06268_ net583 _03010_ vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__o211a_1
X_16362_ clknet_leaf_31_clk _02571_ net1126 vssd1 vssd1 vccd1 vccd1 top.CPU.fetch.current_ra\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10786_ net398 _06323_ _06396_ vssd1 vssd1 vccd1 vccd1 _06397_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_136_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09453__A2 net1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08110__C1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_171_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12525_ net449 _04727_ _04890_ _04918_ _07004_ vssd1 vssd1 vccd1 vccd1 _07034_ sky130_fd_sc_hd__o221a_1
X_15313_ net1647 _01523_ net1189 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[113\]
+ sky130_fd_sc_hd__dfrtp_1
X_16293_ clknet_leaf_108_clk _02502_ net1246 vssd1 vssd1 vccd1 vccd1 top.CPU.data_out\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_12_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11260__A2 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12915__A top.CPU.alu.program_counter\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12456_ _03405_ _03439_ _06962_ _06964_ vssd1 vssd1 vccd1 vccd1 _06965_ sky130_fd_sc_hd__o211a_1
X_15244_ net1578 _01454_ net1078 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09205__A2 net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11407_ _06537_ net282 net269 net3204 vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__a22o_1
X_15175_ net1512 _01385_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r1_prev\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_12387_ _06923_ _06924_ vssd1 vssd1 vccd1 vccd1 _06925_ sky130_fd_sc_hd__or2_1
XFILLER_4_550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11338_ net3483 net285 net278 _05963_ vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__a22o_1
XFILLER_125_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_169_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11269_ net519 _06560_ vssd1 vssd1 vccd1 vccd1 _06692_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_37_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08177__C1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13008_ top.SPI.paroutput\[3\] _07429_ _07431_ net2683 vssd1 vssd1 vccd1 vccd1 _01209_
+ sky130_fd_sc_hd__a22o_1
XFILLER_39_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10523__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11720__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07924__C1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11266__A net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12276__A1 _03474_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11079__A2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14959_ clknet_leaf_87_clk _01204_ net1271 vssd1 vssd1 vccd1 vccd1 top.SPI.csx sky130_fd_sc_hd__dfstp_1
XANTENNA__13473__B1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12796__S net1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09677__C1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14148__318 clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 net1787 sky130_fd_sc_hd__inv_2
X_07500_ top.SPI.count\[3\] vssd1 vssd1 vccd1 vccd1 _03140_ sky130_fd_sc_hd__inv_2
XFILLER_35_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08480_ net943 _04097_ _04098_ net958 vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__o211a_1
XFILLER_63_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09170__S net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11205__S net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_28_Left_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09101_ top.CPU.registers.data\[423\] top.CPU.registers.data\[391\] net832 vssd1
+ vssd1 vccd1 vccd1 _04740_ sky130_fd_sc_hd__mux2_1
XANTENNA__11787__B1 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10329__B _05960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08652__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13420__S net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09032_ top.CPU.registers.data\[552\] top.CPU.registers.data\[520\] net811 vssd1
+ vssd1 vccd1 vccd1 _04671_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_96_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15293__RESET_B net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1035 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11003__A2 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold300 top.CPU.registers.data\[370\] vssd1 vssd1 vccd1 vccd1 net2857 sky130_fd_sc_hd__dlygate4sd3_1
Xhold311 top.CPU.registers.data\[167\] vssd1 vssd1 vccd1 vccd1 net2868 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08404__B1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout203_A net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold322 top.CPU.registers.data\[588\] vssd1 vssd1 vccd1 vccd1 net2879 sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 top.SPI.paroutput\[24\] vssd1 vssd1 vccd1 vccd1 net2890 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08955__A1 _04593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07758__A2 net1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold344 top.CPU.registers.data\[842\] vssd1 vssd1 vccd1 vccd1 net2901 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold355 top.CPU.registers.data\[447\] vssd1 vssd1 vccd1 vccd1 net2912 sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 top.CPU.registers.data\[171\] vssd1 vssd1 vccd1 vccd1 net2923 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold377 top.CPU.registers.data\[18\] vssd1 vssd1 vccd1 vccd1 net2934 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold388 top.CPU.registers.data\[603\] vssd1 vssd1 vccd1 vccd1 net2945 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout802 net803 vssd1 vssd1 vccd1 vccd1 net802 sky130_fd_sc_hd__clkbuf_4
X_09934_ _05530_ _05537_ _05566_ vssd1 vssd1 vccd1 vccd1 _05573_ sky130_fd_sc_hd__and3_1
Xhold399 top.CPU.registers.data\[386\] vssd1 vssd1 vccd1 vccd1 net2956 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout813 _03204_ vssd1 vssd1 vccd1 vccd1 net813 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1112_A net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08168__C1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout824 net831 vssd1 vssd1 vccd1 vccd1 net824 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_37_Left_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout835 net836 vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__clkbuf_4
Xfanout846 net854 vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__clkbuf_4
X_09865_ _05436_ _05503_ vssd1 vssd1 vccd1 vccd1 _05504_ sky130_fd_sc_hd__or2_1
XANTENNA_input8_A DAT_I[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout857 net858 vssd1 vssd1 vccd1 vccd1 net857 sky130_fd_sc_hd__clkbuf_4
Xhold1000 top.CPU.registers.data\[451\] vssd1 vssd1 vccd1 vccd1 net3557 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout193_X net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout572_A net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11711__B1 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout868 net870 vssd1 vssd1 vccd1 vccd1 net868 sky130_fd_sc_hd__clkbuf_2
Xfanout879 _03198_ vssd1 vssd1 vccd1 vccd1 net879 sky130_fd_sc_hd__buf_2
Xhold1011 top.CPU.handler.toreg\[4\] vssd1 vssd1 vccd1 vccd1 net3568 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07915__C1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08183__A2 _03819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1022 top.CPU.registers.data\[535\] vssd1 vssd1 vccd1 vccd1 net3579 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1033 top.CPU.registers.data\[501\] vssd1 vssd1 vccd1 vccd1 net3590 sky130_fd_sc_hd__dlygate4sd3_1
X_08816_ top.CPU.registers.data\[588\] net1371 net977 top.CPU.registers.data\[620\]
+ net904 vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__o221a_1
XFILLER_86_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09796_ _05432_ _05433_ vssd1 vssd1 vccd1 vccd1 _05435_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_29_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1044 top.CPU.registers.data\[594\] vssd1 vssd1 vccd1 vccd1 net3601 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1055 top.CPU.registers.data\[931\] vssd1 vssd1 vccd1 vccd1 net3612 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1066 top.CPU.registers.data\[1001\] vssd1 vssd1 vccd1 vccd1 net3623 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07930__A2 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_90_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13464__A0 top.CPU.handler.toreg\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12267__A1 _06391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08747_ net1366 _04382_ _04385_ _03116_ vssd1 vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__o211a_1
Xhold1077 top.CPU.registers.data\[944\] vssd1 vssd1 vccd1 vccd1 net3634 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout360_X net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1088 top.CPU.registers.data\[844\] vssd1 vssd1 vccd1 vccd1 net3645 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1099 top.CPU.registers.data\[714\] vssd1 vssd1 vccd1 vccd1 net3656 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09668__C1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10278__A0 _05332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout837_A net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout458_X net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08678_ net908 _04314_ _04316_ net1368 vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__a211o_1
XFILLER_27_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09080__S net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07629_ net1398 _03259_ vssd1 vssd1 vccd1 vccd1 _03268_ sky130_fd_sc_hd__nand2_1
XFILLER_54_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12019__A1 _05960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11490__A2 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08891__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout625_X net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1367_X net1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_46_Left_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10640_ _04601_ net503 _05685_ _04602_ net443 vssd1 vssd1 vccd1 vccd1 _06258_ sky130_fd_sc_hd__o221a_1
XFILLER_13_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_153_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11778__B1 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10571_ net527 _06192_ vssd1 vssd1 vccd1 vccd1 _06193_ sky130_fd_sc_hd__nor2_1
XANTENNA__12735__A top.CPU.alu.program_counter\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09840__C1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12310_ net2592 _03439_ net1240 vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__mux2_1
XFILLER_158_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07997__A2 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13290_ top.mmio.mem_data_i\[1\] top.mmio.mem_data_i\[3\] top.mmio.mem_data_i\[2\]
+ top.mmio.mem_data_i\[0\] vssd1 vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__or4b_1
XFILLER_155_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08424__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout994_X net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12454__B _03369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09199__A1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12241_ net3167 _05808_ net432 vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__mux2_1
XANTENNA__10255__A net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_163_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14292__462 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 net1931 sky130_fd_sc_hd__inv_2
X_12172_ top.CPU.registers.data\[66\] net651 net245 vssd1 vssd1 vccd1 vccd1 _06854_
+ sky130_fd_sc_hd__o21a_1
X_14589__759 clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 net2228 sky130_fd_sc_hd__inv_2
XFILLER_122_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11950__B1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11123_ net487 net465 _06619_ net303 net3285 vssd1 vssd1 vccd1 vccd1 _02291_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_55_Left_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_43_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12470__A net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08159__C1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15931_ net2265 _02141_ net1208 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[731\]
+ sky130_fd_sc_hd__dfrtp_1
X_14918__1088 clknet_leaf_123_clk vssd1 vssd1 vccd1 vccd1 net2557 sky130_fd_sc_hd__inv_2
X_11054_ net3513 net366 _06585_ net324 vssd1 vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__a22o_1
XFILLER_104_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_178_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11702__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10005_ _03958_ _04020_ net378 vssd1 vssd1 vccd1 vccd1 _05644_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09371__A1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15862_ net2196 _02072_ net1228 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[662\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_97_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_58_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13864__34 clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 net1503 sky130_fd_sc_hd__inv_2
XANTENNA__07921__A2 net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12258__A1 _06212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13455__B1 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15793_ net2127 _02003_ net1177 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[593\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09123__A1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_101_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11956_ _06503_ net344 net229 net3437 vssd1 vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__a22o_1
XANTENNA__08331__C1 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14846__1016 clknet_leaf_153_clk vssd1 vssd1 vccd1 vccd1 net2485 sky130_fd_sc_hd__inv_2
XFILLER_33_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10907_ net481 net458 _06496_ net220 net2886 vssd1 vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__a32o_1
XANTENNA__08882__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11887_ net145 net3304 net188 vssd1 vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__mux2_1
XANTENNA__11481__A2 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16414_ clknet_leaf_56_clk net2614 net1141 vssd1 vssd1 vccd1 vccd1 top.I2C.I2C_state\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13626_ net2659 _03041_ net581 vssd1 vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__mux2_1
X_10838_ net601 _06445_ _06446_ vssd1 vssd1 vccd1 vccd1 _06447_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_15_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09426__A2 net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_116_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11769__B1 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16345_ clknet_leaf_68_clk _02554_ net1168 vssd1 vssd1 vccd1 vccd1 top.CPU.addressnew\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11233__A2 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13557_ net4006 _03000_ net580 vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__mux2_1
X_10769_ _06219_ _06380_ net400 vssd1 vssd1 vccd1 vccd1 _06381_ sky130_fd_sc_hd__mux2_1
XANTENNA__10717__X _06332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10441__A0 _03683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12508_ _04222_ _04255_ _04291_ _04324_ vssd1 vssd1 vccd1 vccd1 _07017_ sky130_fd_sc_hd__a22o_1
XANTENNA__07739__A net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16276_ clknet_leaf_44_clk _02486_ net1124 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.toreg\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13488_ top.CPU.data_out\[2\] _05084_ net590 vssd1 vssd1 vccd1 vccd1 _02500_ sky130_fd_sc_hd__mux2_1
XANTENNA__08334__S net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14533__703 clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 net2172 sky130_fd_sc_hd__inv_2
XFILLER_145_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12439_ net1341 top.I2C.output_state\[6\] net2926 vssd1 vssd1 vccd1 vccd1 _06956_
+ sky130_fd_sc_hd__a21oi_1
X_15227_ net1561 _01437_ net1215 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12194__B1 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08398__C1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11536__A3 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15158_ clknet_leaf_44_clk _01368_ net1124 vssd1 vssd1 vccd1 vccd1 top.I2C.data_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_153_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11941__B1 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07980_ top.CPU.registers.data\[248\] net1378 net983 top.CPU.registers.data\[216\]
+ net907 vssd1 vssd1 vccd1 vccd1 _03619_ sky130_fd_sc_hd__a221o_1
X_15089_ net1471 _01302_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r2_prev\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07474__A net1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12497__B2 _05265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09650_ _05280_ _05287_ _05288_ vssd1 vssd1 vccd1 vccd1 _05289_ sky130_fd_sc_hd__a21oi_1
XFILLER_110_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08570__C1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08601_ net617 _04232_ _04238_ _04239_ vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__o22a_1
X_09581_ net676 _05217_ _05219_ net902 vssd1 vssd1 vccd1 vccd1 _05220_ sky130_fd_sc_hd__o211a_1
XANTENNA__12249__A1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08532_ top.CPU.registers.data\[240\] top.CPU.registers.data\[208\] net983 vssd1
+ vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__mux2_1
XANTENNA__16295__Q top.CPU.data_out\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08463_ top.CPU.registers.data\[337\] net1296 net1016 top.CPU.registers.data\[369\]
+ net949 vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__a221o_1
XANTENNA__08873__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout153_A net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07771__S1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08394_ net626 _04032_ net616 vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__a21o_1
XFILLER_10_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10059__B _03185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout320_A net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08625__B1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12555__A top.CPU.done vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09822__C1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_30_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07979__A2 net1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10432__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11775__A3 net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14276__446 clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 net1915 sky130_fd_sc_hd__inv_2
X_09015_ _04652_ _04653_ net672 vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__o21a_1
XANTENNA__10983__B2 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout206_X net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1327_A _03109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold130 net107 vssd1 vssd1 vccd1 vccd1 net2687 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07936__X _03575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09050__B1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold141 top.CPU.registers.data\[300\] vssd1 vssd1 vccd1 vccd1 net2698 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14020__190 clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 net1659 sky130_fd_sc_hd__inv_2
XANTENNA__10735__A1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold152 top.CPU.registers.data\[548\] vssd1 vssd1 vccd1 vccd1 net2709 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_72_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11932__B1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout787_A net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold163 top.CPU.registers.data\[430\] vssd1 vssd1 vccd1 vccd1 net2720 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13386__A _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold174 top.CPU.registers.data\[434\] vssd1 vssd1 vccd1 vccd1 net2731 sky130_fd_sc_hd__dlygate4sd3_1
X_14317__487 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 net1956 sky130_fd_sc_hd__inv_2
Xhold185 top.SPI.paroutput\[19\] vssd1 vssd1 vccd1 vccd1 net2742 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07600__A1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold196 top.CPU.registers.data\[900\] vssd1 vssd1 vccd1 vccd1 net2753 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout610 net611 vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__buf_4
Xfanout621 net623 vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__buf_4
Xfanout632 _03291_ vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__buf_2
X_09917_ _04991_ _05545_ _05554_ _04987_ net412 vssd1 vssd1 vccd1 vccd1 _05556_ sky130_fd_sc_hd__a32o_1
Xfanout643 net644 vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__clkbuf_8
Xfanout654 net658 vssd1 vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__buf_2
XANTENNA_fanout954_A net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout575_X net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout665 net666 vssd1 vssd1 vccd1 vccd1 net665 sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_97_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_97_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08156__A2 net1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout676 _03336_ vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_146_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout687 _03332_ vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__clkbuf_8
X_09848_ net945 _05485_ _05486_ net960 vssd1 vssd1 vccd1 vccd1 _05487_ sky130_fd_sc_hd__o211a_1
Xfanout698 net699 vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11160__B2 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08561__C1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout742_X net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ net939 _05415_ _05417_ net956 vssd1 vssd1 vccd1 vccd1 _05418_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_107_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11558__A_N _06731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11810_ net1402 _06651_ net238 net157 net2985 vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__a32o_1
X_12790_ top.CPU.alu.program_counter\[15\] _04256_ vssd1 vssd1 vccd1 vccd1 _07245_
+ sky130_fd_sc_hd__nand2_1
XFILLER_15_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_87_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08313__C1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11999__B1 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _06586_ net238 net194 net3055 vssd1 vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__a22o_1
XFILLER_15_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08864__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11672_ net517 _06488_ net204 net167 net3061 vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_120_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09408__A2 net1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13411_ top.I2C.data_out\[28\] net555 _02925_ net598 vssd1 vssd1 vccd1 vccd1 _02926_
+ sky130_fd_sc_hd__a22o_1
X_10623_ net385 _06241_ vssd1 vssd1 vccd1 vccd1 _06242_ sky130_fd_sc_hd__nor2_1
XFILLER_169_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09813__C1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13060__S net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_21_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_155_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13342_ top.CPU.control_unit.instruction\[9\] _02875_ net667 vssd1 vssd1 vccd1 vccd1
+ _02443_ sky130_fd_sc_hd__mux2_1
X_16130_ net2464 _02340_ net1171 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[930\]
+ sky130_fd_sc_hd__dfrtp_1
X_10554_ _04330_ _06153_ vssd1 vssd1 vccd1 vccd1 _06176_ sky130_fd_sc_hd__nand2_1
XANTENNA__11766__A3 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12184__B net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10974__B2 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13273_ net3926 _02814_ _02821_ net1053 vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__a22o_1
XFILLER_127_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16061_ net2395 _02271_ net1114 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[861\]
+ sky130_fd_sc_hd__dfrtp_1
X_10485_ net395 _06022_ vssd1 vssd1 vccd1 vccd1 _06110_ sky130_fd_sc_hd__nand2_1
XFILLER_5_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07993__S net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15012_ clknet_leaf_100_clk _01257_ net1255 vssd1 vssd1 vccd1 vccd1 top.SPI.parameters\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_12224_ net477 _06692_ _06878_ net170 net3393 vssd1 vssd1 vccd1 vccd1 _01449_ sky130_fd_sc_hd__a32o_1
XFILLER_151_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11923__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09592__A1 top.CPU.control_unit.instruction\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12155_ net3963 net172 _06845_ _06656_ vssd1 vssd1 vccd1 vccd1 _01485_ sky130_fd_sc_hd__a22o_1
XFILLER_64_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_166_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10272__X _05906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11106_ _05933_ net531 net575 vssd1 vssd1 vccd1 vccd1 _06611_ sky130_fd_sc_hd__and3b_1
X_12086_ net3993 net647 _06811_ vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__o21a_1
XANTENNA__13676__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_88_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_88_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_127_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09344__A1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15914_ net2248 _02124_ net1084 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[714\]
+ sky130_fd_sc_hd__dfrtp_1
X_11037_ _05808_ net536 vssd1 vssd1 vccd1 vccd1 _06578_ sky130_fd_sc_hd__and2_1
X_15845_ net2179 _02055_ net1062 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[645\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_64_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15776_ net2110 _01986_ net1091 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[576\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_64_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12988_ _03135_ _06945_ vssd1 vssd1 vccd1 vccd1 _07418_ sky130_fd_sc_hd__nor2_2
XANTENNA__12100__B1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11939_ net135 net3480 net231 vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__mux2_1
XFILLER_33_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13609_ net2982 net579 _03031_ _03032_ vssd1 vssd1 vccd1 vccd1 _02553_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_31_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xteam_08_1421 vssd1 vssd1 vccd1 vccd1 team_08_1421/HI gpio_oeb[7] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_31_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xteam_08_1432 vssd1 vssd1 vccd1 vccd1 team_08_1432/HI gpio_out[17] sky130_fd_sc_hd__conb_1
Xclkbuf_leaf_12_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_8
Xteam_08_1443 vssd1 vssd1 vccd1 vccd1 team_08_1443/HI gpio_out[28] sky130_fd_sc_hd__conb_1
X_16328_ clknet_leaf_80_clk _02537_ net1241 vssd1 vssd1 vccd1 vccd1 top.CPU.addressnew\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12954__A2 _03409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07469__A net1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_08_1454 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] team_08_1454/LO sky130_fd_sc_hd__conb_1
XANTENNA__08064__S net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_08_1465 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] team_08_1465/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_93_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16259_ clknet_leaf_28_clk _02469_ net1149 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.toreg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_14004__174 clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 net1643 sky130_fd_sc_hd__inv_2
XFILLER_145_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11914__B1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12182__A3 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10623__A net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07963_ top.CPU.registers.data\[600\] net1319 net850 top.CPU.registers.data\[632\]
+ net704 vssd1 vssd1 vccd1 vccd1 _03602_ sky130_fd_sc_hd__a221o_1
XANTENNA__13667__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07635__C net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09702_ top.CPU.registers.data\[57\] top.CPU.registers.data\[25\] net1001 vssd1 vssd1
+ vccd1 vccd1 _05341_ sky130_fd_sc_hd__mux2_1
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07894_ top.CPU.registers.data\[348\] net1338 net870 top.CPU.registers.data\[380\]
+ net778 vssd1 vssd1 vccd1 vccd1 _03533_ sky130_fd_sc_hd__a221o_1
XFILLER_96_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11142__B2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14661__831 clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 net2300 sky130_fd_sc_hd__inv_2
XANTENNA__08543__C1 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09633_ _04990_ _05057_ _05271_ vssd1 vssd1 vccd1 vccd1 _05272_ sky130_fd_sc_hd__and3_1
XANTENNA__12890__A1 top.CPU.alu.program_counter\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10769__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11693__A2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout368_A net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11454__A net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09564_ top.CPU.registers.data\[960\] net1293 net1005 top.CPU.registers.data\[992\]
+ net902 vssd1 vssd1 vccd1 vccd1 _05203_ sky130_fd_sc_hd__a221o_1
XFILLER_83_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08515_ _04151_ _04153_ net644 vssd1 vssd1 vccd1 vccd1 _04154_ sky130_fd_sc_hd__a21o_1
XANTENNA__07649__A1 _03152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14702__872 clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 net2341 sky130_fd_sc_hd__inv_2
XANTENNA__11445__A2 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09495_ top.CPU.registers.data\[545\] top.CPU.registers.data\[513\] net1000 vssd1
+ vssd1 vccd1 vccd1 _05134_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout156_X net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout535_A net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08446_ top.CPU.registers.data\[817\] top.CPU.registers.data\[785\] net832 vssd1
+ vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1030 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08377_ net792 _04012_ _04013_ net720 vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout323_X net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout702_A net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14917__1087 clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 net2556 sky130_fd_sc_hd__inv_2
XFILLER_23_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11748__A3 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10517__B _06139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10009__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12158__B1 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09594__A _05232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10270_ _05852_ _05903_ _05902_ _05882_ vssd1 vssd1 vccd1 vccd1 _05904_ sky130_fd_sc_hd__a211o_1
XANTENNA__16443__RESET_B net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout692_X net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11905__B1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13370__A2 _07089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14845__1015 clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 net2484 sky130_fd_sc_hd__inv_2
XANTENNA__11381__A1 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08782__C1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1405 net1407 vssd1 vssd1 vccd1 vccd1 net1405 sky130_fd_sc_hd__buf_4
Xfanout440 net441 vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09326__A1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout957_X net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13122__A2 net1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout462 net463 vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__clkbuf_4
Xfanout473 _03193_ vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__buf_4
XFILLER_19_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout484 net485 vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout495 net496 vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_161_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12911_ top.CPU.alu.program_counter\[26\] _07354_ net1362 vssd1 vssd1 vccd1 vccd1
+ _01189_ sky130_fd_sc_hd__mux2_1
XFILLER_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13055__S net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15630_ net1964 _01840_ net1105 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[430\]
+ sky130_fd_sc_hd__dfrtp_1
X_12842_ _07291_ vssd1 vssd1 vccd1 vccd1 _07292_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_122_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11083__B _05694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15561_ net1895 _01771_ net1055 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[361\]
+ sky130_fd_sc_hd__dfrtp_1
X_12773_ _07228_ _07229_ vssd1 vssd1 vccd1 vccd1 _07230_ sky130_fd_sc_hd__nor2_1
XANTENNA__08837__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11724_ _06568_ net204 net422 net3109 vssd1 vssd1 vccd1 vccd1 _01829_ sky130_fd_sc_hd__a22o_1
X_15492_ net1826 _01702_ net1219 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[292\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08673__A net1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11655_ _06357_ net201 net425 net3724 vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__a22o_1
XFILLER_80_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10606_ _05643_ _05824_ _06223_ _06225_ vssd1 vssd1 vccd1 vccd1 _06226_ sky130_fd_sc_hd__o211a_1
XFILLER_127_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09262__B1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11586_ _06697_ net280 net246 net2671 vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__a22o_1
XFILLER_167_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10427__B _06054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10947__B2 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16113_ net2447 _02323_ net1190 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[913\]
+ sky130_fd_sc_hd__dfrtp_1
X_10537_ _06159_ _06157_ _04260_ vssd1 vssd1 vccd1 vccd1 _06160_ sky130_fd_sc_hd__mux2_1
X_13325_ top.I2C.data_out\[5\] net553 _02862_ vssd1 vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__a21oi_1
XFILLER_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16044_ net2378 _02254_ net1069 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[844\]
+ sky130_fd_sc_hd__dfrtp_1
X_10468_ net549 _05297_ net509 _05296_ _06093_ vssd1 vssd1 vccd1 vccd1 _06094_ sky130_fd_sc_hd__o221a_1
X_13256_ net3878 _02805_ _02812_ _02803_ vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__a22o_1
XANTENNA__09014__B1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08368__A2 net1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13361__A2 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12207_ net564 net365 _06678_ net169 top.CPU.registers.data\[48\] vssd1 vssd1 vccd1
+ vccd1 _06871_ sky130_fd_sc_hd__a32o_1
X_13187_ top.I2C.output_state\[2\] top.I2C.byte_manager_state\[2\] vssd1 vssd1 vccd1
+ vccd1 _02768_ sky130_fd_sc_hd__nand2_1
X_10399_ net414 _06025_ _06027_ net224 _06020_ vssd1 vssd1 vccd1 vccd1 _06028_ sky130_fd_sc_hd__o221a_2
XFILLER_123_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07576__B1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10175__A2 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12138_ top.CPU.registers.data\[83\] net651 net244 vssd1 vssd1 vccd1 vccd1 _06837_
+ sky130_fd_sc_hd__o21a_1
XFILLER_123_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14645__815 clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 net2284 sky130_fd_sc_hd__inv_2
X_12069_ top.CPU.registers.data\[119\] net651 vssd1 vssd1 vccd1 vccd1 _06804_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_1_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08525__C1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15828_ net2162 _02038_ net1074 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[628\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_53_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11427__A2 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15759_ net2093 _01969_ net1104 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[559\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08300_ net695 _03937_ _03938_ vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_47_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09280_ top.CPU.control_unit.instruction\[25\] _04596_ _04597_ vssd1 vssd1 vccd1
+ vccd1 _04919_ sky130_fd_sc_hd__o21a_1
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08231_ net798 _03866_ _03867_ net753 vssd1 vssd1 vccd1 vccd1 _03870_ sky130_fd_sc_hd__o211a_1
XFILLER_166_719 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08162_ net795 _03790_ _03791_ net724 vssd1 vssd1 vccd1 vccd1 _03801_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_60_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08093_ top.CPU.registers.data\[181\] top.CPU.registers.data\[149\] net830 vssd1
+ vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__mux2_1
XANTENNA__10056__C net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload50 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 clkload50/Y sky130_fd_sc_hd__inv_8
XFILLER_118_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09618__S net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload61 clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 clkload61/Y sky130_fd_sc_hd__clkinv_1
XFILLER_161_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload72 clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 clkload72/Y sky130_fd_sc_hd__inv_6
Xclkload83 clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 clkload83/Y sky130_fd_sc_hd__clkinv_4
XFILLER_115_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload94 clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 clkload94/Y sky130_fd_sc_hd__inv_16
XANTENNA__08359__A2 net1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11449__A net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07567__B1 net1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1025_A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14091__261 clknet_leaf_148_clk vssd1 vssd1 vccd1 vccd1 net1730 sky130_fd_sc_hd__inv_2
XFILLER_134_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08995_ top.CPU.alu.program_counter\[9\] _04633_ net1033 vssd1 vssd1 vccd1 vccd1
+ _04634_ sky130_fd_sc_hd__mux2_4
XFILLER_76_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_10_Left_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09308__A1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout485_A net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14388__558 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 net2027 sky130_fd_sc_hd__inv_2
XFILLER_69_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07946_ top.CPU.registers.data\[88\] net1321 net852 top.CPU.registers.data\[120\]
+ net770 vssd1 vssd1 vccd1 vccd1 _03585_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_143_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11115__A1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09353__S net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11455__Y _06726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07877_ top.CPU.registers.data\[668\] net1338 net870 top.CPU.registers.data\[700\]
+ net730 vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout273_X net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout652_A net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1394_A net1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11184__A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08531__A2 net1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09616_ top.CPU.registers.data\[544\] top.CPU.registers.data\[512\] net810 vssd1
+ vssd1 vccd1 vccd1 _05255_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14429__599 clknet_leaf_130_clk vssd1 vssd1 vccd1 vccd1 net2068 sky130_fd_sc_hd__inv_2
XFILLER_141_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11418__A2 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout440_X net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09547_ top.CPU.registers.data\[321\] net1334 net866 top.CPU.registers.data\[353\]
+ net780 vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__a221o_1
XFILLER_93_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout538_X net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout917_A net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09589__A net1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08295__A1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09478_ net748 _05115_ _05116_ net707 vssd1 vssd1 vccd1 vccd1 _05117_ sky130_fd_sc_hd__o211a_1
XANTENNA__12091__A2 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08429_ top.CPU.registers.data\[465\] net1326 net857 top.CPU.registers.data\[497\]
+ net774 vssd1 vssd1 vccd1 vccd1 _04068_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout705_X net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload0 clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clkload0/Y sky130_fd_sc_hd__inv_8
X_11440_ net567 net494 _06581_ _06720_ vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_22_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09244__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10929__B2 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08598__A2 net1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13591__A2 _03137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11371_ net494 net476 _06484_ net274 net2835 vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__a32o_1
XFILLER_164_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13110_ top.SPI.command\[1\] net1410 top.SPI.paroutput\[25\] net1357 vssd1 vssd1
+ vccd1 vccd1 _02720_ sky130_fd_sc_hd__a22o_1
X_10322_ _03648_ _05685_ _05947_ _05952_ _05953_ vssd1 vssd1 vccd1 vccd1 _05954_ sky130_fd_sc_hd__o2111ai_1
XFILLER_3_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09528__S net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12462__B _05428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13996__166 clknet_leaf_191_clk vssd1 vssd1 vccd1 vccd1 net1635 sky130_fd_sc_hd__inv_2
X_14332__502 clknet_leaf_139_clk vssd1 vssd1 vccd1 vccd1 net1971 sky130_fd_sc_hd__inv_2
X_13041_ top.SPI.parameters\[22\] top.SPI.paroutput\[14\] net1355 vssd1 vssd1 vccd1
+ vccd1 _07446_ sky130_fd_sc_hd__mux2_1
XFILLER_4_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10253_ _05738_ _05886_ net391 vssd1 vssd1 vccd1 vccd1 _05887_ sky130_fd_sc_hd__mux2_1
XFILLER_152_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07556__B net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10157__A2 _05793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10184_ _05819_ vssd1 vssd1 vccd1 vccd1 _05820_ sky130_fd_sc_hd__inv_2
Xfanout1202 net1204 vssd1 vssd1 vccd1 vccd1 net1202 sky130_fd_sc_hd__clkbuf_2
Xfanout1213 net1214 vssd1 vssd1 vccd1 vccd1 net1213 sky130_fd_sc_hd__clkbuf_4
XFILLER_132_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1224 net1225 vssd1 vssd1 vccd1 vccd1 net1224 sky130_fd_sc_hd__clkbuf_4
Xfanout1235 net1236 vssd1 vssd1 vccd1 vccd1 net1235 sky130_fd_sc_hd__clkbuf_4
Xfanout1246 net1249 vssd1 vssd1 vccd1 vccd1 net1246 sky130_fd_sc_hd__clkbuf_4
XFILLER_120_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08770__A2 net1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10550__X _06173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1257 net1258 vssd1 vssd1 vccd1 vccd1 net1257 sky130_fd_sc_hd__buf_2
X_14992_ clknet_leaf_98_clk _01237_ net1256 vssd1 vssd1 vccd1 vccd1 top.SPI.paroutput\[31\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1268 net1275 vssd1 vssd1 vccd1 vccd1 net1268 sky130_fd_sc_hd__clkbuf_4
Xfanout270 _06716_ vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__buf_4
XANTENNA__08507__C1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1279 _03145_ vssd1 vssd1 vccd1 vccd1 net1279 sky130_fd_sc_hd__clkbuf_4
Xfanout281 net284 vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__buf_4
Xfanout292 _06700_ vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__clkbuf_8
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11657__A2 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11094__A net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09180__C1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08522__A2 net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07730__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15613_ net1947 _01823_ net1119 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[413\]
+ sky130_fd_sc_hd__dfrtp_1
X_12825_ _07275_ _07276_ vssd1 vssd1 vccd1 vccd1 _07277_ sky130_fd_sc_hd__or2_1
XANTENNA__11409__A2 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12918__A top.CPU.alu.program_counter\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11244__D net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15544_ net1878 _01754_ net1101 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[344\]
+ sky130_fd_sc_hd__dfrtp_1
X_12756_ top.CPU.alu.program_counter\[12\] _04462_ vssd1 vssd1 vccd1 vccd1 _07214_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__12082__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11290__A0 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11541__B net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11707_ _06540_ net201 net421 net3032 vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_139_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15475_ net1809 _01685_ net1191 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[275\]
+ sky130_fd_sc_hd__dfrtp_1
X_12687_ top.CPU.alu.program_counter\[5\] _07142_ vssd1 vssd1 vccd1 vccd1 _07152_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_42_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09235__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11638_ _05991_ net205 net426 net3889 vssd1 vssd1 vccd1 vccd1 _01913_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_42_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13940__110 clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 net1579 sky130_fd_sc_hd__inv_2
XFILLER_129_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09786__A1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12653__A net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11569_ net2842 net246 _06743_ net481 vssd1 vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__a22o_1
XANTENNA__07797__B1 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold707 top.CPU.fetch.current_ra\[9\] vssd1 vssd1 vccd1 vccd1 net3264 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold718 top.CPU.fetch.current_ra\[13\] vssd1 vssd1 vccd1 vccd1 net3275 sky130_fd_sc_hd__dlygate4sd3_1
X_13308_ net1343 top.mmio.mem_data_i\[1\] net596 vssd1 vssd1 vccd1 vccd1 _02850_ sky130_fd_sc_hd__o21a_1
Xhold729 top.CPU.registers.data\[505\] vssd1 vssd1 vccd1 vccd1 net3286 sky130_fd_sc_hd__dlygate4sd3_1
X_16027_ net2361 _02237_ net1214 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[827\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11269__A net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14075__245 clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 net1714 sky130_fd_sc_hd__inv_2
X_13239_ top.I2C.which_data_address\[0\] _02772_ vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__and2_4
XFILLER_41_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10173__A net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11896__A2 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08761__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07800_ net683 _03432_ _03438_ _03416_ _03426_ vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__a32o_4
Xhold1407 top.CPU.registers.data\[96\] vssd1 vssd1 vccd1 vccd1 net3964 sky130_fd_sc_hd__dlygate4sd3_1
X_08780_ top.CPU.registers.data\[332\] net1316 net847 top.CPU.registers.data\[364\]
+ net762 vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_88_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1418 top.I2C.output_state\[6\] vssd1 vssd1 vccd1 vccd1 net3975 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_127_Right_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10901__A net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14116__286 clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 net1755 sky130_fd_sc_hd__inv_2
Xhold1429 top.CPU.handler.toreg\[25\] vssd1 vssd1 vccd1 vccd1 net3986 sky130_fd_sc_hd__dlygate4sd3_1
X_14916__1086 clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 net2555 sky130_fd_sc_hd__inv_2
X_07731_ _03369_ vssd1 vssd1 vccd1 vccd1 _03370_ sky130_fd_sc_hd__inv_2
XFILLER_78_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11648__A2 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10112__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07662_ top.CPU.control_unit.instruction\[14\] net1398 vssd1 vssd1 vccd1 vccd1 _03301_
+ sky130_fd_sc_hd__nand2_1
XFILLER_37_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10320__A2 _03650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09401_ top.CPU.registers.data\[579\] net1328 net859 top.CPU.registers.data\[611\]
+ net751 vssd1 vssd1 vccd1 vccd1 _05040_ sky130_fd_sc_hd__a221o_1
XFILLER_52_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07593_ net802 _03227_ _03228_ _03231_ vssd1 vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__o31a_1
XANTENNA__11291__X _06704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08277__A1 net1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09332_ net752 _04969_ _04970_ net708 vssd1 vssd1 vccd1 vccd1 _04971_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_62_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14844__1014 clknet_leaf_139_clk vssd1 vssd1 vccd1 vccd1 net2483 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_62_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12073__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09263_ top.CPU.registers.data\[165\] net1370 net966 top.CPU.registers.data\[133\]
+ net672 vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__a221o_1
X_14773__943 clknet_leaf_173_clk vssd1 vssd1 vccd1 vccd1 net2412 sky130_fd_sc_hd__inv_2
XFILLER_33_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12039__S net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout233_A net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08214_ net627 _03844_ _03852_ vssd1 vssd1 vccd1 vccd1 _03853_ sky130_fd_sc_hd__and3_1
XFILLER_21_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09194_ top.CPU.registers.data\[550\] top.CPU.registers.data\[518\] net978 vssd1
+ vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__mux2_1
XANTENNA__11878__S net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08145_ _03783_ _03756_ net454 vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__mux2_1
X_14814__984 clknet_leaf_155_clk vssd1 vssd1 vccd1 vccd1 net2453 sky130_fd_sc_hd__inv_2
XANTENNA_fanout400_A net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07788__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08985__C1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload150 clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 clkload150/Y sky130_fd_sc_hd__inv_6
X_08076_ _03711_ _03714_ net618 _03706_ vssd1 vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__a211oi_1
XFILLER_101_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload161 clknet_leaf_114_clk vssd1 vssd1 vccd1 vccd1 clkload161/Y sky130_fd_sc_hd__inv_8
XFILLER_162_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload172 clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 clkload172/Y sky130_fd_sc_hd__inv_8
XFILLER_106_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload183 clknet_leaf_84_clk vssd1 vssd1 vccd1 vccd1 clkload183/Y sky130_fd_sc_hd__clkinv_4
XFILLER_122_608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload194 clknet_leaf_95_clk vssd1 vssd1 vccd1 vccd1 clkload194/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_8_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13665__Y _03047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout488_X net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout867_A net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold12 top.CPU.registers.data_out_r2_prev\[11\] vssd1 vssd1 vccd1 vccd1 net2569 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold23 top.CPU.registers.data_out_r1_prev\[9\] vssd1 vssd1 vccd1 vccd1 net2580 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08752__A2 _04390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10811__A net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08978_ net737 _04612_ _04613_ _04616_ net635 vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__a311o_1
XFILLER_60_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold34 top.CPU.registers.data_out_r2_prev\[20\] vssd1 vssd1 vccd1 vccd1 net2591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 top.I2C.I2C_state\[17\] vssd1 vssd1 vccd1 vccd1 net2602 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold56 top.I2C.I2C_state\[14\] vssd1 vssd1 vccd1 vccd1 net2613 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07960__B1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold67 top.I2C.I2C_state\[16\] vssd1 vssd1 vccd1 vccd1 net2624 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold78 top.CPU.registers.data_out_r1_prev\[29\] vssd1 vssd1 vccd1 vccd1 net2635 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11639__A2 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07929_ top.CPU.registers.data\[316\] net1026 net948 vssd1 vssd1 vccd1 vccd1 _03568_
+ sky130_fd_sc_hd__a21o_1
XFILLER_152_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout655_X net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold89 top.CPU.registers.data\[569\] vssd1 vssd1 vccd1 vccd1 net2646 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1397_X net1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09162__C1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08504__A2 net1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10847__B1 _05754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10940_ _03167_ _06447_ vssd1 vssd1 vccd1 vccd1 _06517_ sky130_fd_sc_hd__or2_1
XFILLER_17_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07712__B1 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout822_X net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10871_ net484 net460 _06475_ net220 net2983 vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__a32o_1
XFILLER_72_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12610_ _07106_ _07107_ _07108_ _07109_ vssd1 vssd1 vccd1 vccd1 _07110_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_27_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13590_ net1352 _06124_ vssd1 vssd1 vccd1 vccd1 _03020_ sky130_fd_sc_hd__nand2_1
XANTENNA__12064__A2 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13261__B2 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10075__A1 _04634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09112__A net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12541_ _03309_ net547 _03322_ _05609_ _07049_ vssd1 vssd1 vccd1 vccd1 _07050_ sky130_fd_sc_hd__a41o_1
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11272__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15260_ net1594 _01470_ net1235 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[60\]
+ sky130_fd_sc_hd__dfrtp_1
X_12472_ _03955_ _03984_ vssd1 vssd1 vccd1 vccd1 _06981_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_117_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11423_ _06563_ net277 net268 net3295 vssd1 vssd1 vccd1 vccd1 _02088_ sky130_fd_sc_hd__a22o_1
X_15191_ net1528 _01401_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r1_prev\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12473__A _04019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07779__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12772__B1 top.CPU.alu.program_counter\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08976__C1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11575__B2 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14059__229 clknet_leaf_134_clk vssd1 vssd1 vccd1 vccd1 net1698 sky130_fd_sc_hd__inv_2
X_11354_ net3713 net285 net275 _06314_ vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__a22o_1
X_10305_ net394 _05814_ vssd1 vssd1 vccd1 vccd1 _05937_ sky130_fd_sc_hd__or2_1
XANTENNA__08991__A2 net1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12119__A3 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11285_ net562 _06603_ _03183_ vssd1 vssd1 vccd1 vccd1 _06700_ sky130_fd_sc_hd__or3b_1
XFILLER_3_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08728__C1 net1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11327__B2 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10236_ _05631_ _05636_ net387 vssd1 vssd1 vccd1 vccd1 _05871_ sky130_fd_sc_hd__mux2_1
X_13024_ net2801 _07437_ net894 vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__mux2_1
XFILLER_112_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1010 net1012 vssd1 vssd1 vccd1 vccd1 net1010 sky130_fd_sc_hd__clkbuf_4
Xfanout1021 net1022 vssd1 vssd1 vccd1 vccd1 net1021 sky130_fd_sc_hd__buf_2
XFILLER_6_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10167_ _05512_ _05522_ _05611_ net445 vssd1 vssd1 vccd1 vccd1 _05804_ sky130_fd_sc_hd__a31o_1
Xfanout1032 _03333_ vssd1 vssd1 vccd1 vccd1 net1032 sky130_fd_sc_hd__clkbuf_4
Xfanout1043 _03165_ vssd1 vssd1 vccd1 vccd1 net1043 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10721__A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1054 _06891_ vssd1 vssd1 vccd1 vccd1 net1054 sky130_fd_sc_hd__buf_2
XFILLER_0_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1065 net1067 vssd1 vssd1 vccd1 vccd1 net1065 sky130_fd_sc_hd__clkbuf_4
XFILLER_66_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07951__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1076 net1079 vssd1 vssd1 vccd1 vccd1 net1076 sky130_fd_sc_hd__clkbuf_4
X_10098_ _03315_ _03444_ _05735_ vssd1 vssd1 vccd1 vccd1 _05736_ sky130_fd_sc_hd__a21oi_1
X_14975_ clknet_leaf_96_clk _01220_ net1258 vssd1 vssd1 vccd1 vccd1 top.SPI.paroutput\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1087 net1089 vssd1 vssd1 vccd1 vccd1 net1087 sky130_fd_sc_hd__clkbuf_4
Xfanout1098 net1100 vssd1 vssd1 vccd1 vccd1 net1098 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11255__C net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08900__C1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14460__630 clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 net2099 sky130_fd_sc_hd__inv_2
XFILLER_74_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10853__A3 _06139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14757__927 clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 net2396 sky130_fd_sc_hd__inv_2
XFILLER_34_157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12808_ _07260_ _07261_ vssd1 vssd1 vccd1 vccd1 _07262_ sky130_fd_sc_hd__nor2_1
XFILLER_50_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16546__RESET_B net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13788_ net17 net1050 net885 net2853 vssd1 vssd1 vccd1 vccd1 _02669_ sky130_fd_sc_hd__o22a_1
XANTENNA__13252__B2 _02803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09022__A net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15527_ net1861 _01737_ net1191 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[327\]
+ sky130_fd_sc_hd__dfrtp_1
X_12739_ _07196_ _07198_ vssd1 vssd1 vccd1 vccd1 _07199_ sky130_fd_sc_hd__xor2_1
X_14501__671 clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 net2140 sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15458_ net1792 _01668_ net1172 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[258\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09208__B1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13555__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10455__X _06082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15389_ net1723 _01599_ net1119 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[189\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08967__C1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold504 top.CPU.registers.data\[470\] vssd1 vssd1 vccd1 vccd1 net3061 sky130_fd_sc_hd__dlygate4sd3_1
Xhold515 top.CPU.registers.data\[356\] vssd1 vssd1 vccd1 vccd1 net3072 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08431__A1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10615__B net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold526 top.CPU.registers.data\[780\] vssd1 vssd1 vccd1 vccd1 net3083 sky130_fd_sc_hd__dlygate4sd3_1
Xhold537 top.CPU.registers.data\[887\] vssd1 vssd1 vccd1 vccd1 net3094 sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 top.CPU.registers.data\[483\] vssd1 vssd1 vccd1 vccd1 net3105 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09950_ _05579_ _05588_ _05582_ _03789_ vssd1 vssd1 vccd1 vccd1 _05589_ sky130_fd_sc_hd__a2bb2o_1
Xhold559 top.CPU.registers.data\[707\] vssd1 vssd1 vccd1 vccd1 net3116 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11318__B2 _06311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08719__C1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09692__A _05330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08901_ top.CPU.registers.data\[682\] top.CPU.registers.data\[650\] net809 vssd1
+ vssd1 vccd1 vccd1 _04540_ sky130_fd_sc_hd__mux2_1
XFILLER_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_9_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09881_ _03310_ _03313_ net547 vssd1 vssd1 vccd1 vccd1 _05520_ sky130_fd_sc_hd__and3_1
XANTENNA__08800__S net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15428__RESET_B net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08832_ top.CPU.registers.data\[555\] top.CPU.registers.data\[523\] net966 vssd1
+ vssd1 vccd1 vccd1 _04471_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1204 top.CPU.registers.data_out_r1_prev\[7\] vssd1 vssd1 vccd1 vccd1 net3761
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1215 top.CPU.data_out\[28\] vssd1 vssd1 vccd1 vccd1 net3772 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1226 top.CPU.registers.data\[747\] vssd1 vssd1 vccd1 vccd1 net3783 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16298__Q top.CPU.data_out\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11446__B _06033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1237 top.CPU.registers.data\[124\] vssd1 vssd1 vccd1 vccd1 net3794 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1248 top.CPU.handler.toreg\[12\] vssd1 vssd1 vccd1 vccd1 net3805 sky130_fd_sc_hd__dlygate4sd3_1
X_08763_ top.CPU.registers.data\[588\] net1316 net847 top.CPU.registers.data\[620\]
+ net767 vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout183_A _06777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1259 top.CPU.registers.data\[893\] vssd1 vssd1 vccd1 vccd1 net3816 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09144__C1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07714_ net1409 _03154_ net1278 net1282 _03104_ vssd1 vssd1 vccd1 vccd1 _03353_ sky130_fd_sc_hd__a2111o_2
XANTENNA__08498__A1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13491__A1 _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09695__B1 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08694_ top.CPU.registers.data\[813\] top.CPU.registers.data\[781\] net807 vssd1
+ vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__mux2_1
XANTENNA__07940__A _03544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13661__B _03152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07645_ _03277_ _03280_ _03282_ vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__a21o_2
XANTENNA_fanout350_A net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07576_ top.CPU.registers.data\[639\] net1337 net866 top.CPU.registers.data\[607\]
+ net802 vssd1 vssd1 vccd1 vccd1 _03215_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_24_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09998__A1 _04294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09315_ top.CPU.control_unit.instruction\[24\] _04595_ vssd1 vssd1 vccd1 vccd1 _04954_
+ sky130_fd_sc_hd__or2_1
XANTENNA__11181__B net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13794__A2 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout236_X net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout615_A net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1357_A top.SPI.state\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09246_ top.CPU.registers.data\[453\] net1310 net841 top.CPU.registers.data\[485\]
+ net713 vssd1 vssd1 vccd1 vccd1 _04885_ sky130_fd_sc_hd__a221o_1
XANTENNA__08670__A1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09177_ top.CPU.registers.data\[646\] net1317 net848 top.CPU.registers.data\[678\]
+ net722 vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_79_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1145_X net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08128_ net917 _03764_ _03766_ net620 vssd1 vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__o211a_1
XFILLER_147_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout984_A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08059_ net932 _03696_ _03697_ net952 vssd1 vssd1 vccd1 vccd1 _03698_ sky130_fd_sc_hd__o211a_1
XFILLER_134_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1312_X net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput46 net46 vssd1 vssd1 vccd1 vccd1 ADR_O[16] sky130_fd_sc_hd__buf_2
XANTENNA__11309__B2 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput57 net57 vssd1 vssd1 vccd1 vccd1 ADR_O[28] sky130_fd_sc_hd__buf_2
X_11070_ net3169 net366 _06590_ net323 vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__a22o_1
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 DAT_O[0] sky130_fd_sc_hd__buf_2
XANTENNA__08710__S net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 DAT_O[1] sky130_fd_sc_hd__buf_2
XANTENNA_fanout772_X net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10021_ net308 _05658_ _05659_ vssd1 vssd1 vccd1 vccd1 _05660_ sky130_fd_sc_hd__o21ai_1
XFILLER_103_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08725__A2 _04361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07933__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14444__614 clknet_leaf_195_clk vssd1 vssd1 vccd1 vccd1 net2083 sky130_fd_sc_hd__inv_2
XFILLER_91_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11972_ _06527_ net350 net183 net2812 vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__a22o_1
X_13711_ _03060_ _03061_ vssd1 vssd1 vccd1 vccd1 _02626_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_2_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11493__B1 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10923_ _06313_ _06468_ vssd1 vssd1 vccd1 vccd1 _06507_ sky130_fd_sc_hd__nor2_1
XFILLER_72_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16430_ clknet_leaf_56_clk _00012_ net1141 vssd1 vssd1 vccd1 vccd1 top.I2C.I2C_state\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13642_ net2889 _07242_ net665 vssd1 vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__mux2_1
X_10854_ _03314_ _06451_ _06461_ vssd1 vssd1 vccd1 vccd1 _06462_ sky130_fd_sc_hd__o21ai_2
XANTENNA__09438__B1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08157__S net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11091__B net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13785__A2 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16361_ clknet_leaf_31_clk _02570_ net1126 vssd1 vssd1 vccd1 vccd1 top.CPU.fetch.current_ra\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11245__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13573_ top.CPU.alu.program_counter\[10\] top.CPU.handler.state\[3\] vssd1 vssd1
+ vccd1 vccd1 _03010_ sky130_fd_sc_hd__or2_1
X_10785_ net381 _06394_ _06395_ net386 vssd1 vssd1 vccd1 vccd1 _06396_ sky130_fd_sc_hd__o211a_1
XFILLER_72_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15312_ net1646 _01522_ net1156 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[112\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_171_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12524_ _06998_ _07008_ vssd1 vssd1 vccd1 vccd1 _07033_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_171_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16292_ clknet_leaf_96_clk _02501_ net1247 vssd1 vssd1 vccd1 vccd1 top.CPU.data_out\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_13_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08681__A net1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12915__B _05429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14915__1085 clknet_leaf_171_clk vssd1 vssd1 vccd1 vccd1 net2554 sky130_fd_sc_hd__inv_2
X_15243_ net1577 _01453_ net1065 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[43\]
+ sky130_fd_sc_hd__dfrtp_1
X_12455_ _03475_ _03508_ _06963_ vssd1 vssd1 vccd1 vccd1 _06964_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_10_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11406_ _06536_ net280 net269 net3504 vssd1 vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__a22o_1
X_15174_ net1511 _01384_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r1_prev\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_12386_ top.CPU.addressnew\[25\] top.CPU.addressnew\[24\] top.CPU.addressnew\[27\]
+ top.CPU.addressnew\[26\] vssd1 vssd1 vccd1 vccd1 _06924_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10220__A1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11337_ net3687 net288 net282 _05935_ vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__a22o_1
XFILLER_153_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11268_ net3273 net293 _06691_ net481 vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14843__1013 clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 net2482 sky130_fd_sc_hd__inv_2
XFILLER_95_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13007_ top.SPI.paroutput\[2\] _07429_ _07431_ net2702 vssd1 vssd1 vccd1 vccd1 _01208_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08716__A2 net1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10219_ _05502_ net447 _05850_ _05436_ vssd1 vssd1 vccd1 vccd1 _05854_ sky130_fd_sc_hd__a31o_1
X_11199_ net660 _06270_ net429 vssd1 vssd1 vccd1 vccd1 _06657_ sky130_fd_sc_hd__and3_1
XANTENNA__07924__B1 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14958_ clknet_leaf_87_clk _01203_ net1264 vssd1 vssd1 vccd1 vccd1 top.SPI.busy sky130_fd_sc_hd__dfrtp_4
XFILLER_36_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11079__A3 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14187__357 clknet_leaf_134_clk vssd1 vssd1 vccd1 vccd1 net1826 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_50_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13473__A1 net1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09451__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09141__A2 net1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11484__B1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10597__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07601__B1_N net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10169__Y _05806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14228__398 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 net1867 sky130_fd_sc_hd__inv_2
XFILLER_50_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11787__A1 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09100_ top.CPU.registers.data\[231\] net1393 net832 top.CPU.registers.data\[199\]
+ net778 vssd1 vssd1 vccd1 vccd1 _04739_ sky130_fd_sc_hd__a221o_1
X_09031_ top.CPU.registers.data\[648\] net1314 net845 top.CPU.registers.data\[680\]
+ net716 vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__a221o_1
XFILLER_30_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07478__Y _03118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11539__B2 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold301 top.CPU.registers.data\[299\] vssd1 vssd1 vccd1 vccd1 net2858 sky130_fd_sc_hd__dlygate4sd3_1
Xhold312 top.CPU.registers.data\[923\] vssd1 vssd1 vccd1 vccd1 net2869 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold323 top.CPU.registers.data\[7\] vssd1 vssd1 vccd1 vccd1 net2880 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10211__A1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13496__X _02967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold334 top.CPU.registers.data\[596\] vssd1 vssd1 vccd1 vccd1 net2891 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09693__Y _05332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold345 top.CPU.registers.data\[15\] vssd1 vssd1 vccd1 vccd1 net2902 sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 top.CPU.addressnew\[27\] vssd1 vssd1 vccd1 vccd1 net2913 sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 top.CPU.registers.data\[95\] vssd1 vssd1 vccd1 vccd1 net2924 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold378 top.CPU.fetch.current_ra\[10\] vssd1 vssd1 vccd1 vccd1 net2935 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09933_ _04226_ _04257_ vssd1 vssd1 vccd1 vccd1 _05572_ sky130_fd_sc_hd__nor2_1
XANTENNA__07935__A net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold389 top.CPU.registers.data\[468\] vssd1 vssd1 vccd1 vccd1 net2946 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout803 net804 vssd1 vssd1 vccd1 vccd1 net803 sky130_fd_sc_hd__buf_2
XANTENNA__12560__B _05767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10632__Y _06251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout814 net822 vssd1 vssd1 vccd1 vccd1 net814 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08168__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout825 net831 vssd1 vssd1 vccd1 vccd1 net825 sky130_fd_sc_hd__buf_4
XANTENNA__09365__C1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11457__A net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout836 net839 vssd1 vssd1 vccd1 vccd1 net836 sky130_fd_sc_hd__clkbuf_4
X_09864_ _05501_ _05502_ vssd1 vssd1 vccd1 vccd1 _05503_ sky130_fd_sc_hd__nand2b_2
X_14131__301 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 net1770 sky130_fd_sc_hd__inv_2
Xfanout847 net848 vssd1 vssd1 vccd1 vccd1 net847 sky130_fd_sc_hd__clkbuf_4
Xfanout858 _03203_ vssd1 vssd1 vccd1 vccd1 net858 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1105_A net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07915__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1001 top.CPU.registers.data\[242\] vssd1 vssd1 vccd1 vccd1 net3558 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout869 net870 vssd1 vssd1 vccd1 vccd1 net869 sky130_fd_sc_hd__buf_2
Xhold1012 top.CPU.registers.data\[183\] vssd1 vssd1 vccd1 vccd1 net3569 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08815_ top.CPU.registers.data\[716\] net1372 net977 top.CPU.registers.data\[748\]
+ net930 vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__o221a_1
Xhold1023 top.CPU.registers.data\[961\] vssd1 vssd1 vccd1 vccd1 net3580 sky130_fd_sc_hd__dlygate4sd3_1
X_09795_ _05399_ _05430_ vssd1 vssd1 vccd1 vccd1 _05434_ sky130_fd_sc_hd__nand2_1
Xhold1034 top.CPU.registers.data\[475\] vssd1 vssd1 vccd1 vccd1 net3591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1045 top.CPU.registers.data\[739\] vssd1 vssd1 vccd1 vccd1 net3602 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout565_A net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout186_X net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11891__S net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1056 top.CPU.registers.data\[911\] vssd1 vssd1 vccd1 vccd1 net3613 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09117__C1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1067 net99 vssd1 vssd1 vccd1 vccd1 net3624 sky130_fd_sc_hd__dlygate4sd3_1
X_08746_ net1283 _04383_ _04384_ vssd1 vssd1 vccd1 vccd1 _04385_ sky130_fd_sc_hd__or3_1
XFILLER_26_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1078 top.CPU.registers.data\[663\] vssd1 vssd1 vccd1 vccd1 net3635 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1089 top.CPU.registers.data\[646\] vssd1 vssd1 vccd1 vccd1 net3646 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09361__S net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09132__A2 net1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11475__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout732_A net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout353_X net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08677_ top.CPU.registers.data\[654\] net1012 net934 _04315_ vssd1 vssd1 vccd1 vccd1
+ _04316_ sky130_fd_sc_hd__o211a_1
XANTENNA__08340__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07628_ top.CPU.control_unit.instruction\[30\] _03258_ _03266_ vssd1 vssd1 vccd1
+ vccd1 _03267_ sky130_fd_sc_hd__a21bo_1
XANTENNA__12019__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11227__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout520_X net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12575__X _07080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07559_ net1408 net1045 vssd1 vssd1 vccd1 vccd1 _03198_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_153_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout618_X net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10570_ net552 _06190_ vssd1 vssd1 vccd1 vccd1 _06192_ sky130_fd_sc_hd__or2_1
XFILLER_42_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12735__B _04598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09229_ net635 _04865_ _04867_ vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__o21a_1
XFILLER_155_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07851__C1 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12240_ net2844 _05771_ net433 vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__mux2_1
XFILLER_107_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout987_X net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12171_ net3731 net174 _06853_ vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__a21o_1
XFILLER_150_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Left_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11122_ net1405 net576 net528 net139 vssd1 vssd1 vccd1 vccd1 _06619_ sky130_fd_sc_hd__and4_1
XFILLER_122_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold890 top.CPU.registers.data\[658\] vssd1 vssd1 vccd1 vccd1 net3447 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13058__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09356__C1 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15930_ net2264 _02140_ net1253 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[730\]
+ sky130_fd_sc_hd__dfrtp_1
X_11053_ _06056_ net536 vssd1 vssd1 vccd1 vccd1 _06585_ sky130_fd_sc_hd__and2_1
XANTENNA__07906__B1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10004_ net413 _05616_ vssd1 vssd1 vccd1 vccd1 _05643_ sky130_fd_sc_hd__or2_4
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_129_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15861_ net2195 _02071_ net1216 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[661\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_88_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_129_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13455__A1 net1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15792_ net2126 _02002_ net1106 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[592\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11466__A0 _06354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11955_ _06502_ net341 net229 net3413 vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__a22o_1
XFILLER_33_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08331__B1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10906_ _06174_ _06466_ vssd1 vssd1 vccd1 vccd1 _06497_ sky130_fd_sc_hd__nor2_1
X_11886_ net142 net3028 net188 vssd1 vssd1 vccd1 vccd1 _01677_ sky130_fd_sc_hd__mux2_1
XFILLER_60_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16413_ clknet_leaf_56_clk _00037_ net1142 vssd1 vssd1 vccd1 vccd1 top.I2C.I2C_state\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13625_ top.CPU.alu.program_counter\[31\] _05688_ net1350 vssd1 vssd1 vccd1 vccd1
+ _03041_ sky130_fd_sc_hd__mux2_1
X_10837_ top.CPU.fetch.current_ra\[1\] net1041 net883 top.CPU.handler.toreg\[1\] vssd1
+ vssd1 vccd1 vccd1 _06446_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_15_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16344_ clknet_leaf_74_clk _02553_ net1159 vssd1 vssd1 vccd1 vccd1 top.CPU.addressnew\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_13556_ top.CPU.alu.program_counter\[3\] _06410_ net1348 vssd1 vssd1 vccd1 vccd1
+ _03000_ sky130_fd_sc_hd__mux2_1
XANTENNA__08095__C1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08634__A1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10768_ _06295_ _06379_ net386 vssd1 vssd1 vccd1 vccd1 _06380_ sky130_fd_sc_hd__mux2_1
XANTENNA__09831__B1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12645__B _06941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12507_ _06997_ _07015_ _06996_ vssd1 vssd1 vccd1 vccd1 _07016_ sky130_fd_sc_hd__o21ai_1
XFILLER_145_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16275_ clknet_leaf_33_clk _02485_ net1123 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.toreg\[19\]
+ sky130_fd_sc_hd__dfrtp_2
X_13487_ top.CPU.data_out\[1\] _05154_ net587 vssd1 vssd1 vccd1 vccd1 _02499_ sky130_fd_sc_hd__mux2_1
X_14572__742 clknet_leaf_195_clk vssd1 vssd1 vccd1 vccd1 net2211 sky130_fd_sc_hd__inv_2
X_10699_ net3880 net225 net315 _06314_ vssd1 vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__a22o_1
X_15226_ net1560 _01436_ net1254 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12438_ net1054 _06955_ vssd1 vssd1 vccd1 vccd1 _00054_ sky130_fd_sc_hd__and2_1
XFILLER_145_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10490__B1_N net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08398__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08937__A2 net1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15157_ clknet_leaf_40_clk _01367_ net1117 vssd1 vssd1 vccd1 vccd1 top.I2C.data_out\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_12369_ top.I2C.I2C_state\[24\] top.I2C.I2C_state\[22\] vssd1 vssd1 vccd1 vccd1 _06910_
+ sky130_fd_sc_hd__or2_1
XFILLER_153_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10733__X _06347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10744__A2 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14613__783 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 net2252 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_91_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15088_ net1470 _01301_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r2_prev\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_35_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11277__A net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09362__A2 net1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08570__B1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08600_ net963 _04235_ net624 vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__a21o_1
XFILLER_110_997 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09580_ net951 _05218_ vssd1 vssd1 vccd1 vccd1 _05219_ sky130_fd_sc_hd__or2_1
XANTENNA__12249__A2 _06010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07490__A net1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09114__A2 net1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08531_ top.CPU.registers.data\[176\] net1380 net983 top.CPU.registers.data\[144\]
+ net675 vssd1 vssd1 vccd1 vccd1 _04170_ sky130_fd_sc_hd__a221o_1
XFILLER_36_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08462_ top.CPU.registers.data\[465\] net1296 net1016 top.CPU.registers.data\[497\]
+ net913 vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__a221o_1
XANTENNA__11209__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08393_ top.CPU.registers.data\[946\] top.CPU.registers.data\[914\] top.CPU.registers.data\[818\]
+ top.CPU.registers.data\[786\] net982 net908 vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout146_A _06149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12421__A2 _06941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10356__A _05983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout313_A net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09014_ top.CPU.registers.data\[201\] net1369 net964 top.CPU.registers.data\[233\]
+ net926 vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__o221a_1
XANTENNA__10983__A2 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12185__A1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11886__S net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08928__A2 _04566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold120 top.CPU.registers.data\[297\] vssd1 vssd1 vccd1 vccd1 net2677 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12571__A _06462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold131 top.CPU.registers.data\[906\] vssd1 vssd1 vccd1 vccd1 net2688 sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 net48 vssd1 vssd1 vccd1 vccd1 net2699 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10196__B1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1222_A net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold153 top.CPU.fetch.current_ra\[30\] vssd1 vssd1 vccd1 vccd1 net2710 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_72_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold164 top.CPU.registers.data\[424\] vssd1 vssd1 vccd1 vccd1 net2721 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 top.CPU.registers.data\[560\] vssd1 vssd1 vccd1 vccd1 net2732 sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 top.CPU.registers.data\[407\] vssd1 vssd1 vccd1 vccd1 net2743 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout682_A net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout600 _05690_ vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__buf_4
Xhold197 top.CPU.registers.data\[411\] vssd1 vssd1 vccd1 vccd1 net2754 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout611 net616 vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__clkbuf_8
XFILLER_120_728 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09916_ _04990_ _05544_ _05554_ vssd1 vssd1 vccd1 vccd1 _05555_ sky130_fd_sc_hd__or3b_1
Xfanout622 net623 vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__clkbuf_4
Xfanout633 net634 vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1010_X net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout644 _03202_ vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__buf_4
XFILLER_113_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1108_X net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout655 net657 vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_146_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout666 _03042_ vssd1 vssd1 vccd1 vccd1 net666 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_146_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout677 net684 vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11696__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09847_ top.CPU.registers.data\[922\] net1305 net1027 top.CPU.registers.data\[954\]
+ net921 vssd1 vssd1 vccd1 vccd1 _05486_ sky130_fd_sc_hd__a221o_1
Xfanout688 _03332_ vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__buf_4
XANTENNA_fanout470_X net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout699 net701 vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__buf_4
XANTENNA_fanout947_A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout568_X net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11160__A2 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13606__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14914__1084 clknet_leaf_143_clk vssd1 vssd1 vccd1 vccd1 net2553 sky130_fd_sc_hd__inv_2
X_09778_ net915 _05416_ vssd1 vssd1 vccd1 vccd1 _05417_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_107_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11448__A0 _06056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08729_ top.CPU.registers.data\[333\] net1371 net967 top.CPU.registers.data\[365\]
+ net1280 vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout735_X net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09510__C1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _06585_ net499 net193 net3178 vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__a22o_1
XANTENNA__10120__B1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout902_X net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11671_ net464 _06486_ net238 net166 net2979 vssd1 vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_120_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10818__X _06428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_970 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13410_ top.mmio.mem_data_i\[28\] net593 net67 vssd1 vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_12_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10622_ _04430_ _04532_ net376 vssd1 vssd1 vccd1 vccd1 _06241_ sky130_fd_sc_hd__mux2_1
X_14556__726 clknet_leaf_140_clk vssd1 vssd1 vccd1 vccd1 net2195 sky130_fd_sc_hd__inv_2
X_14842__1012 clknet_leaf_164_clk vssd1 vssd1 vccd1 vccd1 net2481 sky130_fd_sc_hd__inv_2
XFILLER_169_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13341_ net888 _02874_ vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__and2_1
XANTENNA__11620__B1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_839 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10553_ net3806 net226 net315 _06175_ vssd1 vssd1 vccd1 vccd1 _02417_ sky130_fd_sc_hd__a22o_1
XFILLER_155_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10974__A2 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14300__470 clknet_leaf_139_clk vssd1 vssd1 vccd1 vccd1 net1939 sky130_fd_sc_hd__inv_2
X_16060_ net2394 _02270_ net1193 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[860\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_143_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13272_ top.I2C.data_out\[0\] net891 _06948_ vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__mux2_1
X_10484_ _05293_ _06108_ vssd1 vssd1 vccd1 vccd1 _06109_ sky130_fd_sc_hd__xnor2_1
XFILLER_170_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15011_ clknet_leaf_96_clk _01256_ net1253 vssd1 vssd1 vccd1 vccd1 top.SPI.parameters\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09577__C1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12223_ top.CPU.registers.data\[39\] net657 _03185_ vssd1 vssd1 vccd1 vccd1 _06878_
+ sky130_fd_sc_hd__o21a_1
XFILLER_170_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09592__A2 _03152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12154_ top.CPU.registers.data\[75\] net645 net244 vssd1 vssd1 vccd1 vccd1 _06845_
+ sky130_fd_sc_hd__o21a_1
X_13924__94 clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 net1563 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_166_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09329__C1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11105_ net494 net469 _06610_ net304 net3066 vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__a32o_1
XFILLER_151_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12085_ net564 net360 _06622_ net176 top.CPU.registers.data\[110\] vssd1 vssd1 vccd1
+ vccd1 _06811_ sky130_fd_sc_hd__a32o_1
XFILLER_96_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11036_ net3303 net368 _06577_ net321 vssd1 vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__a22o_1
X_15913_ net2247 _02123_ net1055 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[713\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11687__B1 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08001__C1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15844_ net2178 _02054_ net1198 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[644\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13428__A1 _02855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15775_ net2109 _01985_ net1223 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[575\]
+ sky130_fd_sc_hd__dfrtp_1
X_12987_ net3715 _07415_ _07417_ vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__o21a_1
XFILLER_73_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12100__A1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09501__C1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09789__X _05428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11938_ _06476_ net353 net232 net3236 vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__a22o_1
XFILLER_60_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12656__A top.CPU.alu.program_counter\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11869_ net135 net3225 net190 vssd1 vssd1 vccd1 vccd1 _01693_ sky130_fd_sc_hd__mux2_1
XFILLER_32_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12939__B1 top.CPU.alu.program_counter\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13251__S _02780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13608_ top.CPU.alu.program_counter\[23\] net1348 net583 vssd1 vssd1 vccd1 vccd1
+ _03032_ sky130_fd_sc_hd__o21a_1
XFILLER_159_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14299__469 clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 net1938 sky130_fd_sc_hd__inv_2
XANTENNA__09804__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xteam_08_1422 vssd1 vssd1 vccd1 vccd1 team_08_1422/HI gpio_oeb[8] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_31_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16327_ clknet_leaf_80_clk _02536_ net1241 vssd1 vssd1 vccd1 vccd1 top.CPU.addressnew\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xteam_08_1433 vssd1 vssd1 vccd1 vccd1 team_08_1433/HI gpio_out[18] sky130_fd_sc_hd__conb_1
XANTENNA__11611__A0 _06149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_08_1444 vssd1 vssd1 vccd1 vccd1 team_08_1444/HI gpio_out[29] sky130_fd_sc_hd__conb_1
X_13539_ _03575_ net585 vssd1 vssd1 vccd1 vccd1 _02990_ sky130_fd_sc_hd__and2_1
Xteam_08_1455 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] team_08_1455/LO sky130_fd_sc_hd__conb_1
XANTENNA__09280__A1 top.CPU.control_unit.instruction\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_71_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xteam_08_1466 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] team_08_1466/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_93_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16258_ clknet_leaf_29_clk _02468_ net1153 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.toreg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_145_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15209_ net1543 _01419_ net1061 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09568__C1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12391__A top.CPU.addressnew\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16189_ net2523 _02399_ net1114 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[989\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_141_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11390__A2 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07962_ top.CPU.registers.data\[824\] net1390 net820 top.CPU.registers.data\[792\]
+ net694 vssd1 vssd1 vccd1 vccd1 _03601_ sky130_fd_sc_hd__a221o_1
XFILLER_101_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09701_ top.CPU.registers.data\[345\] net1306 net1029 top.CPU.registers.data\[377\]
+ net946 vssd1 vssd1 vccd1 vccd1 _05340_ sky130_fd_sc_hd__a221o_1
XANTENNA__09335__A2 net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11678__B1 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10910__Y _06500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07893_ top.CPU.registers.data\[316\] top.CPU.registers.data\[284\] net833 vssd1
+ vssd1 vccd1 vccd1 _03532_ sky130_fd_sc_hd__mux2_1
XANTENNA__11142__A2 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13426__S net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09632_ _05127_ _05269_ _05058_ _05124_ vssd1 vssd1 vccd1 vccd1 _05271_ sky130_fd_sc_hd__o211ai_2
XANTENNA__09740__C1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_74_Left_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12330__S net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12890__A2 _03118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10996__D net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09563_ top.CPU.registers.data\[832\] net1293 net1005 top.CPU.registers.data\[864\]
+ net928 vssd1 vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_69_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout263_A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08514_ net793 _04141_ _04142_ _04152_ net706 vssd1 vssd1 vccd1 vccd1 _04153_ sky130_fd_sc_hd__a311o_1
XANTENNA_clkbuf_leaf_162_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14243__413 clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 net1882 sky130_fd_sc_hd__inv_2
X_09494_ net628 _05132_ _05131_ net608 vssd1 vssd1 vccd1 vccd1 _05133_ sky130_fd_sc_hd__a211o_1
XFILLER_23_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08445_ net754 _04082_ _04083_ net700 vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_102_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout430_A _06642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11850__B1 net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_42_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12566__A _06309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1172_A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout528_A net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08059__C1 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08376_ net744 _04006_ _04007_ net706 vssd1 vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__a31o_1
XFILLER_143_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10357__Y _05988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12285__B _06887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_177_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_83_Left_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11602__B1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09271__A1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout316_X net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_57_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09559__C1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_100_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_148_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_148_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11629__B net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08231__C1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout685_X net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11381__A2 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1406 net1407 vssd1 vssd1 vccd1 vccd1 net1406 sky130_fd_sc_hd__buf_4
XANTENNA__13658__A1 _07391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout430 _06642_ vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__clkbuf_4
XFILLER_24_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout441 net442 vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__clkbuf_4
Xfanout452 net453 vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__clkbuf_4
Xfanout463 _03194_ vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_115_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11669__B1 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_92_Left_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout852_X net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout474 _03193_ vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__buf_4
Xfanout485 net486 vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_161_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12910_ _07347_ _07353_ net129 vssd1 vssd1 vccd1 vccd1 _07354_ sky130_fd_sc_hd__mux2_1
XFILLER_111_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09731__C1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout496 net497 vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12240__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07888__A2 net1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11684__A3 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12841_ top.CPU.alu.program_counter\[20\] _03685_ vssd1 vssd1 vccd1 vccd1 _07291_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__11364__B net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07561__C net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10892__B2 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15560_ net1894 _01770_ net1098 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[360\]
+ sky130_fd_sc_hd__dfrtp_1
X_12772_ top.CPU.alu.program_counter\[12\] _07208_ top.CPU.alu.program_counter\[13\]
+ vssd1 vssd1 vccd1 vccd1 _07229_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11083__C _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11723_ _06566_ net203 net422 net3317 vssd1 vssd1 vccd1 vccd1 _01830_ sky130_fd_sc_hd__a22o_1
X_15491_ net1825 _01701_ net1209 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[291\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11841__B1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11654_ _06336_ net206 net427 net3339 vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__a22o_1
XFILLER_70_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13594__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10605_ net548 _04469_ net503 _04465_ _06224_ vssd1 vssd1 vccd1 vccd1 _06225_ sky130_fd_sc_hd__o221a_1
X_14027__197 clknet_leaf_134_clk vssd1 vssd1 vccd1 vccd1 net1666 sky130_fd_sc_hd__inv_2
XANTENNA__09798__C1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08065__A2 net1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11585_ _06696_ net260 net248 net2704 vssd1 vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__a22o_1
XFILLER_127_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10947__A2 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16112_ net2446 _02322_ net1154 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[912\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_167_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13324_ net1343 top.mmio.mem_data_i\[5\] net596 vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__o21a_1
XFILLER_6_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10536_ net371 _06155_ _06158_ net511 vssd1 vssd1 vccd1 vccd1 _06159_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_116_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07812__A2 net1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13346__A0 net1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire897 _07422_ vssd1 vssd1 vccd1 vccd1 net897 sky130_fd_sc_hd__buf_2
XFILLER_143_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12149__B2 _06500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16043_ net2377 _02253_ net1058 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[843\]
+ sky130_fd_sc_hd__dfrtp_1
X_13255_ top.I2C.data_out\[8\] net893 _06948_ vssd1 vssd1 vccd1 vccd1 _02812_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_108_Right_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10467_ _04052_ _05680_ vssd1 vssd1 vccd1 vccd1 _06093_ sky130_fd_sc_hd__nand2_1
XFILLER_124_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12206_ net3828 net652 _06870_ vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__o21a_1
X_13186_ _03124_ _02758_ _02765_ _02766_ vssd1 vssd1 vccd1 vccd1 _02767_ sky130_fd_sc_hd__a31o_1
XFILLER_89_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10398_ _06026_ vssd1 vssd1 vccd1 vccd1 _06027_ sky130_fd_sc_hd__inv_2
XFILLER_9_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11372__A2 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12137_ net3902 net649 _06836_ vssd1 vssd1 vccd1 vccd1 _01494_ sky130_fd_sc_hd__o21a_1
X_14684__854 clknet_leaf_138_clk vssd1 vssd1 vccd1 vccd1 net2323 sky130_fd_sc_hd__inv_2
XANTENNA__09724__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12068_ top.CPU.registers.data\[119\] net178 vssd1 vssd1 vccd1 vccd1 _06803_ sky130_fd_sc_hd__and2_1
XFILLER_38_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12321__A1 _03984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11019_ net3223 net218 _06566_ net322 vssd1 vssd1 vccd1 vccd1 _02342_ sky130_fd_sc_hd__a22o_1
XANTENNA__10332__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11675__A3 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14725__895 clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 net2364 sky130_fd_sc_hd__inv_2
XANTENNA__09025__A _04634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15827_ net2161 _02037_ net1177 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[627\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_92_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12085__B1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15758_ net2092 _01968_ net1193 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[558\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11832__B1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15689_ net2023 _01899_ net1056 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[489\]
+ sky130_fd_sc_hd__dfrtp_1
X_08230_ net802 _03864_ _03865_ net756 vssd1 vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__o211a_1
XFILLER_165_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08161_ net707 _03798_ _03799_ vssd1 vssd1 vccd1 vccd1 _03800_ sky130_fd_sc_hd__or3_1
XFILLER_147_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08092_ net643 _03727_ _03730_ vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__or3_1
XANTENNA__08461__C1 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14913__1083 clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 net2552 sky130_fd_sc_hd__inv_2
XANTENNA__12833__B _03986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload40 clknet_leaf_181_clk vssd1 vssd1 vccd1 vccd1 clkload40/Y sky130_fd_sc_hd__inv_16
XANTENNA__07486__Y _03126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10056__D net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload51 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 clkload51/Y sky130_fd_sc_hd__inv_4
Xclkload62 clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 clkload62/Y sky130_fd_sc_hd__clkinv_8
Xclkload73 clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 clkload73/Y sky130_fd_sc_hd__clkinv_4
XFILLER_161_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload84 clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 clkload84/Y sky130_fd_sc_hd__clkinv_4
Xclkload95 clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 clkload95/Y sky130_fd_sc_hd__inv_16
XFILLER_115_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11449__B net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11899__B1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_1035 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08994_ _04618_ _04632_ vssd1 vssd1 vccd1 vccd1 _04633_ sky130_fd_sc_hd__or2_4
XFILLER_125_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1018_A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07945_ top.CPU.registers.data\[56\] top.CPU.registers.data\[24\] net820 vssd1 vssd1
+ vccd1 vccd1 _03584_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_143_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14841__1011 clknet_leaf_177_clk vssd1 vssd1 vccd1 vccd1 net2480 sky130_fd_sc_hd__inv_2
XANTENNA__11115__A2 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12312__A1 _03575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout478_A net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09713__C1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07876_ net755 _03513_ _03514_ net712 vssd1 vssd1 vccd1 vccd1 _03515_ sky130_fd_sc_hd__o211a_1
XANTENNA__11666__A3 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09615_ top.CPU.registers.data\[960\] net1315 net846 top.CPU.registers.data\[992\]
+ net715 vssd1 vssd1 vccd1 vccd1 _05254_ sky130_fd_sc_hd__a221o_1
XANTENNA__11184__B net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout645_A net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout266_X net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1387_A net1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12076__B1 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09546_ top.CPU.registers.data\[289\] top.CPU.registers.data\[257\] net835 vssd1
+ vssd1 vccd1 vccd1 _05185_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_84_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08819__A1 _03116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15805__RESET_B net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11823__B1 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09477_ top.CPU.registers.data\[898\] net1324 net855 top.CPU.registers.data\[930\]
+ net723 vssd1 vssd1 vccd1 vccd1 _05116_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout812_A net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11300__A1_N _05960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout433_X net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09492__A1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08428_ top.CPU.registers.data\[433\] top.CPU.registers.data\[401\] net825 vssd1
+ vssd1 vccd1 vccd1 _04067_ sky130_fd_sc_hd__mux2_1
XFILLER_157_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload1 clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clkload1/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA_fanout600_X net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08359_ top.CPU.registers.data\[754\] net1389 net815 top.CPU.registers.data\[722\]
+ net718 vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_22_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10929__A2 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11370_ net495 net476 _06481_ net274 net3405 vssd1 vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__a32o_1
XANTENNA__08713__S net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10321_ _05643_ _05949_ _05950_ _05687_ _05945_ vssd1 vssd1 vccd1 vccd1 _05953_ sky130_fd_sc_hd__o32a_1
XFILLER_137_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14371__541 clknet_leaf_171_clk vssd1 vssd1 vccd1 vccd1 net2010 sky130_fd_sc_hd__inv_2
X_13040_ net2892 _07445_ net896 vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_115_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09547__A2 net1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10252_ _05825_ _05885_ net309 vssd1 vssd1 vccd1 vccd1 _05886_ sky130_fd_sc_hd__mux2_1
XANTENNA__12000__B1 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08204__C1 net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14668__838 clknet_leaf_195_clk vssd1 vssd1 vccd1 vccd1 net2307 sky130_fd_sc_hd__inv_2
XFILLER_3_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07558__A1 net1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11354__A2 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10183_ net382 _05716_ _05818_ vssd1 vssd1 vccd1 vccd1 _05819_ sky130_fd_sc_hd__o21ai_1
XFILLER_78_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1203 net1204 vssd1 vssd1 vccd1 vccd1 net1203 sky130_fd_sc_hd__clkbuf_4
Xfanout1214 net1218 vssd1 vssd1 vccd1 vccd1 net1214 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09544__S net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1225 net1226 vssd1 vssd1 vccd1 vccd1 net1225 sky130_fd_sc_hd__buf_2
Xfanout1236 net1276 vssd1 vssd1 vccd1 vccd1 net1236 sky130_fd_sc_hd__buf_2
X_14412__582 clknet_leaf_195_clk vssd1 vssd1 vccd1 vccd1 net2051 sky130_fd_sc_hd__inv_2
XFILLER_78_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14991_ clknet_leaf_93_clk _01236_ net1268 vssd1 vssd1 vccd1 vccd1 top.SPI.paroutput\[30\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1247 net1249 vssd1 vssd1 vccd1 vccd1 net1247 sky130_fd_sc_hd__clkbuf_4
Xfanout1258 net1259 vssd1 vssd1 vccd1 vccd1 net1258 sky130_fd_sc_hd__clkbuf_2
Xfanout260 net261 vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__buf_4
Xfanout1269 net1270 vssd1 vssd1 vccd1 vccd1 net1269 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12303__A1 _04889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout271 _06714_ vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__clkbuf_8
X_14709__879 clknet_leaf_172_clk vssd1 vssd1 vccd1 vccd1 net2348 sky130_fd_sc_hd__inv_2
XANTENNA__08507__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout282 net283 vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__buf_4
XFILLER_87_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout293 _06662_ vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12854__A2 _03685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09180__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11094__B net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15612_ net1946 _01822_ net1234 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[412\]
+ sky130_fd_sc_hd__dfrtp_1
X_12824_ top.CPU.alu.program_counter\[18\] _04050_ vssd1 vssd1 vccd1 vccd1 _07276_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__12067__B1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15546__RESET_B net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15543_ net1877 _01753_ net1181 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[343\]
+ sky130_fd_sc_hd__dfrtp_1
X_12755_ top.CPU.alu.program_counter\[12\] _04462_ vssd1 vssd1 vccd1 vccd1 _07213_
+ sky130_fd_sc_hd__and2_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10719__A _06333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11706_ _06538_ net203 net422 net3123 vssd1 vssd1 vccd1 vccd1 _01847_ sky130_fd_sc_hd__a22o_1
X_15474_ net1808 _01684_ net1102 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[274\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_139_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ _07149_ _07150_ vssd1 vssd1 vccd1 vccd1 _07151_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_139_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08038__A2 net1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11637_ _05963_ net202 net424 net3330 vssd1 vssd1 vccd1 vccd1 _01914_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_42_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12934__A top.CPU.alu.program_counter\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11568_ net571 _06679_ vssd1 vssd1 vccd1 vccd1 _06743_ sky130_fd_sc_hd__nor2_1
Xhold708 top.I2C.data_out\[28\] vssd1 vssd1 vccd1 vccd1 net3265 sky130_fd_sc_hd__dlygate4sd3_1
X_13307_ top.CPU.control_unit.instruction\[0\] _02849_ net669 vssd1 vssd1 vccd1 vccd1
+ _02434_ sky130_fd_sc_hd__mux2_1
XFILLER_116_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14922__Q top.CPU.alu.program_counter\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10519_ _04192_ net505 vssd1 vssd1 vccd1 vccd1 _06143_ sky130_fd_sc_hd__nor2_1
XFILLER_7_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold719 top.CPU.registers.data\[358\] vssd1 vssd1 vccd1 vccd1 net3276 sky130_fd_sc_hd__dlygate4sd3_1
X_11499_ _06632_ net261 net256 net3107 vssd1 vssd1 vccd1 vccd1 _02025_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_139_Left_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmax_cap449 _04696_ vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__clkbuf_4
X_16026_ net2360 _02236_ net1250 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[826\]
+ sky130_fd_sc_hd__dfrtp_1
X_13238_ net3790 _02779_ _02802_ _02773_ vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__a22o_1
XANTENNA__10173__B net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12542__A1 _03252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11345__A2 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13169_ _06947_ _02752_ _02751_ vssd1 vssd1 vccd1 vccd1 _02754_ sky130_fd_sc_hd__a21o_1
XANTENNA__08210__A2 net1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10553__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09454__S net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1408 top.CPU.registers.data\[91\] vssd1 vssd1 vccd1 vccd1 net3965 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1419 top.CPU.addressnew\[4\] vssd1 vssd1 vccd1 vccd1 net3976 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10901__B net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11285__A net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07730_ _03098_ net688 net608 _03361_ _03368_ vssd1 vssd1 vccd1 vccd1 _03369_ sky130_fd_sc_hd__o221a_4
XANTENNA__12845__A2 _03986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10856__A1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07661_ _03161_ _03272_ vssd1 vssd1 vccd1 vccd1 _03300_ sky130_fd_sc_hd__nand2b_1
XFILLER_77_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07721__A1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_148_Left_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09400_ _05035_ _05038_ net637 vssd1 vssd1 vccd1 vccd1 _05039_ sky130_fd_sc_hd__a21o_1
XANTENNA__12058__B1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07592_ net779 _03229_ _03230_ net711 vssd1 vssd1 vccd1 vccd1 _03231_ sky130_fd_sc_hd__o31a_1
XFILLER_18_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10608__A1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09331_ top.CPU.registers.data\[900\] net1329 net860 top.CPU.registers.data\[932\]
+ net726 vssd1 vssd1 vccd1 vccd1 _04970_ sky130_fd_sc_hd__a221o_1
XANTENNA__10188__X _05824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_5_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09262_ top.CPU.registers.data\[69\] net1286 net1004 top.CPU.registers.data\[101\]
+ net950 vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__a221o_1
XANTENNA__08682__C1 top.CPU.control_unit.instruction\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11820__A3 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08213_ net954 _03846_ _03848_ _03851_ vssd1 vssd1 vccd1 vccd1 _03852_ sky130_fd_sc_hd__a31o_1
XANTENNA__09226__A1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09193_ top.CPU.registers.data\[934\] top.CPU.registers.data\[902\] top.CPU.registers.data\[806\]
+ top.CPU.registers.data\[774\] net978 net904 vssd1 vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__mux4_1
XANTENNA__08029__A2 net1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout226_A net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08144_ net680 _03776_ _03782_ _03770_ vssd1 vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__a31o_4
XFILLER_162_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12563__B _06081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14355__525 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 net1994 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_157_Left_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11584__A2 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload140 clknet_leaf_148_clk vssd1 vssd1 vccd1 vccd1 clkload140/Y sky130_fd_sc_hd__inv_12
X_08075_ net675 _03712_ _03713_ net604 vssd1 vssd1 vccd1 vccd1 _03714_ sky130_fd_sc_hd__a31oi_1
XFILLER_161_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload151 clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 clkload151/Y sky130_fd_sc_hd__inv_6
XANTENNA_fanout1135_A net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload162 clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 clkload162/Y sky130_fd_sc_hd__clkinv_16
Xclkload173 clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 clkload173/Y sky130_fd_sc_hd__clkinv_8
Xclkload184 clknet_leaf_85_clk vssd1 vssd1 vccd1 vccd1 clkload184/Y sky130_fd_sc_hd__clkinv_4
XFILLER_106_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload195 clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 clkload195/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_8_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12850__Y _07300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11336__A2 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11894__S net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08737__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08201__A2 net1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1302_A net1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09217__X _04856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold13 top.CPU.registers.data_out_r2_prev\[22\] vssd1 vssd1 vccd1 vccd1 net2570 sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ net783 _04614_ _04615_ net713 vssd1 vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__o211a_1
Xhold24 top.CPU.registers.data_out_r1_prev\[10\] vssd1 vssd1 vccd1 vccd1 net2581 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout383_X net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold35 top.CPU.registers.data_out_r2_prev\[30\] vssd1 vssd1 vccd1 vccd1 net2592 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout762_A net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold46 _00027_ vssd1 vssd1 vccd1 vccd1 net2603 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold57 _00038_ vssd1 vssd1 vccd1 vccd1 net2614 sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ top.CPU.registers.data\[412\] net996 _03566_ vssd1 vssd1 vccd1 vccd1 _03567_
+ sky130_fd_sc_hd__a21o_1
Xhold68 _00030_ vssd1 vssd1 vccd1 vccd1 net2625 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 net54 vssd1 vssd1 vccd1 vccd1 net2636 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_166_Left_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09701__A2 net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout550_X net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10847__B2 _05937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07859_ net674 _03493_ _03494_ _03497_ net610 vssd1 vssd1 vccd1 vccd1 _03498_ sky130_fd_sc_hd__a311o_1
XANTENNA_fanout1292_X net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout648_X net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12049__B1 _06780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10870_ net659 _05808_ net435 vssd1 vssd1 vccd1 vccd1 _06475_ sky130_fd_sc_hd__and3_1
XANTENNA__08708__S net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09529_ top.CPU.registers.data\[673\] top.CPU.registers.data\[641\] net838 vssd1
+ vssd1 vccd1 vccd1 _05168_ sky130_fd_sc_hd__mux2_1
XFILLER_25_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout815_X net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12540_ _03309_ _07041_ _07048_ _03252_ vssd1 vssd1 vccd1 vccd1 _07049_ sky130_fd_sc_hd__a22o_1
XANTENNA__11272__A1 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13963__133 clknet_leaf_149_clk vssd1 vssd1 vccd1 vccd1 net1602 sky130_fd_sc_hd__inv_2
XANTENNA__13549__A0 top.CPU.alu.program_counter\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08009__A _03613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11811__A3 net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12471_ _04019_ _04048_ vssd1 vssd1 vccd1 vccd1 _06980_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_173_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11422_ _06561_ net283 net270 net2739 vssd1 vssd1 vccd1 vccd1 _02089_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_117_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15190_ net1527 _01400_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r1_prev\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11024__B2 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12221__B1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08425__C1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08443__S net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12473__B _04048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12772__A1 top.CPU.alu.program_counter\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11575__A2 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08976__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14098__268 clknet_leaf_201_clk vssd1 vssd1 vccd1 vccd1 net1737 sky130_fd_sc_hd__inv_2
XFILLER_125_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11353_ net3711 net285 net275 _06293_ vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__a22o_1
XANTENNA__08440__A2 net1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10274__A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10304_ _03650_ _04060_ _05299_ vssd1 vssd1 vccd1 vccd1 _05936_ sky130_fd_sc_hd__nand3_1
XANTENNA__11089__B net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11284_ net312 net525 _06572_ net293 net2693 vssd1 vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__a32o_1
XFILLER_79_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11327__A2 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13023_ top.SPI.parameters\[13\] top.SPI.paroutput\[5\] net1355 vssd1 vssd1 vccd1
+ vccd1 _07437_ sky130_fd_sc_hd__mux2_1
X_10235_ _05869_ vssd1 vssd1 vccd1 vccd1 _05870_ sky130_fd_sc_hd__inv_2
Xfanout1000 net1001 vssd1 vssd1 vccd1 vccd1 net1000 sky130_fd_sc_hd__clkbuf_4
Xfanout1011 net1012 vssd1 vssd1 vccd1 vccd1 net1011 sky130_fd_sc_hd__clkbuf_2
Xfanout1022 net1032 vssd1 vssd1 vccd1 vccd1 net1022 sky130_fd_sc_hd__clkbuf_4
X_10166_ _05642_ _05802_ vssd1 vssd1 vccd1 vccd1 _05803_ sky130_fd_sc_hd__nand2_1
Xfanout1033 net1037 vssd1 vssd1 vccd1 vccd1 net1033 sky130_fd_sc_hd__buf_4
XFILLER_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1044 _03165_ vssd1 vssd1 vccd1 vccd1 net1044 sky130_fd_sc_hd__clkbuf_2
XFILLER_121_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1055 net1056 vssd1 vssd1 vccd1 vccd1 net1055 sky130_fd_sc_hd__clkbuf_4
Xfanout1066 net1067 vssd1 vssd1 vccd1 vccd1 net1066 sky130_fd_sc_hd__clkbuf_2
Xfanout1077 net1079 vssd1 vssd1 vccd1 vccd1 net1077 sky130_fd_sc_hd__clkbuf_4
X_10097_ _03443_ _05670_ net507 _03409_ _05734_ vssd1 vssd1 vccd1 vccd1 _05735_ sky130_fd_sc_hd__a221o_1
X_14974_ clknet_leaf_98_clk _01219_ net1254 vssd1 vssd1 vccd1 vccd1 top.SPI.paroutput\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1088 net1089 vssd1 vssd1 vccd1 vccd1 net1088 sky130_fd_sc_hd__clkbuf_4
Xfanout1099 net1100 vssd1 vssd1 vccd1 vccd1 net1099 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10838__A1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08685__Y _04324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14912__1082 clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 net2551 sky130_fd_sc_hd__inv_2
XANTENNA_clkload4_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08618__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14796__966 clknet_leaf_195_clk vssd1 vssd1 vccd1 vccd1 net2435 sky130_fd_sc_hd__inv_2
X_12807_ top.CPU.alu.program_counter\[15\] _07240_ top.CPU.alu.program_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 _07261_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13788__B1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13787_ net16 net1050 net885 net3859 vssd1 vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__o22a_1
XANTENNA__08259__A2 net1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10999_ net524 _06553_ vssd1 vssd1 vccd1 vccd1 _06554_ sky130_fd_sc_hd__nor2_1
XANTENNA__12055__A3 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12738_ _07185_ _07197_ vssd1 vssd1 vccd1 vccd1 _07198_ sky130_fd_sc_hd__or2_1
X_15526_ net1860 _01736_ net1073 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[326\]
+ sky130_fd_sc_hd__dfrtp_1
X_14042__212 clknet_leaf_150_clk vssd1 vssd1 vccd1 vccd1 net1681 sky130_fd_sc_hd__inv_2
XFILLER_124_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09208__A1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15457_ net1791 _01667_ net1231 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[257\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13841__11_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12669_ _07135_ _07134_ net125 vssd1 vssd1 vccd1 vccd1 _07136_ sky130_fd_sc_hd__mux2_1
X_14339__509 clknet_leaf_114_clk vssd1 vssd1 vccd1 vccd1 net1978 sky130_fd_sc_hd__inv_2
XANTENNA__12664__A top.CPU.alu.program_counter\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14840__1010 clknet_leaf_168_clk vssd1 vssd1 vccd1 vccd1 net2479 sky130_fd_sc_hd__inv_2
XANTENNA__12212__B1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_160_Right_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15388_ net1722 _01598_ net1236 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[188\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_144_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11566__A2 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold505 top.CPU.registers.data\[384\] vssd1 vssd1 vccd1 vccd1 net3062 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10774__B1 _05680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold516 top.CPU.registers.data\[316\] vssd1 vssd1 vccd1 vccd1 net3073 sky130_fd_sc_hd__dlygate4sd3_1
Xhold527 top.CPU.registers.data\[520\] vssd1 vssd1 vccd1 vccd1 net3084 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold538 top.CPU.registers.data\[12\] vssd1 vssd1 vccd1 vccd1 net3095 sky130_fd_sc_hd__dlygate4sd3_1
Xhold549 top.CPU.registers.data\[670\] vssd1 vssd1 vccd1 vccd1 net3106 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11318__A2 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08900_ net787 _04537_ _04538_ net715 vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__o211a_1
X_16009_ net2343 _02219_ net1060 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[809\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_98_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09880_ _03374_ _03442_ _05514_ _05515_ net371 vssd1 vssd1 vccd1 vccd1 _05519_ sky130_fd_sc_hd__a311oi_1
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07493__A top.SPI.busy vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08831_ _04331_ _04397_ _04469_ vssd1 vssd1 vccd1 vccd1 _04470_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_55_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11286__Y _06701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1205 top.CPU.registers.data\[413\] vssd1 vssd1 vccd1 vccd1 net3762 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1216 _02706_ vssd1 vssd1 vccd1 vccd1 net3773 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1227 top.I2C.data_out\[18\] vssd1 vssd1 vccd1 vccd1 net3784 sky130_fd_sc_hd__dlygate4sd3_1
X_08762_ net789 _04399_ _04400_ net742 vssd1 vssd1 vccd1 vccd1 _04401_ sky130_fd_sc_hd__o211a_1
X_13885__55 clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 net1524 sky130_fd_sc_hd__inv_2
Xhold1238 top.SPI.state\[3\] vssd1 vssd1 vccd1 vccd1 net3795 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11446__C net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1249 top.CPU.registers.data\[1007\] vssd1 vssd1 vccd1 vccd1 net3806 sky130_fd_sc_hd__dlygate4sd3_1
X_14740__910 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 net2379 sky130_fd_sc_hd__inv_2
XANTENNA__10829__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07713_ _03103_ _03153_ net1279 net1365 net1408 vssd1 vssd1 vccd1 vccd1 _03352_ sky130_fd_sc_hd__o2111a_1
X_08693_ top.CPU.alu.program_counter\[13\] net1037 vssd1 vssd1 vccd1 vccd1 _04332_
+ sky130_fd_sc_hd__or2_1
XFILLER_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout176_A _06795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07644_ _03277_ _03280_ _03282_ vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__a21oi_2
XFILLER_80_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07575_ top.CPU.registers.data\[575\] top.CPU.registers.data\[543\] net836 vssd1
+ vssd1 vccd1 vccd1 _03214_ sky130_fd_sc_hd__mux2_1
X_13947__117 clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 net1586 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_24_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout343_A _06771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09314_ net1363 net1041 net1039 net1047 vssd1 vssd1 vccd1 vccd1 _04953_ sky130_fd_sc_hd__o31a_1
XANTENNA__10057__A2 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11254__B2 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11889__S net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09245_ top.CPU.registers.data\[325\] net1310 net841 top.CPU.registers.data\[357\]
+ net737 vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout510_A _05669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_898 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1252_A net1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout229_X net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout608_A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11006__B2 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09176_ top.CPU.registers.data\[902\] net1316 net847 top.CPU.registers.data\[934\]
+ net718 vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_79_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16256__RESET_B net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12754__A1 top.CPU.alu.program_counter\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11557__A2 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08127_ net940 _03765_ vssd1 vssd1 vccd1 vccd1 _03766_ sky130_fd_sc_hd__or2_1
XFILLER_147_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07630__B1 _03262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08058_ top.CPU.registers.data\[660\] net1289 net1009 top.CPU.registers.data\[692\]
+ net906 vssd1 vssd1 vccd1 vccd1 _03697_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_112_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout598_X net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout977_A net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11309__A2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput47 net47 vssd1 vssd1 vccd1 vccd1 ADR_O[17] sky130_fd_sc_hd__buf_2
XFILLER_1_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput58 net58 vssd1 vssd1 vccd1 vccd1 ADR_O[29] sky130_fd_sc_hd__buf_2
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 DAT_O[10] sky130_fd_sc_hd__buf_2
XFILLER_115_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1305_X net1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10020_ net384 _05657_ vssd1 vssd1 vccd1 vccd1 _05659_ sky130_fd_sc_hd__or2_1
XFILLER_1_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout765_X net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07933__A1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14483__653 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 net2122 sky130_fd_sc_hd__inv_2
X_11971_ _06526_ net351 net182 net3145 vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout932_X net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12749__A top.CPU.alu.program_counter\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13710_ top.SPI.timem\[7\] _03058_ _07113_ vssd1 vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__o21ai_1
X_10922_ net478 net456 _06506_ net220 net2777 vssd1 vssd1 vccd1 vccd1 _02379_ sky130_fd_sc_hd__a32o_1
XANTENNA__11493__A1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07697__B1 net1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13641_ net3275 _07230_ net665 vssd1 vssd1 vccd1 vccd1 _02575_ sky130_fd_sc_hd__mux2_1
X_10853_ net410 _06138_ _06139_ _06455_ _06460_ vssd1 vssd1 vccd1 vccd1 _06461_ sky130_fd_sc_hd__o311a_1
X_14524__694 clknet_leaf_134_clk vssd1 vssd1 vccd1 vccd1 net2163 sky130_fd_sc_hd__inv_2
XFILLER_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16360_ clknet_leaf_32_clk _02569_ net1125 vssd1 vssd1 vccd1 vccd1 top.CPU.fetch.current_ra\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11245__A1 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13572_ top.CPU.addressnew\[9\] _03009_ net580 vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__mux2_1
XFILLER_13_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08646__C1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10784_ _05626_ _05628_ net382 vssd1 vssd1 vccd1 vccd1 _06395_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08110__A1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15311_ net1645 _01521_ net1097 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[111\]
+ sky130_fd_sc_hd__dfrtp_1
X_12523_ _06965_ _06966_ _07025_ _07030_ vssd1 vssd1 vccd1 vccd1 _07032_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_171_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16291_ clknet_leaf_109_clk _02500_ net1240 vssd1 vssd1 vccd1 vccd1 top.CPU.data_out\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_15242_ net1576 _01452_ net1094 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[42\]
+ sky130_fd_sc_hd__dfrtp_1
X_12454_ _03241_ _03369_ vssd1 vssd1 vccd1 vccd1 _06963_ sky130_fd_sc_hd__and2_1
XFILLER_126_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11405_ _06535_ net278 net268 net3355 vssd1 vssd1 vccd1 vccd1 _02106_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_10_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15173_ net1510 _01383_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r1_prev\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_12385_ top.CPU.addressnew\[29\] top.CPU.addressnew\[28\] top.CPU.addressnew\[31\]
+ top.CPU.addressnew\[30\] vssd1 vssd1 vccd1 vccd1 _06923_ sky130_fd_sc_hd__or4_1
XFILLER_125_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10756__B1 _06367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09793__A _05399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11336_ net3374 net288 net282 _05908_ vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__a22o_1
XANTENNA__08901__S net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11267_ net472 _06690_ vssd1 vssd1 vccd1 vccd1 _06691_ sky130_fd_sc_hd__nor2_1
XFILLER_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08177__A1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13006_ top.SPI.paroutput\[1\] _07429_ _07431_ net2669 vssd1 vssd1 vccd1 vccd1 _01207_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16399__Q top.CPU.handler.state\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10218_ net512 _05599_ _05851_ net447 _05435_ vssd1 vssd1 vccd1 vccd1 _05853_ sky130_fd_sc_hd__a221o_1
X_11198_ net3458 net297 _06656_ net323 vssd1 vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__a22o_1
XFILLER_94_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11720__A2 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10149_ net384 _05654_ _05785_ vssd1 vssd1 vccd1 vccd1 _05786_ sky130_fd_sc_hd__a21o_1
XANTENNA__11266__C net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09732__S net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14957_ clknet_leaf_89_clk top.SPI.nextwrx net1273 vssd1 vssd1 vccd1 vccd1 top.SPI.wrx
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13473__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11484__A1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08348__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15509_ net1843 _01719_ net1216 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[309\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12394__A net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16489_ clknet_leaf_41_clk _02651_ net1115 vssd1 vssd1 vccd1 vccd1 top.mmio.mem_data_i\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08652__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_695 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09030_ top.CPU.registers.data\[904\] net1314 net845 top.CPU.registers.data\[936\]
+ net716 vssd1 vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__a221o_1
XANTENNA__07860__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11539__A2 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09062__C1 net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold302 net50 vssd1 vssd1 vccd1 vccd1 net2859 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08404__A2 net1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold313 top.CPU.registers.data\[526\] vssd1 vssd1 vccd1 vccd1 net2870 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold324 top.CPU.registers.data\[558\] vssd1 vssd1 vccd1 vccd1 net2881 sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 top.SPI.paroutput\[21\] vssd1 vssd1 vccd1 vccd1 net2892 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08811__S net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold346 top.CPU.registers.data\[184\] vssd1 vssd1 vccd1 vccd1 net2903 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12841__B _03685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold357 top.CPU.registers.data\[555\] vssd1 vssd1 vccd1 vccd1 net2914 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09932_ _04295_ _04326_ vssd1 vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__or2_1
XANTENNA__13429__S net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold368 top.CPU.registers.data\[976\] vssd1 vssd1 vccd1 vccd1 net2925 sky130_fd_sc_hd__dlygate4sd3_1
Xhold379 top.CPU.registers.data\[3\] vssd1 vssd1 vccd1 vccd1 net2936 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout804 _03205_ vssd1 vssd1 vccd1 vccd1 net804 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09365__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout815 net822 vssd1 vssd1 vccd1 vccd1 net815 sky130_fd_sc_hd__buf_2
Xfanout826 net831 vssd1 vssd1 vccd1 vccd1 net826 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09863_ _05467_ _05500_ vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__nand2_2
Xfanout837 net839 vssd1 vssd1 vccd1 vccd1 net837 sky130_fd_sc_hd__clkbuf_4
X_14170__340 clknet_leaf_166_clk vssd1 vssd1 vccd1 vccd1 net1809 sky130_fd_sc_hd__inv_2
Xfanout848 net854 vssd1 vssd1 vccd1 vccd1 net848 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout293_A _06662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11172__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout859 net862 vssd1 vssd1 vccd1 vccd1 net859 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14467__637 clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 net2106 sky130_fd_sc_hd__inv_2
Xhold1002 top.CPU.registers.data\[936\] vssd1 vssd1 vccd1 vccd1 net3559 sky130_fd_sc_hd__dlygate4sd3_1
X_08814_ net904 _04450_ _04452_ net1366 vssd1 vssd1 vccd1 vccd1 _04453_ sky130_fd_sc_hd__a211o_1
XANTENNA__11711__A2 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1013 top.CPU.registers.data\[838\] vssd1 vssd1 vccd1 vccd1 net3570 sky130_fd_sc_hd__dlygate4sd3_1
X_09794_ _05399_ _05430_ vssd1 vssd1 vccd1 vccd1 _05433_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout1000_A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1024 top.CPU.registers.data\[882\] vssd1 vssd1 vccd1 vccd1 net3581 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1035 top.CPU.registers.data\[511\] vssd1 vssd1 vccd1 vccd1 net3592 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09117__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1046 top.CPU.registers.data\[612\] vssd1 vssd1 vccd1 vccd1 net3603 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1057 top.I2C.data_out\[15\] vssd1 vssd1 vccd1 vccd1 net3614 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08745_ top.CPU.registers.data\[589\] net1371 net968 top.CPU.registers.data\[621\]
+ net910 vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__o221a_1
XFILLER_39_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1068 top.CPU.registers.data\[135\] vssd1 vssd1 vccd1 vccd1 net3625 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout460_A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12569__A _06124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1079 top.CPU.registers.data\[992\] vssd1 vssd1 vccd1 vccd1 net3636 sky130_fd_sc_hd__dlygate4sd3_1
X_14211__381 clknet_leaf_114_clk vssd1 vssd1 vccd1 vccd1 net1850 sky130_fd_sc_hd__inv_2
XANTENNA_fanout558_A net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11473__A net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout179_X net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14508__678 clknet_leaf_190_clk vssd1 vssd1 vccd1 vccd1 net2147 sky130_fd_sc_hd__inv_2
XANTENNA__08876__C1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08258__S net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08676_ top.CPU.registers.data\[686\] net1291 vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__or2_1
XFILLER_27_979 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07627_ net1397 _03263_ vssd1 vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__nor2_1
XANTENNA__10089__A _03889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout725_A net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout346_X net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11227__A1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07558_ net1403 _03180_ _03183_ vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_153_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11778__A2 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07489_ top.I2C.read_byte_done vssd1 vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__inv_2
XANTENNA__10817__A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout513_X net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09228_ top.CPU.registers.data_out_r1_prev\[5\] net871 net640 _04866_ net713 vssd1
+ vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__o221a_1
XFILLER_42_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10095__Y _05733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09159_ _04797_ vssd1 vssd1 vccd1 vccd1 _04798_ sky130_fd_sc_hd__inv_2
XANTENNA__09053__C1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07603__A0 top.CPU.alu.program_counter\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14911__1081 clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 net2550 sky130_fd_sc_hd__inv_2
X_12170_ top.CPU.registers.data\[67\] net653 net149 net363 net356 vssd1 vssd1 vccd1
+ vccd1 _06853_ sky130_fd_sc_hd__o2111a_1
XFILLER_101_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout882_X net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11950__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11121_ net3581 net302 _06618_ net325 vssd1 vssd1 vccd1 vccd1 _02292_ sky130_fd_sc_hd__a22o_1
XFILLER_150_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12243__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10552__A net1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08159__A1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold880 top.CPU.registers.data\[204\] vssd1 vssd1 vccd1 vccd1 net3437 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13152__A1 net1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold891 top.CPU.registers.data\[689\] vssd1 vssd1 vccd1 vccd1 net3448 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_168_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09356__B1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13152__B2 top.CPU.alu.program_counter\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11052_ net3515 net368 _06584_ net318 vssd1 vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__a22o_1
XFILLER_153_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10003_ net413 _05616_ vssd1 vssd1 vccd1 vccd1 _05642_ sky130_fd_sc_hd__nor2_4
XANTENNA__11702__A2 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15860_ net2194 _02070_ net1120 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[660\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_130_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input21_A DAT_I[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15791_ net2125 _02001_ net1105 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[591\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13455__A2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08676__B net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_13_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09124__Y _04763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11954_ net516 _06500_ net345 _06775_ vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__a31o_1
XANTENNA__12198__B net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10905_ _06174_ _06468_ vssd1 vssd1 vccd1 vccd1 _06496_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_142_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_192_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_192_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11885_ _06230_ net3683 net189 vssd1 vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__mux2_1
XANTENNA__08882__A2 net1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_103_Left_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16412_ clknet_leaf_54_clk net2628 net1135 vssd1 vssd1 vccd1 vccd1 top.I2C.I2C_state\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13624_ net2666 _03040_ net581 vssd1 vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__mux2_1
X_10836_ net413 _06431_ _06439_ _06444_ vssd1 vssd1 vccd1 vccd1 _06445_ sky130_fd_sc_hd__a211o_2
XANTENNA__09788__A net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11769__A2 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13555_ top.CPU.addressnew\[2\] net579 _02998_ _02999_ vssd1 vssd1 vccd1 vccd1 _02532_
+ sky130_fd_sc_hd__a22o_1
XFILLER_158_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16343_ clknet_leaf_74_clk _02552_ net1158 vssd1 vssd1 vccd1 vccd1 top.CPU.addressnew\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_160_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10767_ _06342_ _06378_ net305 vssd1 vssd1 vccd1 vccd1 _06379_ sky130_fd_sc_hd__mux2_1
XFILLER_160_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12506_ _06999_ _07014_ _06998_ vssd1 vssd1 vccd1 vccd1 _07015_ sky130_fd_sc_hd__o21a_1
X_16274_ clknet_leaf_46_clk _02484_ net1137 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.toreg\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_173_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13486_ top.CPU.data_out\[0\] _05226_ net590 vssd1 vssd1 vccd1 vccd1 _02498_ sky130_fd_sc_hd__mux2_1
X_10698_ net572 net514 _06312_ vssd1 vssd1 vccd1 vccd1 _06314_ sky130_fd_sc_hd__and3_1
X_15225_ net1559 _01435_ net1238 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_12437_ net1340 top.I2C.output_state\[8\] top.I2C.output_state\[22\] vssd1 vssd1
+ vccd1 vccd1 _06955_ sky130_fd_sc_hd__a21o_1
XFILLER_32_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09595__A0 _05226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12194__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15156_ clknet_leaf_44_clk _01366_ net1124 vssd1 vssd1 vccd1 vccd1 top.I2C.data_out\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_12368_ top.I2C.I2C_state\[24\] top.I2C.I2C_state\[22\] vssd1 vssd1 vccd1 vccd1 _06909_
+ sky130_fd_sc_hd__nor2_1
XFILLER_5_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14930__Q top.CPU.alu.program_counter\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13249__S _02782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_112_Left_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14154__324 clknet_leaf_146_clk vssd1 vssd1 vccd1 vccd1 net1793 sky130_fd_sc_hd__inv_2
XFILLER_5_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11319_ net477 net519 _05694_ _06509_ vssd1 vssd1 vccd1 vccd1 _06710_ sky130_fd_sc_hd__and4_1
XANTENNA__11941__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15087_ clknet_leaf_53_clk _01300_ net1133 vssd1 vssd1 vccd1 vccd1 top.I2C.bit_timer_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12299_ net2580 _04633_ net1061 vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__mux2_1
XANTENNA__12006__X _06781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09028__A top.CPU.alu.program_counter\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13855__25 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 net1494 sky130_fd_sc_hd__inv_2
X_15989_ net2323 _02199_ net1217 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[789\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12249__A3 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08530_ top.CPU.registers.data\[80\] net1291 net1011 top.CPU.registers.data\[112\]
+ net953 vssd1 vssd1 vccd1 vccd1 _04169_ sky130_fd_sc_hd__a221o_1
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_121_Left_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08461_ top.CPU.registers.data\[977\] net1296 net1016 top.CPU.registers.data\[1009\]
+ net913 vssd1 vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_183_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_183_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08873__A2 net1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11209__A1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08392_ net908 _04030_ vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_34_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08625__A2 net1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout139_A _06126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08107__A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09013_ top.CPU.registers.data\[73\] net1369 net964 top.CPU.registers.data\[105\]
+ net900 vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__o221a_1
XFILLER_128_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09035__C1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12185__A2 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold110 net42 vssd1 vssd1 vccd1 vccd1 net2667 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold121 top.CPU.registers.data\[290\] vssd1 vssd1 vccd1 vccd1 net2678 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08541__S net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09050__A2 net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold132 top.CPU.registers.data\[302\] vssd1 vssd1 vccd1 vccd1 net2689 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11393__B1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_1_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07597__C1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold143 top.SPI.percount\[1\] vssd1 vssd1 vccd1 vccd1 net2700 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11932__A2 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold154 top.CPU.registers.data\[693\] vssd1 vssd1 vccd1 vccd1 net2711 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 top.CPU.registers.data\[47\] vssd1 vssd1 vccd1 vccd1 net2722 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold176 top.CPU.registers.data\[641\] vssd1 vssd1 vccd1 vccd1 net2733 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold187 top.CPU.handler.toreg\[29\] vssd1 vssd1 vccd1 vccd1 net2744 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout601 net603 vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__buf_4
XANTENNA__09338__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold198 top.SPI.parameters\[21\] vssd1 vssd1 vccd1 vccd1 net2755 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout612 net615 vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__buf_4
X_09915_ net401 _05055_ _05127_ _05550_ _05552_ vssd1 vssd1 vccd1 vccd1 _05554_ sky130_fd_sc_hd__a221o_1
XFILLER_132_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout623 _03340_ vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__buf_4
Xfanout634 _03244_ vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10091__B net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout645 net646 vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__clkbuf_4
XFILLER_58_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout296_X net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout675_A net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout656 net657 vssd1 vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__buf_2
XANTENNA__15412__RESET_B net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout667 net669 vssd1 vssd1 vccd1 vccd1 net667 sky130_fd_sc_hd__clkbuf_4
X_09846_ top.CPU.registers.data\[826\] top.CPU.registers.data\[794\] net1000 vssd1
+ vssd1 vccd1 vccd1 _05485_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_146_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout678 net684 vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1003_X net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout689 _03331_ vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08561__A1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09777_ top.CPU.registers.data\[699\] top.CPU.registers.data\[667\] net991 vssd1
+ vssd1 vccd1 vccd1 _05416_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout842_A net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout463_X net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_107_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08728_ top.CPU.registers.data\[461\] net1371 net967 top.CPU.registers.data\[493\]
+ net1364 vssd1 vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__o221a_1
XANTENNA__08849__C1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08313__A1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09510__B1 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11999__A2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08659_ top.CPU.registers.data\[462\] net1375 net981 top.CPU.registers.data\[494\]
+ net1364 vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout630_X net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10120__A1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_174_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_174_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08864__A2 net1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout728_X net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11670_ net462 _06485_ net237 net165 net2826 vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_120_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10621_ net444 _06236_ _06238_ _05283_ vssd1 vssd1 vccd1 vccd1 _06240_ sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_12_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14595__765 clknet_leaf_114_clk vssd1 vssd1 vccd1 vccd1 net2234 sky130_fd_sc_hd__inv_2
XANTENNA__08616__A2 _04254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13340_ top.I2C.data_out\[9\] net553 _02873_ net596 vssd1 vssd1 vccd1 vccd1 _02874_
+ sky130_fd_sc_hd__a22o_1
X_10552_ net1405 net576 net523 net143 vssd1 vssd1 vccd1 vccd1 _06175_ sky130_fd_sc_hd__and4_1
X_13271_ net3870 _02814_ _02820_ net1053 vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__a22o_1
X_10483_ _04192_ _05290_ vssd1 vssd1 vccd1 vccd1 _06108_ sky130_fd_sc_hd__nand2_1
X_15010_ clknet_leaf_97_clk _01255_ net1253 vssd1 vssd1 vccd1 vccd1 top.SPI.parameters\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_14138__308 clknet_leaf_163_clk vssd1 vssd1 vccd1 vccd1 net1777 sky130_fd_sc_hd__inv_2
X_12222_ net3899 net645 _06877_ vssd1 vssd1 vccd1 vccd1 _01450_ sky130_fd_sc_hd__o21a_1
XFILLER_135_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11384__B1 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11923__A2 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12153_ net3930 net646 _06844_ vssd1 vssd1 vccd1 vccd1 _01486_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_166_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11104_ net521 _05907_ vssd1 vssd1 vccd1 vccd1 _06610_ sky130_fd_sc_hd__nor2_1
X_12084_ net4020 net647 _06810_ vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__o21a_1
XFILLER_49_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11035_ _05768_ _05769_ _05770_ net536 vssd1 vssd1 vccd1 vccd1 _06577_ sky130_fd_sc_hd__o31a_2
X_15912_ net2246 _02122_ net1077 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[712\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08001__B1 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11687__A1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15843_ net2177 _02053_ net1206 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[643\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_94_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07760__C1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12986_ net3715 _07415_ net1342 vssd1 vssd1 vccd1 vccd1 _07417_ sky130_fd_sc_hd__a21oi_1
X_15774_ net2108 _01984_ net1240 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[574\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07738__S0 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12100__A2 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10111__A1 _03407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_165_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_165_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11937_ _06475_ net344 net229 net3209 vssd1 vssd1 vccd1 vccd1 _01631_ sky130_fd_sc_hd__a22o_1
X_11868_ _05847_ net3335 net191 vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__mux2_1
XANTENNA__12656__B _05156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14925__Q top.CPU.alu.program_counter\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13607_ net1348 _05988_ vssd1 vssd1 vccd1 vccd1 _03031_ sky130_fd_sc_hd__nand2_1
X_10819_ net440 _06428_ vssd1 vssd1 vccd1 vccd1 _06429_ sky130_fd_sc_hd__and2_1
XFILLER_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11799_ top.CPU.registers.data\[349\] net159 vssd1 vssd1 vccd1 vccd1 _06764_ sky130_fd_sc_hd__and2_1
XANTENNA__10457__A _06082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09804__A1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_08_1412 vssd1 vssd1 vccd1 vccd1 team_08_1412/HI ADR_O[26] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_31_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xteam_08_1423 vssd1 vssd1 vccd1 vccd1 team_08_1423/HI gpio_oeb[9] sky130_fd_sc_hd__conb_1
X_16326_ clknet_leaf_74_clk _02535_ net1159 vssd1 vssd1 vccd1 vccd1 top.CPU.addressnew\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_31_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13538_ top.CPU.data_out\[27\] net590 net339 _02989_ vssd1 vssd1 vccd1 vccd1 _02525_
+ sky130_fd_sc_hd__o22a_1
XFILLER_119_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xteam_08_1434 vssd1 vssd1 vccd1 vccd1 team_08_1434/HI gpio_out[19] sky130_fd_sc_hd__conb_1
XFILLER_158_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xteam_08_1445 vssd1 vssd1 vccd1 vccd1 team_08_1445/HI gpio_out[30] sky130_fd_sc_hd__conb_1
Xteam_08_1456 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] team_08_1456/LO sky130_fd_sc_hd__conb_1
Xteam_08_1467 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] team_08_1467/LO sky130_fd_sc_hd__conb_1
XFILLER_145_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09965__B _03371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13469_ net1396 net872 _02915_ net418 vssd1 vssd1 vccd1 vccd1 _02956_ sky130_fd_sc_hd__a31o_1
X_16257_ clknet_leaf_33_clk _02467_ net1123 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.toreg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12672__A top.CPU.alu.program_counter\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12167__A2 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15208_ net1542 _01418_ net1065 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_161_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16188_ net2522 _02398_ net1193 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[988\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11375__B1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11914__A2 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11288__A net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15139_ clknet_leaf_59_clk _01349_ net1140 vssd1 vssd1 vccd1 vccd1 top.I2C.data_out\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08791__A1 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09981__A _05123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07961_ top.CPU.registers.data\[568\] top.CPU.registers.data\[536\] net820 vssd1
+ vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__mux2_1
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11127__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09700_ top.CPU.registers.data\[473\] net1306 net1029 top.CPU.registers.data\[505\]
+ net922 vssd1 vssd1 vccd1 vccd1 _05339_ sky130_fd_sc_hd__a221o_1
XANTENNA__11678__A1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07892_ top.CPU.registers.data\[92\] net1332 net863 top.CPU.registers.data\[124\]
+ net778 vssd1 vssd1 vccd1 vccd1 _03531_ sky130_fd_sc_hd__a221o_1
XFILLER_67_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08543__A1 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09631_ _05127_ _05269_ vssd1 vssd1 vccd1 vccd1 _05270_ sky130_fd_sc_hd__or2_1
XFILLER_167_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09562_ net928 _05199_ _05200_ net951 vssd1 vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_69_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08513_ net745 _04145_ _04146_ net770 vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__o211a_1
X_14282__452 clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 net1921 sky130_fd_sc_hd__inv_2
X_14910__1080 clknet_leaf_152_clk vssd1 vssd1 vccd1 vccd1 net2549 sky130_fd_sc_hd__inv_2
X_09493_ top.CPU.registers.data\[417\] top.CPU.registers.data\[385\] top.CPU.registers.data\[289\]
+ top.CPU.registers.data\[257\] net998 net923 vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__mux4_1
XFILLER_23_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_156_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_156_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout256_A _06728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14579__749 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 net2218 sky130_fd_sc_hd__inv_2
X_08444_ top.CPU.registers.data\[657\] net1332 net863 top.CPU.registers.data\[689\]
+ net729 vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__a221o_1
XFILLER_169_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09221__A _04829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08375_ net792 _04010_ _04011_ net720 vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__o211a_1
XFILLER_23_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14323__493 clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 net1962 sky130_fd_sc_hd__inv_2
XANTENNA_fanout1165_A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11897__S net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09008__C1 net1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout211_X net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1332_A net1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12158__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09559__B1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08271__S net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout792_A net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11366__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11905__A2 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_148_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1218_X net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08782__A1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07585__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1407 top.CPU.control_unit.instruction\[8\] vssd1 vssd1 vccd1 vccd1 net1407
+ sky130_fd_sc_hd__buf_4
XFILLER_105_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout420 net423 vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__buf_4
Xfanout431 net432 vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout678_X net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout442 _05697_ vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__buf_2
Xfanout453 _03330_ vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__buf_4
XANTENNA__12866__B1 top.CPU.alu.program_counter\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout464 net467 vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_126_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout475 net477 vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout486 net497 vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__clkbuf_4
XFILLER_171_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_161_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09829_ top.CPU.registers.data\[58\] net1027 net945 vssd1 vssd1 vccd1 vccd1 _05468_
+ sky130_fd_sc_hd__a21o_1
XFILLER_19_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout497 _03188_ vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08300__A net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout845_X net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12840_ top.CPU.alu.program_counter\[19\] _07290_ net1360 vssd1 vssd1 vccd1 vccd1
+ _01182_ sky130_fd_sc_hd__mux2_1
XANTENNA__10892__A2 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16452__RESET_B net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10629__C1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12771_ top.CPU.alu.program_counter\[13\] top.CPU.alu.program_counter\[12\] _07208_
+ vssd1 vssd1 vccd1 vccd1 _07228_ sky130_fd_sc_hd__and3_1
XFILLER_15_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_147_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_147_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11722_ _06564_ net197 net420 net2878 vssd1 vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__a22o_1
XANTENNA__08393__S0 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15490_ net1824 _01700_ net1172 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[290\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08446__S net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11653_ _06314_ net196 net424 net3320 vssd1 vssd1 vccd1 vccd1 _01898_ sky130_fd_sc_hd__a22o_1
XFILLER_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10604_ _04467_ net508 _05677_ _04463_ vssd1 vssd1 vccd1 vccd1 _06224_ sky130_fd_sc_hd__o22a_1
XFILLER_156_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11584_ _06695_ net261 net248 net2709 vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__a22o_1
XANTENNA__09262__A2 net1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13323_ net1409 _02861_ net669 vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__mux2_1
XFILLER_10_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16111_ net2445 _02321_ net1095 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[911\]
+ sky130_fd_sc_hd__dfrtp_1
X_10535_ _04330_ _05569_ _05570_ vssd1 vssd1 vccd1 vccd1 _06158_ sky130_fd_sc_hd__a21o_1
XFILLER_11_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12492__A _04763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11600__S net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07586__A top.CPU.control_unit.instruction\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12149__A2 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13254_ net3888 _02805_ _02811_ _02803_ vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__a22o_1
XFILLER_109_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16042_ net2376 _02252_ net1084 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[842\]
+ sky130_fd_sc_hd__dfrtp_1
X_10466_ net415 _06091_ _05762_ vssd1 vssd1 vccd1 vccd1 _06092_ sky130_fd_sc_hd__o21ba_1
XFILLER_143_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11357__B1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12205_ net565 net362 _06677_ net169 top.CPU.registers.data\[49\] vssd1 vssd1 vccd1
+ vccd1 _06870_ sky130_fd_sc_hd__a32o_1
XFILLER_89_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13185_ top.I2C.I2C_state\[23\] top.I2C.I2C_state\[2\] _02765_ vssd1 vssd1 vccd1
+ vccd1 _02766_ sky130_fd_sc_hd__nor3_1
X_10397_ _05791_ _06023_ net402 vssd1 vssd1 vccd1 vccd1 _06026_ sky130_fd_sc_hd__mux2_1
XANTENNA__07576__A2 net1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12136_ _06057_ net361 net355 net173 top.CPU.registers.data\[84\] vssd1 vssd1 vccd1
+ vccd1 _06836_ sky130_fd_sc_hd__a32o_1
XFILLER_97_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12067_ net473 _06612_ _06802_ net177 net3883 vssd1 vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__a32o_1
X_11018_ net528 _06565_ vssd1 vssd1 vccd1 vccd1 _06566_ sky130_fd_sc_hd__nor2_1
XFILLER_65_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14266__436 clknet_leaf_161_clk vssd1 vssd1 vccd1 vccd1 net1905 sky130_fd_sc_hd__inv_2
X_15826_ net2160 _02036_ net1101 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[626\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12085__A1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_138_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_138_clk
+ sky130_fd_sc_hd__clkbuf_8
X_15757_ net2091 _01967_ net1077 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[557\]
+ sky130_fd_sc_hd__dfrtp_1
X_12969_ top.I2C.bit_timer_counter\[1\] top.I2C.bit_timer_counter\[0\] _07401_ top.I2C.bit_timer_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _07405_ sky130_fd_sc_hd__a31o_1
X_14010__180 clknet_leaf_159_clk vssd1 vssd1 vccd1 vccd1 net1649 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_47_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09312__Y _04951_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11832__A1 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15688_ net2022 _01898_ net1077 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[488\]
+ sky130_fd_sc_hd__dfrtp_1
X_14307__477 clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 net1946 sky130_fd_sc_hd__inv_2
XANTENNA__10458__Y _06085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09041__A net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09238__C1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08160_ net795 _03794_ _03795_ net749 vssd1 vssd1 vccd1 vccd1 _03799_ sky130_fd_sc_hd__o211a_1
XFILLER_174_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10399__B2 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11596__B1 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16309_ clknet_leaf_95_clk _02518_ net1247 vssd1 vssd1 vccd1 vccd1 top.CPU.data_out\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08091_ net799 _03728_ _03729_ net753 vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__o211a_1
XANTENNA__08461__B1 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10915__A net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload30 clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 clkload30/Y sky130_fd_sc_hd__inv_12
Xclkload41 clknet_leaf_185_clk vssd1 vssd1 vccd1 vccd1 clkload41/Y sky130_fd_sc_hd__inv_12
XFILLER_146_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload52 clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 clkload52/Y sky130_fd_sc_hd__inv_16
XANTENNA__11348__B1 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload63 clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 clkload63/Y sky130_fd_sc_hd__bufinv_16
Xclkload74 clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 clkload74/Y sky130_fd_sc_hd__inv_6
Xclkload85 clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 clkload85/Y sky130_fd_sc_hd__inv_8
XFILLER_133_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload96 clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 clkload96/Y sky130_fd_sc_hd__inv_16
XANTENNA__11899__A1 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11449__C _06085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_1_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08993_ net640 _04628_ _04631_ net702 _04625_ vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__o311a_1
X_07944_ top.CPU.registers.data\[344\] net1321 net852 top.CPU.registers.data\[376\]
+ net770 vssd1 vssd1 vccd1 vccd1 _03583_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_143_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08120__A net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07875_ top.CPU.registers.data\[924\] net1338 net870 top.CPU.registers.data\[956\]
+ net729 vssd1 vssd1 vccd1 vccd1 _03514_ sky130_fd_sc_hd__a221o_1
XANTENNA__10323__A1 _05793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout373_A net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11520__B1 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09614_ top.CPU.registers.data\[832\] net1315 net844 top.CPU.registers.data\[864\]
+ net741 vssd1 vssd1 vccd1 vccd1 _05253_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_67_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09545_ net803 _05183_ vssd1 vssd1 vccd1 vccd1 _05184_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_84_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_129_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_129_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09477__C1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout540_A net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout161_X net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout259_X net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout638_A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_174_Right_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09476_ top.CPU.registers.data\[802\] top.CPU.registers.data\[770\] net823 vssd1
+ vssd1 vccd1 vccd1 _05115_ sky130_fd_sc_hd__mux2_1
XFILLER_52_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08427_ top.CPU.registers.data\[241\] net1393 net825 top.CPU.registers.data\[209\]
+ net774 vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout805_A net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout426_X net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08358_ top.CPU.registers.data\[594\] net1317 net848 top.CPU.registers.data\[626\]
+ net742 vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__a221o_1
XANTENNA__08790__A top.CPU.alu.program_counter\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload2 clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clkload2/Y sky130_fd_sc_hd__inv_8
XFILLER_165_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09244__A2 net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11587__B1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08289_ top.CPU.registers.data\[51\] top.CPU.registers.data\[19\] net825 vssd1 vssd1
+ vccd1 vccd1 _03928_ sky130_fd_sc_hd__mux2_1
XFILLER_165_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1335_X net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10320_ net550 _03650_ _05679_ _03649_ vssd1 vssd1 vccd1 vccd1 _05952_ sky130_fd_sc_hd__o22a_1
XFILLER_109_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09097__S net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11339__B1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout795_X net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1443_X net4000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10251_ _05399_ _05467_ net374 vssd1 vssd1 vccd1 vccd1 _05885_ sky130_fd_sc_hd__mux2_1
XFILLER_152_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09401__C1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07558__A2 _03180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10182_ _05705_ _05706_ net382 vssd1 vssd1 vccd1 vccd1 _05818_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout962_X net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1204 net1205 vssd1 vssd1 vccd1 vccd1 net1204 sky130_fd_sc_hd__clkbuf_2
Xfanout1215 net1217 vssd1 vssd1 vccd1 vccd1 net1215 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07963__C1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1226 net1233 vssd1 vssd1 vccd1 vccd1 net1226 sky130_fd_sc_hd__clkbuf_2
Xfanout1237 net1240 vssd1 vssd1 vccd1 vccd1 net1237 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12251__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14990_ clknet_leaf_98_clk _01235_ net1254 vssd1 vssd1 vccd1 vccd1 top.SPI.paroutput\[29\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout250 _06733_ vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__clkbuf_8
Xfanout1248 net1249 vssd1 vssd1 vccd1 vccd1 net1248 sky130_fd_sc_hd__clkbuf_4
Xfanout1259 net1276 vssd1 vssd1 vccd1 vccd1 net1259 sky130_fd_sc_hd__clkbuf_4
Xfanout261 net262 vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__clkbuf_8
XFILLER_19_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout272 _06714_ vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__clkbuf_4
XFILLER_87_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout283 net284 vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__buf_4
Xfanout294 _06662_ vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08030__A net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07715__C1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11094__C net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09560__S net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15611_ net1945 _01821_ net1213 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[411\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11662__Y _06757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07730__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13590__B _06124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12823_ top.CPU.alu.program_counter\[18\] _04050_ vssd1 vssd1 vccd1 vccd1 _07275_
+ sky130_fd_sc_hd__and2_1
XANTENNA__12067__A1 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09468__C1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_141_Right_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15542_ net1876 _01752_ net1222 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[342\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11814__A1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12754_ top.CPU.alu.program_counter\[11\] _03118_ _07211_ _07212_ vssd1 vssd1 vccd1
+ vccd1 _01174_ sky130_fd_sc_hd__a22o_1
XANTENNA__08140__C1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11705_ _06537_ net203 net422 net3586 vssd1 vssd1 vccd1 vccd1 _01848_ sky130_fd_sc_hd__a22o_1
X_12685_ _07138_ _07140_ _07137_ vssd1 vssd1 vccd1 vccd1 _07150_ sky130_fd_sc_hd__a21bo_1
X_15473_ net1807 _01683_ net1189 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[273\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_139_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13567__A1 _03006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11636_ _05935_ net209 net427 net3286 vssd1 vssd1 vccd1 vccd1 _01915_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_42_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12934__B _03477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14651__821 clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 net2290 sky130_fd_sc_hd__inv_2
X_11567_ _06678_ net262 net247 net2732 vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__a22o_1
XANTENNA__10250__B1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13319__A1 _02858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07797__A2 net1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10518_ net410 _06138_ _06141_ _05673_ vssd1 vssd1 vccd1 vccd1 _06142_ sky130_fd_sc_hd__o2bb2a_1
X_13306_ net888 _02848_ vssd1 vssd1 vccd1 vccd1 _02849_ sky130_fd_sc_hd__and2_1
Xhold709 top.CPU.registers.data\[382\] vssd1 vssd1 vccd1 vccd1 net3266 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_170_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11498_ net479 net471 _06631_ net254 net3104 vssd1 vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__a32o_1
XFILLER_7_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13237_ top.I2C.data_out\[16\] net892 _06948_ vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__mux2_1
X_16025_ net2359 _02235_ net1244 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[825\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_170_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10449_ _03315_ _05295_ _05670_ _03988_ _06074_ vssd1 vssd1 vccd1 vccd1 _06076_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_161_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10173__C net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09735__S net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13168_ _06947_ _02752_ _02753_ _02751_ top.I2C.within_byte_counter_reading\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__a32o_1
XANTENNA__08859__B net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11750__B1 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07954__C1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_41_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12119_ _05809_ net355 net237 _06827_ vssd1 vssd1 vccd1 vccd1 _01503_ sky130_fd_sc_hd__a31o_1
X_13099_ _02713_ _02712_ top.SPI.count\[0\] vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1409 top.CPU.registers.data\[87\] vssd1 vssd1 vccd1 vccd1 net3966 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11502__B1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_176_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07660_ _03178_ _03288_ _03294_ vssd1 vssd1 vccd1 vccd1 _03299_ sky130_fd_sc_hd__a21o_1
XFILLER_66_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10856__A2 _06462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_56_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12058__A1 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15809_ net2143 _02019_ net1243 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[609\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09459__C1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07591_ top.CPU.registers.data\[383\] net1334 net865 top.CPU.registers.data\[351\]
+ net731 vssd1 vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__o221a_1
XFILLER_92_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09330_ top.CPU.registers.data\[804\] top.CPU.registers.data\[772\] net826 vssd1
+ vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__mux2_1
XFILLER_80_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09261_ top.CPU.registers.data\[37\] top.CPU.registers.data\[5\] net966 vssd1 vssd1
+ vccd1 vccd1 _04900_ sky130_fd_sc_hd__mux2_1
XANTENNA__09977__Y _05616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13007__B1 _07431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08212_ net677 _03849_ _03850_ net606 vssd1 vssd1 vccd1 vccd1 _03851_ sky130_fd_sc_hd__a31o_1
XFILLER_53_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09192_ top.CPU.registers.data\[390\] net1287 net1006 top.CPU.registers.data\[422\]
+ net904 vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__a221o_1
XFILLER_159_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_114_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08143_ net620 _03777_ _03778_ _03781_ vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__a31o_1
XANTENNA__07497__Y _03137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout121_A net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14394__564 clknet_leaf_161_clk vssd1 vssd1 vccd1 vccd1 net2033 sky130_fd_sc_hd__inv_2
XFILLER_162_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07788__A2 net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload130 clknet_leaf_172_clk vssd1 vssd1 vccd1 vccd1 clkload130/Y sky130_fd_sc_hd__inv_6
X_08074_ top.CPU.registers.data\[468\] net1288 net1008 top.CPU.registers.data\[500\]
+ net905 vssd1 vssd1 vccd1 vccd1 _03713_ sky130_fd_sc_hd__a221o_1
XFILLER_134_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload141 clknet_leaf_149_clk vssd1 vssd1 vccd1 vccd1 clkload141/Y sky130_fd_sc_hd__clkinv_8
Xclkload152 clknet_leaf_133_clk vssd1 vssd1 vccd1 vccd1 clkload152/Y sky130_fd_sc_hd__inv_6
XFILLER_134_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload163 clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 clkload163/Y sky130_fd_sc_hd__inv_8
XFILLER_162_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload174 clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 clkload174/Y sky130_fd_sc_hd__inv_12
Xclkload185 clknet_leaf_86_clk vssd1 vssd1 vccd1 vccd1 clkload185/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_129_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_779 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1030_A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1128_A net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08198__C1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout490_A net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11741__B1 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11476__A net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold14 top.CPU.registers.data_out_r2_prev\[21\] vssd1 vssd1 vccd1 vccd1 net2571 sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ top.CPU.registers.data\[73\] net1309 net840 top.CPU.registers.data\[105\]
+ net764 vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__a221o_1
XFILLER_152_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold25 top.CPU.registers.data_out_r1_prev\[15\] vssd1 vssd1 vccd1 vccd1 net2582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 top.CPU.registers.data_out_r2_prev\[25\] vssd1 vssd1 vccd1 vccd1 net2593 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold47 top.CPU.registers.data_out_r2_prev\[29\] vssd1 vssd1 vccd1 vccd1 net2604 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07960__A2 net1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold58 top.I2C.I2C_state\[15\] vssd1 vssd1 vccd1 vccd1 net2615 sky130_fd_sc_hd__dlygate4sd3_1
X_07927_ top.CPU.registers.data\[444\] net1026 net920 vssd1 vssd1 vccd1 vccd1 _03566_
+ sky130_fd_sc_hd__a21o_1
XFILLER_102_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold69 top.CPU.registers.data_out_r1_prev\[18\] vssd1 vssd1 vccd1 vccd1 net2626 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09698__C1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout376_X net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout755_A net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09162__A1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07858_ net932 _03495_ _03496_ net952 vssd1 vssd1 vccd1 vccd1 _03497_ sky130_fd_sc_hd__o211a_1
XANTENNA__07712__A2 net1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08370__C1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12049__A1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07616__D_N net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout922_A net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout543_X net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07789_ top.CPU.registers.data\[990\] net1302 net1023 top.CPU.registers.data\[1022\]
+ net919 vssd1 vssd1 vccd1 vccd1 _03428_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1285_X net1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13797__A1 top.CPU.handler.readout vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09528_ top.CPU.registers.data\[737\] top.CPU.registers.data\[705\] net838 vssd1
+ vssd1 vccd1 vccd1 _05167_ sky130_fd_sc_hd__mux2_1
XFILLER_40_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout710_X net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09459_ top.CPU.registers.data\[450\] net1324 net855 top.CPU.registers.data\[482\]
+ net773 vssd1 vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__a221o_1
XANTENNA__11272__A2 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08791__Y _04430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout808_X net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13630__S net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13549__A1 _06462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14635__805 clknet_leaf_148_clk vssd1 vssd1 vccd1 vccd1 net2274 sky130_fd_sc_hd__inv_2
X_12470_ net451 _03717_ vssd1 vssd1 vccd1 vccd1 _06979_ sky130_fd_sc_hd__nand2_1
XFILLER_40_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11421_ _06559_ net276 net267 net3501 vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_117_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11024__A2 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08425__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07779__A2 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11352_ net3771 net285 net276 _06272_ vssd1 vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__a22o_1
XFILLER_152_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11980__B1 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10303_ net3722 net227 net319 _05935_ vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__a22o_1
XANTENNA__10842__X _06450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11283_ net1405 _03170_ net513 net131 vssd1 vssd1 vccd1 vccd1 _06699_ sky130_fd_sc_hd__or4b_1
X_13022_ net3738 _07436_ net894 vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__mux2_1
XFILLER_112_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10234_ net386 _05624_ vssd1 vssd1 vccd1 vccd1 _05869_ sky130_fd_sc_hd__nand2_1
XANTENNA__11732__B1 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1001 net1002 vssd1 vssd1 vccd1 vccd1 net1001 sky130_fd_sc_hd__clkbuf_4
Xfanout1012 net1013 vssd1 vssd1 vccd1 vccd1 net1012 sky130_fd_sc_hd__clkbuf_4
X_10165_ _05790_ _05801_ net402 vssd1 vssd1 vccd1 vccd1 _05802_ sky130_fd_sc_hd__mux2_1
XFILLER_126_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1023 net1031 vssd1 vssd1 vccd1 vccd1 net1023 sky130_fd_sc_hd__clkbuf_4
Xfanout1034 net1036 vssd1 vssd1 vccd1 vccd1 net1034 sky130_fd_sc_hd__buf_4
Xfanout1045 _03156_ vssd1 vssd1 vccd1 vccd1 net1045 sky130_fd_sc_hd__buf_2
Xfanout1056 net1068 vssd1 vssd1 vccd1 vccd1 net1056 sky130_fd_sc_hd__buf_2
XANTENNA__07951__A2 net1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10096_ _03442_ net505 vssd1 vssd1 vccd1 vccd1 _05734_ sky130_fd_sc_hd__nor2_1
X_14973_ clknet_leaf_96_clk _01218_ net1247 vssd1 vssd1 vccd1 vccd1 top.SPI.paroutput\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1067 net1068 vssd1 vssd1 vccd1 vccd1 net1067 sky130_fd_sc_hd__clkbuf_2
Xfanout1078 net1079 vssd1 vssd1 vccd1 vccd1 net1078 sky130_fd_sc_hd__clkbuf_2
Xfanout1089 net1110 vssd1 vssd1 vccd1 vccd1 net1089 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09153__A1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10299__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10838__A2 _06445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08900__A1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08361__C1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12806_ top.CPU.alu.program_counter\[15\] top.CPU.alu.program_counter\[16\] _07240_
+ vssd1 vssd1 vccd1 vccd1 _07260_ sky130_fd_sc_hd__and3_1
X_13786_ net15 net1052 net887 net3737 vssd1 vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__a22o_1
X_10998_ net1405 _03170_ _06253_ vssd1 vssd1 vccd1 vccd1 _06553_ sky130_fd_sc_hd__or3b_1
XFILLER_37_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08113__C1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15525_ net1859 _01735_ net1086 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[325\]
+ sky130_fd_sc_hd__dfrtp_1
X_12737_ _07167_ _07178_ _07179_ _07183_ _07176_ vssd1 vssd1 vccd1 vccd1 _07197_ sky130_fd_sc_hd__o311a_1
XFILLER_15_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14081__251 clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 net1720 sky130_fd_sc_hd__inv_2
X_15456_ net1790 _01666_ net1094 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[256\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_129_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14378__548 clknet_leaf_145_clk vssd1 vssd1 vccd1 vccd1 net2017 sky130_fd_sc_hd__inv_2
X_12668_ top.CPU.alu.program_counter\[2\] top.CPU.alu.program_counter\[3\] vssd1 vssd1
+ vccd1 vccd1 _07135_ sky130_fd_sc_hd__xor2_1
XANTENNA__12664__B _05021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12212__A1 _06213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11619_ _06311_ net3084 net213 vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__mux2_1
X_15387_ net1721 _01597_ net1214 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[187\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09613__C1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10223__A0 _03544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12599_ _03139_ top.SPI.count\[3\] top.SPI.count\[2\] _03141_ _07099_ vssd1 vssd1
+ vccd1 vccd1 _07100_ sky130_fd_sc_hd__o221a_1
XFILLER_156_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14122__292 clknet_leaf_146_clk vssd1 vssd1 vccd1 vccd1 net1761 sky130_fd_sc_hd__inv_2
Xhold506 top.CPU.registers.data\[317\] vssd1 vssd1 vccd1 vccd1 net3063 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12951__Y _07391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10774__A1 _03315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14419__589 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 net2058 sky130_fd_sc_hd__inv_2
XFILLER_143_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11971__B1 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold517 top.CPU.registers.data\[978\] vssd1 vssd1 vccd1 vccd1 net3074 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold528 top.SPI.paroutput\[14\] vssd1 vssd1 vccd1 vccd1 net3085 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold539 top.CPU.registers.data\[674\] vssd1 vssd1 vccd1 vccd1 net3096 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_98_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16008_ net2342 _02218_ net1088 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[808\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11723__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11296__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08830_ _04466_ _04467_ vssd1 vssd1 vccd1 vccd1 _04469_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_55_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1206 top.CPU.registers.data\[70\] vssd1 vssd1 vccd1 vccd1 net3763 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12279__A1 _05397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08761_ top.CPU.registers.data\[716\] net814 net767 _04398_ vssd1 vssd1 vccd1 vccd1
+ _04400_ sky130_fd_sc_hd__a211o_1
Xhold1217 top.CPU.registers.data\[52\] vssd1 vssd1 vccd1 vccd1 net3774 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1228 top.CPU.registers.data\[341\] vssd1 vssd1 vccd1 vccd1 net3785 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1239 top.CPU.registers.data_out_r1_prev\[17\] vssd1 vssd1 vccd1 vccd1 net3796
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07712_ top.CPU.registers.data\[127\] net1307 net1030 top.CPU.registers.data\[95\]
+ net681 vssd1 vssd1 vccd1 vccd1 _03351_ sky130_fd_sc_hd__o221a_1
X_08692_ _04260_ _04330_ vssd1 vssd1 vccd1 vccd1 _04331_ sky130_fd_sc_hd__or2_1
XANTENNA__09695__A2 net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07643_ _03262_ _03264_ _03281_ vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__nor3_1
XFILLER_53_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout169_A net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14820__990 clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 net2459 sky130_fd_sc_hd__inv_2
X_07574_ net1047 _03163_ net1038 _03112_ vssd1 vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__a31o_1
X_13986__156 clknet_leaf_147_clk vssd1 vssd1 vccd1 vccd1 net1625 sky130_fd_sc_hd__inv_2
XANTENNA__08892__X _04531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09313_ _04944_ _04950_ vssd1 vssd1 vccd1 vccd1 _04952_ sky130_fd_sc_hd__and2_2
XFILLER_80_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11254__A2 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout336_A net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13450__S net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_60_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_166_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09244_ top.CPU.registers.data\[229\] net1387 net806 top.CPU.registers.data\[197\]
+ net715 vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__a221o_1
XFILLER_31_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10585__A1_N _04392_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11006__A2 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09175_ top.CPU.registers.data\[806\] top.CPU.registers.data\[774\] net814 vssd1
+ vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__mux2_1
XANTENNA__08407__B1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09604__C1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout124_X net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout503_A net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08116__Y _03755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1245_A net1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08126_ top.CPU.registers.data\[53\] top.CPU.registers.data\[21\] net993 vssd1 vssd1
+ vccd1 vccd1 _03765_ sky130_fd_sc_hd__mux2_1
XANTENNA__10214__B1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12754__A2 _03118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08057_ top.CPU.registers.data\[564\] top.CPU.registers.data\[532\] net980 vssd1
+ vssd1 vccd1 vccd1 _03696_ sky130_fd_sc_hd__mux2_1
XANTENNA__09883__B _03544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1033_X net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput48 net48 vssd1 vssd1 vccd1 vccd1 ADR_O[18] sky130_fd_sc_hd__buf_2
Xoutput59 net59 vssd1 vssd1 vccd1 vccd1 ADR_O[2] sky130_fd_sc_hd__buf_2
XFILLER_150_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout872_A net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout493_X net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11714__B1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07918__C1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08186__A2 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08591__C1 net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08959_ top.CPU.control_unit.instruction\[30\] _04596_ _04597_ vssd1 vssd1 vccd1
+ vccd1 _04598_ sky130_fd_sc_hd__o21a_1
XANTENNA__13467__B1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout660_X net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout758_X net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13930__100 clknet_leaf_147_clk vssd1 vssd1 vccd1 vccd1 net1569 sky130_fd_sc_hd__inv_2
X_11970_ net570 net540 _06751_ net1403 vssd1 vssd1 vccd1 vccd1 _06777_ sky130_fd_sc_hd__or4b_4
XANTENNA__09686__A2 net1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_16_Left_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08343__C1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10921_ net144 net435 vssd1 vssd1 vccd1 vccd1 _06506_ sky130_fd_sc_hd__and2_1
XFILLER_84_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11493__A2 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout925_X net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13640_ net3953 _07221_ net665 vssd1 vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__mux2_1
X_10852_ net399 _06296_ _06459_ _06141_ vssd1 vssd1 vccd1 vccd1 _06460_ sky130_fd_sc_hd__o211ai_1
X_14065__235 clknet_leaf_186_clk vssd1 vssd1 vccd1 vccd1 net1704 sky130_fd_sc_hd__inv_2
XANTENNA__09438__A2 net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12956__A_N net1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13571_ top.CPU.alu.program_counter\[9\] _06288_ net1349 vssd1 vssd1 vccd1 vccd1
+ _03009_ sky130_fd_sc_hd__mux2_1
X_10783_ _05619_ _05629_ vssd1 vssd1 vccd1 vccd1 _06394_ sky130_fd_sc_hd__nor2_1
XFILLER_25_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11245__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_51_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_157_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15310_ net1644 _01520_ net1104 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[110\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_169_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12522_ _06962_ _06963_ _06968_ _06995_ vssd1 vssd1 vccd1 vccd1 _07031_ sky130_fd_sc_hd__o22a_1
X_16290_ clknet_leaf_107_clk _02499_ net1248 vssd1 vssd1 vccd1 vccd1 top.CPU.data_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_157_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14106__276 clknet_leaf_162_clk vssd1 vssd1 vccd1 vccd1 net1745 sky130_fd_sc_hd__inv_2
X_15241_ net1575 _01451_ net1063 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12453_ _03405_ _03439_ _03241_ _03369_ vssd1 vssd1 vccd1 vccd1 _06962_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__07578__B net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11404_ _06534_ net284 net270 net3033 vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__a22o_1
XFILLER_166_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12384_ _06918_ _06920_ _06921_ vssd1 vssd1 vccd1 vccd1 _06922_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_10_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09071__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15172_ net1509 _01382_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r1_prev\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_10_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10756__A1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11335_ net3854 net287 net281 _05880_ vssd1 vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__a22o_1
XFILLER_141_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09285__S net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11266_ net513 _06313_ net540 vssd1 vssd1 vccd1 vccd1 _06690_ sky130_fd_sc_hd__or3_1
XANTENNA__11705__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10217_ _05503_ _05598_ net445 vssd1 vssd1 vccd1 vccd1 _05852_ sky130_fd_sc_hd__a21oi_1
XFILLER_140_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13005_ top.SPI.paroutput\[0\] _07429_ _07431_ net2718 vssd1 vssd1 vccd1 vccd1 _01206_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11197_ net142 net429 vssd1 vssd1 vccd1 vccd1 _06656_ sky130_fd_sc_hd__and2_1
XANTENNA__12005__A net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14763__933 clknet_leaf_149_clk vssd1 vssd1 vccd1 vccd1 net2402 sky130_fd_sc_hd__inv_2
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07924__A2 net1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10148_ net308 _05784_ vssd1 vssd1 vccd1 vccd1 _05785_ sky130_fd_sc_hd__and2_1
XANTENNA__13458__A0 top.CPU.handler.toreg\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14956_ clknet_leaf_53_clk _01202_ net1133 vssd1 vssd1 vccd1 vccd1 top.I2C.bit_timer_counter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10079_ _05713_ _05716_ net383 vssd1 vssd1 vccd1 vccd1 _05717_ sky130_fd_sc_hd__mux2_1
XANTENNA__09677__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12130__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14804__974 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 net2443 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_50_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14928__Q top.CPU.alu.program_counter\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12681__A1 top.CPU.alu.program_counter\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11484__A2 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16626_ top.SPI.dcx vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__clkbuf_1
XFILLER_35_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13769_ net28 net1049 net884 net3968 vssd1 vssd1 vccd1 vccd1 _02650_ sky130_fd_sc_hd__o22a_1
XANTENNA__09834__C1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_42_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_94_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15508_ net1842 _01718_ net1120 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[308\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11787__A3 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16488_ clknet_leaf_41_clk _02650_ net1115 vssd1 vssd1 vccd1 vccd1 top.mmio.mem_data_i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_148_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10995__B2 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15439_ net1773 _01649_ net1096 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[239\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_96_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09062__B1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold303 top.CPU.fetch.current_ra\[31\] vssd1 vssd1 vccd1 vccd1 net2860 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold314 top.CPU.registers.data\[27\] vssd1 vssd1 vccd1 vccd1 net2871 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold325 top.SPI.parameters\[24\] vssd1 vssd1 vccd1 vccd1 net2882 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold336 top.CPU.registers.data\[327\] vssd1 vssd1 vccd1 vccd1 net2893 sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 top.CPU.registers.data\[813\] vssd1 vssd1 vccd1 vccd1 net2904 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold358 top.CPU.registers.data\[476\] vssd1 vssd1 vccd1 vccd1 net2915 sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 top.I2C.output_state\[21\] vssd1 vssd1 vccd1 vccd1 net2926 sky130_fd_sc_hd__dlygate4sd3_1
X_09931_ _04295_ _04326_ vssd1 vssd1 vccd1 vccd1 _05570_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_74_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout805 net806 vssd1 vssd1 vccd1 vccd1 net805 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08168__A2 net1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout816 net817 vssd1 vssd1 vccd1 vccd1 net816 sky130_fd_sc_hd__clkbuf_4
X_09862_ _05467_ _05500_ vssd1 vssd1 vccd1 vccd1 _05501_ sky130_fd_sc_hd__nor2_1
Xfanout827 net828 vssd1 vssd1 vccd1 vccd1 net827 sky130_fd_sc_hd__clkbuf_4
Xfanout838 net839 vssd1 vssd1 vccd1 vccd1 net838 sky130_fd_sc_hd__buf_2
XANTENNA__11172__A1 net1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout849 net850 vssd1 vssd1 vccd1 vccd1 net849 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08573__C1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07915__A2 net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08813_ top.CPU.registers.data\[652\] net1013 net935 _04451_ vssd1 vssd1 vccd1 vccd1
+ _04452_ sky130_fd_sc_hd__o211a_1
Xhold1003 top.CPU.registers.data\[210\] vssd1 vssd1 vccd1 vccd1 net3560 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09793_ _05399_ _05430_ vssd1 vssd1 vccd1 vccd1 _05432_ sky130_fd_sc_hd__nor2_1
Xhold1014 top.I2C.data_out\[17\] vssd1 vssd1 vccd1 vccd1 net3571 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1025 top.CPU.registers.data\[640\] vssd1 vssd1 vccd1 vccd1 net3582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1036 top.CPU.registers.data\[704\] vssd1 vssd1 vccd1 vccd1 net3593 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout286_A _06712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1047 top.CPU.registers.data\[320\] vssd1 vssd1 vccd1 vccd1 net3604 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08744_ top.CPU.registers.data\[717\] net1371 net968 top.CPU.registers.data\[749\]
+ net926 vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__o221a_1
Xhold1058 top.CPU.registers.data\[764\] vssd1 vssd1 vccd1 vccd1 net3615 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1069 top.I2C.I2C_state\[11\] vssd1 vssd1 vccd1 vccd1 net3626 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08325__C1 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09668__A2 net1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12569__B _06210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08675_ top.CPU.registers.data\[558\] top.CPU.registers.data\[526\] net982 vssd1
+ vssd1 vccd1 vccd1 _04314_ sky130_fd_sc_hd__mux2_1
X_14049__219 clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 net1688 sky130_fd_sc_hd__inv_2
XANTENNA__08876__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11475__A2 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10683__B1 _06139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08340__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07626_ _03263_ _03264_ vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__nand2_1
X_13836__6 clknet_leaf_190_clk vssd1 vssd1 vccd1 vccd1 net1475 sky130_fd_sc_hd__inv_2
XFILLER_26_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10089__B net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13621__A0 top.CPU.alu.program_counter\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07557_ net1403 _03180_ _03183_ vssd1 vssd1 vccd1 vccd1 _03196_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11227__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout620_A net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout241_X net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout339_X net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_33_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout718_A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07488_ net3838 vssd1 vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__inv_2
XFILLER_50_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10817__B _06426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09840__A2 net1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09227_ top.CPU.registers.data\[805\] top.CPU.registers.data\[773\] top.CPU.registers.data\[549\]
+ top.CPU.registers.data\[517\] net806 net690 vssd1 vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__mux4_1
XANTENNA__10309__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07851__A1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout506_X net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12188__B1 _03185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09158_ _04765_ _04794_ vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_131_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08109_ top.CPU.registers.data\[853\] net1330 net861 top.CPU.registers.data\[885\]
+ net776 vssd1 vssd1 vccd1 vccd1 _03748_ sky130_fd_sc_hd__a221o_1
XANTENNA__07603__A1 _03241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_863 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09089_ top.CPU.control_unit.instruction\[28\] _04596_ _04597_ vssd1 vssd1 vccd1
+ vccd1 _04728_ sky130_fd_sc_hd__o21a_1
XFILLER_174_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14450__620 clknet_leaf_193_clk vssd1 vssd1 vccd1 vccd1 net2089 sky130_fd_sc_hd__inv_2
XFILLER_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11120_ net516 _06106_ vssd1 vssd1 vccd1 vccd1 _06618_ sky130_fd_sc_hd__nor2_1
XFILLER_174_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14747__917 clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 net2386 sky130_fd_sc_hd__inv_2
Xhold870 top.CPU.registers.data\[387\] vssd1 vssd1 vccd1 vccd1 net3427 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10552__B net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout875_X net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold881 top.SPI.parameters\[4\] vssd1 vssd1 vccd1 vccd1 net3438 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_168_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13152__A2 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11051_ _06033_ net538 vssd1 vssd1 vccd1 vccd1 _06584_ sky130_fd_sc_hd__and2_1
Xhold892 top.CPU.registers.data\[784\] vssd1 vssd1 vccd1 vccd1 net3449 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_168_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10002_ _05632_ _05640_ net401 vssd1 vssd1 vccd1 vccd1 _05641_ sky130_fd_sc_hd__mux2_1
XANTENNA__08564__C1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07906__A2 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_129_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15790_ net2124 _02000_ net1106 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[590\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_18_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12112__B1 _06770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input14_A DAT_I[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08867__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11953_ top.CPU.registers.data\[206\] net230 vssd1 vssd1 vccd1 vccd1 _06775_ sky130_fd_sc_hd__and2_1
XFILLER_91_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08331__A2 net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10904_ net486 net462 _06495_ net221 net2925 vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_142_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11884_ _06212_ net3445 net188 vssd1 vssd1 vccd1 vccd1 _01679_ sky130_fd_sc_hd__mux2_1
XFILLER_60_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16411_ clknet_leaf_53_clk net2781 net1135 vssd1 vssd1 vccd1 vccd1 top.I2C.I2C_state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_13623_ top.CPU.alu.program_counter\[30\] _05767_ net1350 vssd1 vssd1 vccd1 vccd1
+ _03040_ sky130_fd_sc_hd__mux2_1
X_10835_ _06442_ _06443_ _06140_ vssd1 vssd1 vccd1 vccd1 _06444_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12495__A _05084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13090__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_24_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_15_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11603__S net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16342_ clknet_leaf_75_clk _02551_ net1158 vssd1 vssd1 vccd1 vccd1 top.CPU.addressnew\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13554_ _03100_ _03137_ net579 vssd1 vssd1 vccd1 vccd1 _02999_ sky130_fd_sc_hd__a21oi_1
XFILLER_34_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10766_ _05706_ _05708_ vssd1 vssd1 vccd1 vccd1 _06378_ sky130_fd_sc_hd__nor2_1
XANTENNA__09292__B1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10977__B2 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12505_ _07009_ _07010_ _07013_ _07012_ _07000_ vssd1 vssd1 vccd1 vccd1 _07014_ sky130_fd_sc_hd__o311a_1
X_16273_ clknet_leaf_45_clk _02483_ net1138 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.toreg\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13485_ _03137_ _03246_ _03288_ vssd1 vssd1 vccd1 vccd1 _02964_ sky130_fd_sc_hd__nor3_1
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10697_ net438 _06311_ vssd1 vssd1 vccd1 vccd1 _06313_ sky130_fd_sc_hd__nand2_1
XANTENNA__12179__B1 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15224_ net1558 _01434_ net1102 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_12436_ net1054 _06954_ vssd1 vssd1 vccd1 vccd1 _00055_ sky130_fd_sc_hd__and2_1
XANTENNA__14923__RESET_B net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11926__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08398__A2 net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15155_ clknet_leaf_42_clk _01365_ net1117 vssd1 vssd1 vccd1 vccd1 top.I2C.data_out\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12367_ top.I2C.initiate_read_bit _06902_ vssd1 vssd1 vccd1 vccd1 _06908_ sky130_fd_sc_hd__nor2_1
XANTENNA__10743__A net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14193__363 clknet_leaf_180_clk vssd1 vssd1 vccd1 vccd1 net1832 sky130_fd_sc_hd__inv_2
X_11318_ net3460 net289 net357 _06311_ vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__a22o_1
XANTENNA__11558__B _05990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15086_ clknet_leaf_53_clk _01299_ net1133 vssd1 vssd1 vccd1 vccd1 top.I2C.bit_timer_state\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_12298_ _04566_ _06887_ _06890_ vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_91_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09347__A1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11249_ net472 _06679_ vssd1 vssd1 vccd1 vccd1 _06680_ sky130_fd_sc_hd__nor2_1
XANTENNA__12351__B1 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10362__C1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11574__A net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08570__A2 net1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15782__RESET_B net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15988_ net2322 _02198_ net1120 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[788\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12103__B1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14939_ clknet_leaf_75_clk _01185_ net1158 vssd1 vssd1 vccd1 vccd1 top.CPU.alu.program_counter\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11106__A_N _05933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15029__RESET_B net1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08460_ top.CPU.registers.data\[849\] net1296 net1016 top.CPU.registers.data\[881\]
+ net938 vssd1 vssd1 vccd1 vccd1 _04099_ sky130_fd_sc_hd__a221o_1
XANTENNA__09979__A net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11209__A2 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08391_ top.CPU.registers.data\[690\] top.CPU.registers.data\[658\] net982 vssd1
+ vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_15_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_50_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10968__B2 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09822__A2 net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09012_ top.CPU.registers.data\[169\] top.CPU.registers.data\[137\] top.CPU.registers.data\[41\]
+ top.CPU.registers.data\[9\] net965 net900 vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__mux4_1
XFILLER_136_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09035__B1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14434__604 clknet_leaf_140_clk vssd1 vssd1 vccd1 vccd1 net2073 sky130_fd_sc_hd__inv_2
XFILLER_145_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11917__B1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09586__A1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold100 top.CPU.registers.data\[394\] vssd1 vssd1 vccd1 vccd1 net2657 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09130__S0 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10653__A net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold111 top.CPU.registers.data\[703\] vssd1 vssd1 vccd1 vccd1 net2668 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout201_A net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold122 top.CPU.registers.data\[63\] vssd1 vssd1 vccd1 vccd1 net2679 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_160_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold133 top.SPI.paroutput\[8\] vssd1 vssd1 vccd1 vccd1 net2690 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07597__B1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold144 top.CPU.registers.data\[305\] vssd1 vssd1 vccd1 vccd1 net2701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 top.CPU.registers.data\[557\] vssd1 vssd1 vccd1 vccd1 net2712 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 top.SPI.parameters\[26\] vssd1 vssd1 vccd1 vccd1 net2723 sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 top.I2C.bit_timer_counter\[5\] vssd1 vssd1 vccd1 vccd1 net2734 sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 net68 vssd1 vssd1 vccd1 vccd1 net2745 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09338__A1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout602 net603 vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__clkbuf_4
Xhold199 top.SPI.parameters\[11\] vssd1 vssd1 vccd1 vccd1 net2756 sky130_fd_sc_hd__dlygate4sd3_1
X_09914_ _05551_ _05552_ vssd1 vssd1 vccd1 vccd1 _05553_ sky130_fd_sc_hd__nor2_1
Xfanout613 net615 vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__clkbuf_4
Xfanout624 net626 vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1110_A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout635 net636 vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__clkbuf_8
XFILLER_98_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08546__C1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout646 net650 vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__buf_2
XANTENNA__13683__B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input6_A DAT_I[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09845_ top.CPU.registers.data\[986\] net1305 net1027 top.CPU.registers.data\[1018\]
+ net921 vssd1 vssd1 vccd1 vccd1 _05484_ sky130_fd_sc_hd__a221o_1
Xfanout657 net658 vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout668 net669 vssd1 vssd1 vccd1 vccd1 net668 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout191_X net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout570_A net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11696__A2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout679 net680 vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout668_A net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout289_X net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09776_ top.CPU.registers.data\[571\] top.CPU.registers.data\[539\] net991 vssd1
+ vssd1 vccd1 vccd1 _05415_ sky130_fd_sc_hd__mux2_1
XANTENNA__08269__S net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08727_ top.CPU.registers.data\[429\] top.CPU.registers.data\[397\] top.CPU.registers.data\[301\]
+ top.CPU.registers.data\[269\] net967 net1280 vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout456_X net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout835_A net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_87_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ top.CPU.registers.data\[430\] top.CPU.registers.data\[398\] top.CPU.registers.data\[302\]
+ top.CPU.registers.data\[270\] net981 net1282 vssd1 vssd1 vccd1 vccd1 _04297_ sky130_fd_sc_hd__mux4_1
XFILLER_14_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07609_ top.CPU.control_unit.instruction\[14\] net1397 vssd1 vssd1 vccd1 vccd1 _03248_
+ sky130_fd_sc_hd__nor2_2
XFILLER_53_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout623_X net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08589_ top.CPU.registers.data\[431\] top.CPU.registers.data\[399\] top.CPU.registers.data\[303\]
+ top.CPU.registers.data\[271\] net974 net1281 vssd1 vssd1 vccd1 vccd1 _04228_ sky130_fd_sc_hd__mux4_1
XFILLER_53_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1365_X net1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10408__B1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10620_ _04603_ _06235_ net444 vssd1 vssd1 vccd1 vccd1 _06239_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_12_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09813__A2 net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10959__B2 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10551_ net439 _06173_ vssd1 vssd1 vccd1 vccd1 _06174_ sky130_fd_sc_hd__nand2_1
XANTENNA__11620__A2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09828__S net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13270_ top.I2C.data_out\[1\] net891 _02774_ vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__mux2_1
XFILLER_108_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08732__S net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10482_ net3554 net228 net313 _06107_ vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout992_X net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11908__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09577__A1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14177__347 clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 net1816 sky130_fd_sc_hd__inv_2
X_12221_ _06312_ net542 _06796_ net168 top.CPU.registers.data\[40\] vssd1 vssd1 vccd1
+ vccd1 _06877_ sky130_fd_sc_hd__a32o_1
XANTENNA__12254__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07588__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08785__C1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12152_ _06231_ net360 net354 net172 top.CPU.registers.data\[76\] vssd1 vssd1 vccd1
+ vccd1 _06844_ sky130_fd_sc_hd__a32o_1
XANTENNA__09129__A net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11103_ net489 net466 _06609_ net303 net3333 vssd1 vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__a32o_1
XANTENNA__09329__A1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14218__388 clknet_leaf_146_clk vssd1 vssd1 vccd1 vccd1 net1857 sky130_fd_sc_hd__inv_2
X_12083_ _06621_ net245 net176 top.CPU.registers.data\[111\] vssd1 vssd1 vccd1 vccd1
+ _06810_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_34_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08537__C1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07872__A _03476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15911_ net2245 _02121_ net1198 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[711\]
+ sky130_fd_sc_hd__dfrtp_1
X_11034_ net325 net138 net539 net368 net2696 vssd1 vssd1 vccd1 vccd1 _02337_ sky130_fd_sc_hd__a32o_1
XFILLER_131_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15842_ net2176 _02052_ net1171 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[642\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07760__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15773_ net2107 _01983_ net1121 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[573\]
+ sky130_fd_sc_hd__dfrtp_1
X_12985_ top.I2C.bit_timer_counter\[3\] top.I2C.bit_timer_counter\[7\] _07406_ vssd1
+ vssd1 vccd1 vccd1 _07416_ sky130_fd_sc_hd__and3_1
XFILLER_18_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07738__S1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11936_ _06474_ net350 net232 net3533 vssd1 vssd1 vccd1 vccd1 _01632_ sky130_fd_sc_hd__a22o_1
XANTENNA__10111__A2 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07811__S net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11867_ _05808_ net3359 net189 vssd1 vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__mux2_1
X_13606_ net2909 _03030_ net583 vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__mux2_1
XANTENNA__13061__A1 top.CPU.data_out\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10818_ top.CPU.fetch.current_ra\[2\] net1041 net633 top.CPU.handler.toreg\[2\] _06427_
+ vssd1 vssd1 vccd1 vccd1 _06428_ sky130_fd_sc_hd__a221o_4
XANTENNA__09265__B1 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11798_ net137 net3540 net158 vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__mux2_1
Xteam_08_1413 vssd1 vssd1 vccd1 vccd1 team_08_1413/HI ADR_O[27] sky130_fd_sc_hd__conb_1
X_16325_ clknet_leaf_67_clk _02534_ net1241 vssd1 vssd1 vccd1 vccd1 top.CPU.addressnew\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_158_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xteam_08_1424 vssd1 vssd1 vccd1 vccd1 team_08_1424/HI gpio_oeb[10] sky130_fd_sc_hd__conb_1
X_13537_ _05428_ net585 vssd1 vssd1 vccd1 vccd1 _02989_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_31_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xteam_08_1435 vssd1 vssd1 vccd1 vccd1 team_08_1435/HI gpio_out[20] sky130_fd_sc_hd__conb_1
X_10749_ net305 _06322_ _06361_ vssd1 vssd1 vccd1 vccd1 _06362_ sky130_fd_sc_hd__o21ai_1
XFILLER_174_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xteam_08_1446 vssd1 vssd1 vccd1 vccd1 team_08_1446/HI gpio_out[31] sky130_fd_sc_hd__conb_1
XFILLER_118_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xteam_08_1457 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] team_08_1457/LO sky130_fd_sc_hd__conb_1
XANTENNA__09738__S net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16256_ clknet_leaf_30_clk _02466_ net1152 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.toreg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xteam_08_1468 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] team_08_1468/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_93_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13468_ top.CPU.handler.toreg\[23\] _02955_ net120 vssd1 vssd1 vccd1 vccd1 _02489_
+ sky130_fd_sc_hd__mux2_1
XFILLER_127_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12672__B _04955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14941__Q top.CPU.alu.program_counter\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09568__A1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15207_ net1541 _01417_ net1191 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12419_ _06935_ _06942_ _06943_ _06944_ vssd1 vssd1 vccd1 vccd1 _06945_ sky130_fd_sc_hd__or4_4
XFILLER_126_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16187_ net2521 _02397_ net1208 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[987\]
+ sky130_fd_sc_hd__dfrtp_1
X_13399_ top.I2C.data_out\[25\] net555 _02916_ net598 vssd1 vssd1 vccd1 vccd1 _02917_
+ sky130_fd_sc_hd__a22o_1
XFILLER_127_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11375__A1 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07579__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08776__C1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15138_ clknet_leaf_47_clk _01348_ net1137 vssd1 vssd1 vccd1 vccd1 top.I2C.data_out\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11288__B net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13915__85 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 net1554 sky130_fd_sc_hd__inv_2
XANTENNA__13116__A2 net1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08791__A2 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15069_ clknet_leaf_55_clk _00047_ net1135 vssd1 vssd1 vccd1 vccd1 top.I2C.output_state\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10760__X _06373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07960_ top.CPU.registers.data\[760\] net1389 net817 top.CPU.registers.data\[728\]
+ net704 vssd1 vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__a221o_1
XANTENNA__11127__A1 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_4_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08528__C1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09473__S net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07782__A net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07891_ top.CPU.registers.data\[60\] top.CPU.registers.data\[28\] net833 vssd1 vssd1
+ vccd1 vccd1 _03530_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_155_Right_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09630_ _05194_ _05267_ _05193_ vssd1 vssd1 vccd1 vccd1 _05269_ sky130_fd_sc_hd__a21boi_2
XANTENNA__09740__A1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10886__B1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10412__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08089__S net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09561_ top.CPU.registers.data\[640\] net1286 net1004 top.CPU.registers.data\[672\]
+ net903 vssd1 vssd1 vccd1 vccd1 _05200_ sky130_fd_sc_hd__a221o_1
XANTENNA__13824__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08512_ net793 _04143_ _04144_ _04150_ vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__a31o_1
X_09492_ net923 _05128_ _05130_ net622 vssd1 vssd1 vccd1 vccd1 _05131_ sky130_fd_sc_hd__o211a_1
XANTENNA__08700__C1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08443_ top.CPU.registers.data\[561\] top.CPU.registers.data\[529\] net832 vssd1
+ vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__mux2_1
XANTENNA__12339__S net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout151_A _06780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11850__A2 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12566__C _06352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08374_ top.CPU.registers.data\[338\] net1320 net851 top.CPU.registers.data\[370\]
+ net769 vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__a221o_1
XANTENNA__08059__A1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11602__A2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1060_A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1158_A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09008__B1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13355__A2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout204_X net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1325_A net1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08767__C1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08231__A1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10574__C1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout785_A net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1113_X net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout410 net411 vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__buf_2
Xfanout1408 top.CPU.control_unit.instruction\[5\] vssd1 vssd1 vccd1 vccd1 net1408
+ sky130_fd_sc_hd__buf_2
Xfanout421 net423 vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__buf_4
XANTENNA__07990__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout432 _06602_ vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__clkbuf_8
XANTENNA__15633__RESET_B net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout443 _05678_ vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__buf_2
Xfanout454 net455 vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11669__A2 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout573_X net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout952_A net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout465 net467 vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_126_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09731__A1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09192__C1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout476 net477 vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_161_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09828_ top.CPU.alu.program_counter\[26\] _05465_ net1036 vssd1 vssd1 vccd1 vccd1
+ _05467_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_122_Right_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout487 net491 vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout498 net500 vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__clkbuf_8
XFILLER_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14562__732 clknet_leaf_140_clk vssd1 vssd1 vccd1 vccd1 net2201 sky130_fd_sc_hd__inv_2
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09759_ top.CPU.alu.program_counter\[27\] net1037 vssd1 vssd1 vccd1 vccd1 _05398_
+ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout740_X net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13815__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout838_X net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10629__B1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13633__S net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08298__A1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12770_ _07225_ _07226_ vssd1 vssd1 vccd1 vccd1 _07227_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12094__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14603__773 clknet_leaf_135_clk vssd1 vssd1 vccd1 vccd1 net2242 sky130_fd_sc_hd__inv_2
X_11721_ _06563_ net201 net421 net2996 vssd1 vssd1 vccd1 vccd1 _01832_ sky130_fd_sc_hd__a22o_1
XANTENNA__08393__S1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11841__A2 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09247__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11652_ _06293_ net197 net424 net3334 vssd1 vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__a22o_1
XFILLER_168_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10603_ net412 _06220_ _06221_ _06222_ vssd1 vssd1 vccd1 vccd1 _06223_ sky130_fd_sc_hd__a31o_1
X_11583_ _06694_ net259 net246 net2789 vssd1 vssd1 vccd1 vccd1 _01959_ sky130_fd_sc_hd__a22o_1
XFILLER_70_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16110_ net2444 _02320_ net1107 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[910\]
+ sky130_fd_sc_hd__dfrtp_1
X_13322_ net888 _02860_ vssd1 vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__and2_1
XANTENNA__10801__B1 _06411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10534_ net447 _06155_ _06156_ _05571_ vssd1 vssd1 vccd1 vccd1 _06157_ sky130_fd_sc_hd__a22o_1
XANTENNA__12492__B _04792_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16041_ net2375 _02251_ net1055 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[841\]
+ sky130_fd_sc_hd__dfrtp_1
X_10465_ _05899_ _06090_ net403 vssd1 vssd1 vccd1 vccd1 _06091_ sky130_fd_sc_hd__mux2_1
X_13253_ top.I2C.data_out\[9\] net893 _02774_ vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__mux2_1
XANTENNA__07586__B _03200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12204_ net3500 net168 _06869_ vssd1 vssd1 vccd1 vccd1 _01460_ sky130_fd_sc_hd__a21bo_1
X_10396_ net408 _05787_ _06024_ _05664_ vssd1 vssd1 vccd1 vccd1 _06025_ sky130_fd_sc_hd__a211o_1
X_13184_ top.I2C.I2C_state\[20\] top.I2C.I2C_state\[25\] top.I2C.I2C_state\[4\] top.I2C.I2C_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__or4_1
XFILLER_151_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12135_ net4003 net174 _06835_ _06650_ vssd1 vssd1 vccd1 vccd1 _01495_ sky130_fd_sc_hd__a22o_1
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09293__S net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07981__B1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11109__B2 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12066_ top.CPU.registers.data\[120\] net649 _03185_ vssd1 vssd1 vccd1 vccd1 _06802_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__10317__C1 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_8_Left_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09183__C1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08525__A2 net1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11017_ net1406 _03170_ net147 vssd1 vssd1 vccd1 vccd1 _06565_ sky130_fd_sc_hd__or3b_1
XANTENNA__09722__B2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10332__A2 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08930__C1 net1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15825_ net2159 _02035_ net1175 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[625\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_38_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12948__A top.CPU.alu.program_counter\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15756_ net2090 _01966_ net1078 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[556\]
+ sky130_fd_sc_hd__dfrtp_1
X_12968_ _07403_ _07404_ vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__nor2_1
XANTENNA__13282__A1 top.CPU.handler.readout vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12085__A2 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_0_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11293__B1 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11919_ net3809 net184 net341 _06214_ vssd1 vssd1 vccd1 vccd1 _01647_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_47_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15687_ net2021 _01897_ net1200 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[487\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12899_ _07338_ _07343_ net128 vssd1 vssd1 vccd1 vccd1 _07344_ sky130_fd_sc_hd__mux2_1
XFILLER_60_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09238__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09789__A1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12683__A top.CPU.alu.program_counter\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16308_ clknet_leaf_95_clk _02517_ net1260 vssd1 vssd1 vccd1 vccd1 top.CPU.data_out\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08997__C1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08090_ top.CPU.registers.data\[757\] net1391 net827 top.CPU.registers.data\[725\]
+ net775 vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_60_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload20 clknet_leaf_196_clk vssd1 vssd1 vccd1 vccd1 clkload20/Y sky130_fd_sc_hd__inv_6
XANTENNA__10915__B _06230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16239_ clknet_leaf_46_clk _02449_ net1137 vssd1 vssd1 vccd1 vccd1 top.CPU.control_unit.instruction\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload31 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 clkload31/Y sky130_fd_sc_hd__clkinv_8
XFILLER_162_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload42 clknet_leaf_186_clk vssd1 vssd1 vccd1 vccd1 clkload42/Y sky130_fd_sc_hd__inv_8
XFILLER_161_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload53 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 clkload53/Y sky130_fd_sc_hd__inv_8
XFILLER_127_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload64 clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 clkload64/X sky130_fd_sc_hd__clkbuf_4
Xclkload75 clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 clkload75/Y sky130_fd_sc_hd__inv_6
XANTENNA__08213__A1 net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload86 clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 clkload86/Y sky130_fd_sc_hd__bufinv_16
XFILLER_47_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload97 clknet_leaf_76_clk vssd1 vssd1 vccd1 vccd1 clkload97/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__11449__D net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09961__A1 _05399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07567__A3 net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08992_ net783 _04629_ _04630_ net737 vssd1 vssd1 vccd1 vccd1 _04631_ sky130_fd_sc_hd__o211a_1
X_07943_ top.CPU.registers.data\[312\] top.CPU.registers.data\[280\] net820 vssd1
+ vssd1 vccd1 vccd1 _03582_ sky130_fd_sc_hd__mux2_1
XFILLER_130_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14546__716 clknet_leaf_193_clk vssd1 vssd1 vccd1 vccd1 net2185 sky130_fd_sc_hd__inv_2
XANTENNA__09174__C1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout199_A net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08516__A2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09713__A1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07874_ top.CPU.registers.data\[828\] top.CPU.registers.data\[796\] net833 vssd1
+ vssd1 vccd1 vccd1 _03513_ sky130_fd_sc_hd__mux2_1
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07724__B1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11520__A1 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09613_ top.CPU.registers.data\[736\] net1387 net810 top.CPU.registers.data\[704\]
+ net715 vssd1 vssd1 vccd1 vccd1 _05252_ sky130_fd_sc_hd__a221o_1
XANTENNA__08921__C1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_104_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout366_A net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13306__X _02849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09544_ top.CPU.registers.data\[417\] top.CPU.registers.data\[385\] net835 vssd1
+ vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__mux2_1
XFILLER_24_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09477__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12076__A2 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13273__B2 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11284__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09475_ top.CPU.registers.data\[642\] net1324 net855 top.CPU.registers.data\[674\]
+ net723 vssd1 vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__a221o_1
XANTENNA__11823__A2 _06648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout154_X net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1275_A net1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08426_ top.CPU.registers.data\[177\] top.CPU.registers.data\[145\] net825 vssd1
+ vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__mux2_1
XFILLER_51_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11036__B1 _06577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout321_X net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08357_ net694 _03995_ vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout700_A net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout419_X net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload3 clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clkload3/Y sky130_fd_sc_hd__inv_8
XANTENNA__11587__A1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08288_ top.CPU.registers.data\[339\] net1326 net857 top.CPU.registers.data\[371\]
+ net773 vssd1 vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_119_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10825__B _05670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10795__C1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13328__A2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11002__A net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1328_X net1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10250_ net550 _05503_ net505 _05502_ _05883_ vssd1 vssd1 vccd1 vccd1 _05884_ sky130_fd_sc_hd__o221a_1
XANTENNA__15814__RESET_B net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09401__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12000__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout690_X net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout788_X net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13628__S net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07693__Y _03332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10181_ _05814_ _05816_ net393 vssd1 vssd1 vccd1 vccd1 _05817_ sky130_fd_sc_hd__mux2_1
XANTENNA__10562__A2 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1205 net1233 vssd1 vssd1 vccd1 vccd1 net1205 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07963__B1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_858 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1216 net1217 vssd1 vssd1 vccd1 vccd1 net1216 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1227 net1229 vssd1 vssd1 vccd1 vccd1 net1227 sky130_fd_sc_hd__clkbuf_4
Xfanout1238 net1240 vssd1 vssd1 vccd1 vccd1 net1238 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout955_X net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout240 net242 vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__clkbuf_4
Xfanout1249 net1259 vssd1 vssd1 vccd1 vccd1 net1249 sky130_fd_sc_hd__clkbuf_2
Xfanout251 _06733_ vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__clkbuf_4
X_14289__459 clknet_leaf_180_clk vssd1 vssd1 vccd1 vccd1 net1928 sky130_fd_sc_hd__inv_2
Xfanout262 _06725_ vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__buf_4
XANTENNA__09165__C1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08507__A2 net1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout273 net274 vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__buf_4
Xfanout284 _06713_ vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__clkbuf_8
Xfanout295 _06662_ vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__buf_6
XANTENNA__09180__A2 net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15610_ net1944 _01820_ net1251 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[410\]
+ sky130_fd_sc_hd__dfrtp_1
X_12822_ top.CPU.alu.program_counter\[18\] _07270_ vssd1 vssd1 vccd1 vccd1 _07274_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__09468__B1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15541_ net1875 _01751_ net1227 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[341\]
+ sky130_fd_sc_hd__dfrtp_1
X_12753_ net125 _07207_ _03118_ vssd1 vssd1 vccd1 vccd1 _07212_ sky130_fd_sc_hd__a21oi_1
X_11704_ _06536_ net205 net422 net2929 vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__a22o_1
XFILLER_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15472_ net1806 _01682_ net1107 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[272\]
+ sky130_fd_sc_hd__dfrtp_1
X_12684_ _07147_ _07148_ vssd1 vssd1 vccd1 vccd1 _07149_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_139_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11635_ _05908_ net210 net427 net3431 vssd1 vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__a22o_1
XANTENNA__12775__A0 top.CPU.alu.program_counter\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11578__B2 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11611__S net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14690__860 clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 net2329 sky130_fd_sc_hd__inv_2
X_11566_ _06677_ net262 net247 net2725 vssd1 vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__a22o_1
XFILLER_11_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10250__A1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13305_ net598 _02844_ net554 top.I2C.data_out\[0\] vssd1 vssd1 vccd1 vccd1 _02848_
+ sky130_fd_sc_hd__a22o_1
X_10517_ net415 _06139_ vssd1 vssd1 vccd1 vccd1 _06141_ sky130_fd_sc_hd__nor2_2
X_11497_ net562 _06630_ net254 net3454 vssd1 vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__a22o_1
XFILLER_143_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16024_ net2358 _02234_ net1108 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[824\]
+ sky130_fd_sc_hd__dfrtp_1
X_13236_ net2799 _02776_ _02801_ vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__mux2_1
X_10448_ _03986_ net506 _05733_ _05871_ vssd1 vssd1 vccd1 vccd1 _06075_ sky130_fd_sc_hd__a22o_1
XANTENNA__08920__S net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14233__403 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 net1872 sky130_fd_sc_hd__inv_2
XANTENNA__10173__D _05808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10751__A net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12542__A3 _06450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13167_ top.I2C.within_byte_counter_reading\[1\] top.I2C.within_byte_counter_reading\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__or2_1
X_10379_ top.CPU.fetch.current_ra\[22\] net1041 net881 top.CPU.handler.toreg\[22\]
+ vssd1 vssd1 vccd1 vccd1 _06009_ sky130_fd_sc_hd__a22o_1
XANTENNA__11750__A1 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10553__A2 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09317__A _04955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12118_ top.CPU.registers.data\[93\] net173 vssd1 vssd1 vccd1 vccd1 _06827_ sky130_fd_sc_hd__and2_1
X_13098_ top.SPI.state\[5\] _07426_ vssd1 vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__nor2_1
XANTENNA__08221__A top.CPU.alu.program_counter\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12049_ net568 _06596_ net364 _06780_ top.CPU.registers.data\[129\] vssd1 vssd1 vccd1
+ vccd1 _06794_ sky130_fd_sc_hd__a32o_1
XANTENNA__07706__B1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08903__C1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15808_ net2142 _02018_ net1091 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[608\]
+ sky130_fd_sc_hd__dfrtp_1
X_07590_ top.CPU.registers.data\[511\] net1334 net865 top.CPU.registers.data\[479\]
+ net756 vssd1 vssd1 vccd1 vccd1 _03229_ sky130_fd_sc_hd__o221a_1
XANTENNA__09459__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15739_ net2073 _01949_ net1216 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[539\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_max_cap586_X net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09987__A _04829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09260_ top.CPU.registers.data\[965\] net1286 net1004 top.CPU.registers.data\[997\]
+ net900 vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_62_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08682__A1 net1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08211_ top.CPU.registers.data\[471\] net1295 net1014 top.CPU.registers.data\[503\]
+ net912 vssd1 vssd1 vccd1 vccd1 _03850_ sky130_fd_sc_hd__a221o_1
XFILLER_60_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09191_ top.CPU.registers.data\[294\] top.CPU.registers.data\[262\] net977 vssd1
+ vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__mux2_1
XANTENNA__07890__C1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11569__B2 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09198__S net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08142_ net627 _03779_ _03780_ net606 vssd1 vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__a31o_1
XANTENNA__08434__A1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12230__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload120 clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 clkload120/Y sky130_fd_sc_hd__inv_6
X_08073_ top.CPU.registers.data\[340\] net1288 net1008 top.CPU.registers.data\[372\]
+ net931 vssd1 vssd1 vccd1 vccd1 _03712_ sky130_fd_sc_hd__a221o_1
XFILLER_174_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload131 clknet_leaf_174_clk vssd1 vssd1 vccd1 vccd1 clkload131/Y sky130_fd_sc_hd__clkinv_8
XFILLER_162_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16613__A net1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload142 clknet_leaf_150_clk vssd1 vssd1 vccd1 vccd1 clkload142/Y sky130_fd_sc_hd__inv_2
Xclkload153 clknet_leaf_135_clk vssd1 vssd1 vccd1 vccd1 clkload153/Y sky130_fd_sc_hd__inv_8
Xclkload164 clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 clkload164/Y sky130_fd_sc_hd__inv_4
XFILLER_106_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload175 clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 clkload175/Y sky130_fd_sc_hd__inv_6
XFILLER_162_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload186 clknet_leaf_87_clk vssd1 vssd1 vccd1 vccd1 clkload186/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__13448__S net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09395__C1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1023_A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11476__B net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08975_ top.CPU.registers.data\[41\] top.CPU.registers.data\[9\] net806 vssd1 vssd1
+ vccd1 vccd1 _04614_ sky130_fd_sc_hd__mux2_1
XANTENNA__08131__A net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout483_A net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold15 top.CPU.registers.data_out_r2_prev\[7\] vssd1 vssd1 vccd1 vccd1 net2572 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09147__C1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold26 top.CPU.registers.data_out_r1_prev\[20\] vssd1 vssd1 vccd1 vccd1 net2583 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 top.I2C.I2C_state\[19\] vssd1 vssd1 vccd1 vccd1 net2594 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07926_ net683 _03560_ _03561_ _03564_ net614 vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__a311o_1
Xhold48 top.CPU.registers.data_out_r2_prev\[26\] vssd1 vssd1 vccd1 vccd1 net2605 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_60_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14017__187 clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 net1656 sky130_fd_sc_hd__inv_2
Xhold59 _00039_ vssd1 vssd1 vccd1 vccd1 net2616 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09698__B1 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout650_A net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07857_ top.CPU.registers.data\[925\] net1289 net1007 top.CPU.registers.data\[957\]
+ net906 vssd1 vssd1 vccd1 vccd1 _03496_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout271_X net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout748_A net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout369_X net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1392_A net1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08370__B1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13246__B2 _02803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07788_ top.CPU.registers.data\[862\] net1302 net1023 top.CPU.registers.data\[894\]
+ net944 vssd1 vssd1 vccd1 vccd1 _03427_ sky130_fd_sc_hd__a221o_1
X_09527_ net780 _05161_ _05162_ _05165_ vssd1 vssd1 vccd1 vccd1 _05166_ sky130_fd_sc_hd__a31o_1
XANTENNA__12875__X _07322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout915_A net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout536_X net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09458_ top.CPU.registers.data\[418\] top.CPU.registers.data\[386\] net823 vssd1
+ vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_156_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14674__844 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 net2313 sky130_fd_sc_hd__inv_2
X_08409_ net675 _04041_ _04047_ _04027_ _04035_ vssd1 vssd1 vccd1 vccd1 _04048_ sky130_fd_sc_hd__a32o_4
XFILLER_101_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07881__C1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09389_ top.CPU.registers.data\[67\] net1328 net859 top.CPU.registers.data\[99\]
+ net775 vssd1 vssd1 vccd1 vccd1 _05028_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout703_X net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11420_ _06558_ net275 net267 net2747 vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__a22o_1
XFILLER_138_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12221__A2 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08976__A2 net1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11351_ net3783 net285 net275 _06255_ vssd1 vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__a22o_1
X_14715__885 clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 net2354 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_134_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12509__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_747 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10302_ _05933_ net575 net521 vssd1 vssd1 vccd1 vccd1 _05935_ sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_89_Left_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11282_ net2948 net296 _06698_ net320 vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__a22o_1
XFILLER_152_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08189__B1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13021_ top.SPI.parameters\[12\] top.SPI.paroutput\[4\] net1355 vssd1 vssd1 vccd1
+ vccd1 _07436_ sky130_fd_sc_hd__mux2_1
XFILLER_4_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10233_ _05642_ _05865_ _05867_ _05863_ vssd1 vssd1 vccd1 vccd1 _05868_ sky130_fd_sc_hd__a31o_1
XFILLER_152_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12262__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10571__A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10164_ _05795_ _05800_ net390 vssd1 vssd1 vccd1 vccd1 _05801_ sky130_fd_sc_hd__mux2_1
Xfanout1002 net1003 vssd1 vssd1 vccd1 vccd1 net1002 sky130_fd_sc_hd__buf_2
XFILLER_79_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1013 net1032 vssd1 vssd1 vccd1 vccd1 net1013 sky130_fd_sc_hd__clkbuf_2
XFILLER_117_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1024 net1031 vssd1 vssd1 vccd1 vccd1 net1024 sky130_fd_sc_hd__clkbuf_2
Xfanout1035 net1036 vssd1 vssd1 vccd1 vccd1 net1035 sky130_fd_sc_hd__clkbuf_4
Xfanout1046 _03156_ vssd1 vssd1 vccd1 vccd1 net1046 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10095_ net403 _05643_ vssd1 vssd1 vccd1 vccd1 _05733_ sky130_fd_sc_hd__nor2_2
X_14972_ clknet_leaf_93_clk _01217_ net1268 vssd1 vssd1 vccd1 vccd1 top.SPI.paroutput\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1057 net1059 vssd1 vssd1 vccd1 vccd1 net1057 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1068 net1111 vssd1 vssd1 vccd1 vccd1 net1068 sky130_fd_sc_hd__buf_2
Xfanout1079 net1111 vssd1 vssd1 vccd1 vccd1 net1079 sky130_fd_sc_hd__buf_2
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11496__B1 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11606__S net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08361__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10510__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_98_Left_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12805_ _07257_ _07258_ vssd1 vssd1 vccd1 vccd1 _07259_ sky130_fd_sc_hd__nor2_1
XANTENNA__13788__A2 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13785_ net14 net1050 net885 net3922 vssd1 vssd1 vccd1 vccd1 _02666_ sky130_fd_sc_hd__o22a_1
XFILLER_76_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10997_ net3397 net217 _06552_ net313 vssd1 vssd1 vccd1 vccd1 _02350_ sky130_fd_sc_hd__a22o_1
XFILLER_163_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15524_ net1858 _01734_ net1186 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[324\]
+ sky130_fd_sc_hd__dfrtp_1
X_12736_ _07194_ _07195_ vssd1 vssd1 vccd1 vccd1 _07196_ sky130_fd_sc_hd__nand2_1
XFILLER_37_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09861__A0 _05498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10471__A1 _05733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15455_ net1789 _01665_ net1220 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[255\]
+ sky130_fd_sc_hd__dfrtp_1
X_12667_ _07132_ _07133_ vssd1 vssd1 vccd1 vccd1 _07134_ sky130_fd_sc_hd__xor2_1
X_11618_ net144 net3583 net212 vssd1 vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__mux2_1
XANTENNA__09613__B1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12212__A2 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15386_ net1720 _01596_ net1251 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[186\]
+ sky130_fd_sc_hd__dfrtp_1
X_12598_ top.SPI.count\[2\] _03141_ top.SPI.count\[1\] _03142_ _07098_ vssd1 vssd1
+ vccd1 vccd1 _07099_ sky130_fd_sc_hd__a221o_1
XFILLER_128_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10223__A1 _05399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11420__B1 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11549_ _06663_ net282 net248 net2875 vssd1 vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__a22o_1
Xhold507 top.SPI.parameters\[7\] vssd1 vssd1 vccd1 vccd1 net3064 sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 top.CPU.registers.data\[185\] vssd1 vssd1 vccd1 vccd1 net3075 sky130_fd_sc_hd__dlygate4sd3_1
Xhold529 top.CPU.registers.data\[821\] vssd1 vssd1 vccd1 vccd1 net3086 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13268__S _02780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16007_ net2341 _02217_ net1203 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[807\]
+ sky130_fd_sc_hd__dfrtp_1
X_13219_ top.I2C.output_state\[28\] _02791_ vssd1 vssd1 vccd1 vccd1 _02792_ sky130_fd_sc_hd__and2_1
XANTENNA__11577__A net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10481__A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07927__B1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1207 top.CPU.registers.data\[53\] vssd1 vssd1 vccd1 vccd1 net3764 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12900__S net1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08760_ top.CPU.registers.data\[684\] top.CPU.registers.data\[652\] net815 vssd1
+ vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__mux2_1
XANTENNA__12279__A2 _06887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1218 top.CPU.registers.data_out_r1_prev\[28\] vssd1 vssd1 vccd1 vccd1 net3775
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1229 top.SPI.timem\[15\] vssd1 vssd1 vccd1 vccd1 net3786 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09144__A2 net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07711_ top.CPU.registers.data\[63\] top.CPU.registers.data\[31\] net999 vssd1 vssd1
+ vccd1 vccd1 _03350_ sky130_fd_sc_hd__mux2_1
XANTENNA__11487__B1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08691_ _04327_ _04329_ vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__nand2_2
XFILLER_54_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_201_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_201_clk
+ sky130_fd_sc_hd__clkbuf_8
X_07642_ net1400 _03108_ _03279_ vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__a21oi_1
XFILLER_38_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14361__531 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 net2000 sky130_fd_sc_hd__inv_2
X_07573_ net1048 _03164_ net1039 top.CPU.control_unit.instruction\[18\] vssd1 vssd1
+ vccd1 vccd1 _03212_ sky130_fd_sc_hd__o31a_4
XTAP_TAPCELL_ROW_24_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14658__828 clknet_leaf_143_clk vssd1 vssd1 vccd1 vccd1 net2297 sky130_fd_sc_hd__inv_2
X_09312_ _04944_ _04950_ vssd1 vssd1 vccd1 vccd1 _04951_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_24_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08825__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09852__B1 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09243_ top.CPU.registers.data\[69\] net1310 net841 top.CPU.registers.data\[101\]
+ net737 vssd1 vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__a221o_1
XFILLER_90_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14402__572 clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 net2041 sky130_fd_sc_hd__inv_2
XANTENNA_fanout231_A _06772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout329_A _03096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12574__C _06054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08407__A1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09174_ _03111_ _04812_ _04805_ net639 vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__a211o_1
XANTENNA__09604__B1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08125_ top.CPU.registers.data\[181\] top.CPU.registers.data\[149\] net993 vssd1
+ vssd1 vccd1 vccd1 _03764_ sky130_fd_sc_hd__mux2_1
XANTENNA__15406__RESET_B net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11411__B1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1140_A net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12871__A top.CPU.alu.program_counter\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11962__A1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08056_ top.CPU.registers.data\[596\] net1288 net1008 top.CPU.registers.data\[628\]
+ net931 vssd1 vssd1 vccd1 vccd1 _03695_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_112_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout698_A net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput49 net49 vssd1 vssd1 vccd1 vccd1 ADR_O[19] sky130_fd_sc_hd__buf_2
XFILLER_163_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12911__A0 top.CPU.alu.program_counter\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1405_A net1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1026_X net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout486_X net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout865_A net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07971__Y _03610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12810__S net1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08958_ net1363 _03150_ net1042 _03177_ vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__or4_2
XANTENNA__13467__A1 net1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13876__46 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 net1515 sky130_fd_sc_hd__inv_2
XFILLER_130_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11478__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07909_ top.CPU.registers.data\[156\] net996 _03547_ vssd1 vssd1 vccd1 vccd1 _03548_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__11934__B net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08889_ net738 _04509_ _04510_ _04513_ net703 vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__a311o_1
XANTENNA_fanout653_X net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1395_X net1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10920_ net480 net457 _06505_ net220 net3011 vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__a32o_1
XANTENNA__07697__A2 _03262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10851_ net394 _06379_ _06458_ net409 vssd1 vssd1 vccd1 vccd1 _06459_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout820_X net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout918_X net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13641__S net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13570_ top.CPU.addressnew\[8\] net578 _03007_ _03008_ vssd1 vssd1 vccd1 vccd1 _02538_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_160_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08646__A1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09843__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10782_ net3651 net226 net318 _06393_ vssd1 vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__a22o_1
XFILLER_24_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12521_ _06968_ _06993_ _07029_ vssd1 vssd1 vccd1 vccd1 _07030_ sky130_fd_sc_hd__or3_1
XANTENNA__11650__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07854__C1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_40_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12257__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15240_ net1574 _01450_ net1065 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[40\]
+ sky130_fd_sc_hd__dfrtp_1
X_12452_ net898 _06961_ vssd1 vssd1 vccd1 vccd1 _00045_ sky130_fd_sc_hd__nor2_1
XFILLER_157_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_175_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11403_ _06533_ net282 net270 net3799 vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__a22o_1
XANTENNA__10205__B2 _05733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11402__B1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15171_ net1508 _01381_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r1_prev\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_12383_ top.CPU.addressnew\[3\] top.CPU.addressnew\[18\] top.CPU.addressnew\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06921_ sky130_fd_sc_hd__and3b_1
XFILLER_153_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10853__X _06461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13596__B net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11334_ net3615 net288 net283 _05849_ vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_55_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09359__C1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11397__A net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07594__B net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11265_ net3049 net293 _06689_ net478 vssd1 vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__a22o_1
XFILLER_134_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13004_ net1358 _07428_ vssd1 vssd1 vccd1 vccd1 _07431_ sky130_fd_sc_hd__nor2_4
X_10216_ _05502_ _05850_ vssd1 vssd1 vccd1 vccd1 _05851_ sky130_fd_sc_hd__nand2_1
XANTENNA__08031__C1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11196_ _06231_ net3645 net297 vssd1 vssd1 vccd1 vccd1 _02254_ sky130_fd_sc_hd__mux2_1
XANTENNA__12005__B _06779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08582__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10147_ _03407_ _03476_ net374 vssd1 vssd1 vccd1 vccd1 _05784_ sky130_fd_sc_hd__mux2_1
XANTENNA__12720__S net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09154__X _04793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11469__A0 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09126__A2 _04763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_113_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14955_ clknet_leaf_53_clk _01201_ net1133 vssd1 vssd1 vccd1 vccd1 top.I2C.bit_timer_counter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10078_ _05714_ _05715_ vssd1 vssd1 vccd1 vccd1 _05716_ sky130_fd_sc_hd__nor2_1
X_14345__515 clknet_leaf_155_clk vssd1 vssd1 vccd1 vccd1 net1984 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_50_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12681__A2 _03118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16625_ top.SPI.csx vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__clkbuf_1
X_13890__60 clknet_leaf_140_clk vssd1 vssd1 vccd1 vccd1 net1529 sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_128_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08098__C1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13768_ net27 net1051 net886 net3995 vssd1 vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__a22o_1
XANTENNA__13630__A1 _03100_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09834__B1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14944__Q top.CPU.alu.program_counter\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12719_ _07178_ _07180_ vssd1 vssd1 vccd1 vccd1 _07181_ sky130_fd_sc_hd__xor2_1
X_15507_ net1841 _01717_ net1191 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[307\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11641__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16487_ clknet_leaf_41_clk _02649_ net1115 vssd1 vssd1 vccd1 vccd1 top.mmio.mem_data_i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_13699_ top.SPI.timem\[3\] top.SPI.timem\[2\] _03052_ vssd1 vssd1 vccd1 vccd1 _03054_
+ sky130_fd_sc_hd__and3_1
XFILLER_87_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10995__A2 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15438_ net1772 _01648_ net1105 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[238\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07860__A2 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13394__A0 top.CPU.control_unit.instruction\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_157_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09598__C1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15369_ net1703 _01579_ net1061 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[169\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_144_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09476__S net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold304 net78 vssd1 vssd1 vccd1 vccd1 net2861 sky130_fd_sc_hd__dlygate4sd3_1
Xhold315 top.CPU.registers.data\[854\] vssd1 vssd1 vccd1 vccd1 net2872 sky130_fd_sc_hd__dlygate4sd3_1
Xhold326 _01266_ vssd1 vssd1 vccd1 vccd1 net2883 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold337 net82 vssd1 vssd1 vccd1 vccd1 net2894 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold348 top.CPU.registers.data\[287\] vssd1 vssd1 vccd1 vccd1 net2905 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09930_ _05537_ _05564_ _05566_ _05540_ vssd1 vssd1 vccd1 vccd1 _05569_ sky130_fd_sc_hd__a31o_1
XFILLER_116_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold359 top.CPU.registers.data\[621\] vssd1 vssd1 vccd1 vccd1 net2916 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11100__A net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09365__A2 net1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout806 net813 vssd1 vssd1 vccd1 vccd1 net806 sky130_fd_sc_hd__clkbuf_4
X_09861_ _05498_ _05499_ net455 vssd1 vssd1 vccd1 vccd1 _05500_ sky130_fd_sc_hd__mux2_1
XANTENNA__08022__C1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout817 net822 vssd1 vssd1 vccd1 vccd1 net817 sky130_fd_sc_hd__clkbuf_4
Xfanout828 net831 vssd1 vssd1 vccd1 vccd1 net828 sky130_fd_sc_hd__buf_4
XFILLER_97_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08573__B1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11172__A2 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout839 _03204_ vssd1 vssd1 vccd1 vccd1 net839 sky130_fd_sc_hd__clkbuf_4
X_13953__123 clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 net1592 sky130_fd_sc_hd__inv_2
XANTENNA__09770__C1 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08812_ top.CPU.registers.data\[684\] net1292 vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__or2_1
XFILLER_140_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09792_ _05430_ vssd1 vssd1 vccd1 vccd1 _05431_ sky130_fd_sc_hd__inv_2
XANTENNA__13449__A1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1004 top.CPU.registers.data\[225\] vssd1 vssd1 vccd1 vccd1 net3561 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1015 top.CPU.registers.data\[841\] vssd1 vssd1 vccd1 vccd1 net3572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1026 top.CPU.registers.data\[521\] vssd1 vssd1 vccd1 vccd1 net3583 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09117__A2 net1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08743_ top.CPU.registers.data\[685\] top.CPU.registers.data\[653\] top.CPU.registers.data\[557\]
+ top.CPU.registers.data\[525\] net970 net901 vssd1 vssd1 vccd1 vccd1 _04382_ sky130_fd_sc_hd__mux4_1
Xhold1037 top.CPU.registers.data\[948\] vssd1 vssd1 vccd1 vccd1 net3594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1048 top.CPU.registers.data\[1013\] vssd1 vssd1 vccd1 vccd1 net3605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1059 top.I2C.bit_timer_state\[1\] vssd1 vssd1 vccd1 vccd1 net3616 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout181_A _06777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08325__B1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout279_A _06713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11473__C net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08674_ top.CPU.registers.data\[942\] top.CPU.registers.data\[910\] top.CPU.registers.data\[814\]
+ top.CPU.registers.data\[782\] net985 net1282 vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__mux4_1
X_14088__258 clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 net1727 sky130_fd_sc_hd__inv_2
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07625_ top.CPU.control_unit.instruction\[26\] top.CPU.control_unit.instruction\[25\]
+ top.CPU.control_unit.instruction\[30\] _03257_ vssd1 vssd1 vccd1 vccd1 _03264_ sky130_fd_sc_hd__or4_2
XANTENNA__11880__A0 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1188_A net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07556_ _03189_ net471 vssd1 vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__nor2_1
XANTENNA__13621__A1 _05806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12585__B net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14129__299 clknet_leaf_190_clk vssd1 vssd1 vccd1 vccd1 net1768 sky130_fd_sc_hd__inv_2
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_153_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11632__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07487_ top.SPI.register\[1\] vssd1 vssd1 vccd1 vccd1 _03127_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_153_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout234_X net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout613_A net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1355_A top.SPI.state\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09226_ net702 _04863_ _04864_ vssd1 vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_170_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09894__B _04567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09157_ _04765_ _04794_ vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout401_X net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10673__X _06290_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11935__A1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09386__S net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08108_ top.CPU.registers.data\[821\] top.CPU.registers.data\[789\] net830 vssd1
+ vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__mux2_1
XANTENNA__08261__C1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09088_ net689 _04726_ _04699_ vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__o21ai_2
XPHY_EDGE_ROW_169_Right_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout982_A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08039_ net746 _03676_ _03677_ net704 vssd1 vssd1 vccd1 vccd1 _03678_ sky130_fd_sc_hd__o211a_1
X_14786__956 clknet_leaf_143_clk vssd1 vssd1 vccd1 vccd1 net2425 sky130_fd_sc_hd__inv_2
XFILLER_174_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold860 top.CPU.registers.data\[524\] vssd1 vssd1 vccd1 vccd1 net3417 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_107_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10552__C net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11010__A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold871 top.CPU.registers.data\[408\] vssd1 vssd1 vccd1 vccd1 net3428 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16446__RESET_B net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold882 _01210_ vssd1 vssd1 vccd1 vccd1 net3439 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold893 top.SPI.timem\[2\] vssd1 vssd1 vccd1 vccd1 net3450 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09356__A2 net1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11050_ net3565 net368 _06583_ net325 vssd1 vssd1 vccd1 vccd1 _02328_ sky130_fd_sc_hd__a22o_1
XANTENNA__11699__B1 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout770_X net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08564__B1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout868_X net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10001_ _05636_ _05639_ net387 vssd1 vssd1 vccd1 vccd1 _05640_ sky130_fd_sc_hd__mux2_1
XANTENNA__13636__S net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14032__202 clknet_leaf_196_clk vssd1 vssd1 vccd1 vccd1 net1671 sky130_fd_sc_hd__inv_2
X_14827__997 clknet_leaf_164_clk vssd1 vssd1 vccd1 vccd1 net2466 sky130_fd_sc_hd__inv_2
XFILLER_88_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_129_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11952_ _06496_ net343 net229 net3433 vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__a22o_1
XFILLER_85_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10903_ net146 net436 vssd1 vssd1 vccd1 vccd1 _06495_ sky130_fd_sc_hd__and2_1
XANTENNA__11871__B1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11883_ _06709_ net240 net189 net3781 vssd1 vssd1 vccd1 vccd1 _01680_ sky130_fd_sc_hd__a22o_1
XANTENNA__12776__A top.CPU.alu.program_counter\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16410_ clknet_leaf_56_clk net2621 net1142 vssd1 vssd1 vccd1 vccd1 top.I2C.I2C_state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13622_ net2800 _03039_ net581 vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__mux2_1
X_10834_ net397 _06279_ _06280_ net406 vssd1 vssd1 vccd1 vccd1 _06443_ sky130_fd_sc_hd__o211ai_1
XANTENNA__09816__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12495__B _05120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10426__A1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16341_ clknet_leaf_74_clk _02550_ net1159 vssd1 vssd1 vccd1 vccd1 top.CPU.addressnew\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11623__A0 _06391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13553_ net1350 _06426_ vssd1 vssd1 vccd1 vccd1 _02998_ sky130_fd_sc_hd__nand2_1
XANTENNA__07827__C1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10765_ _05272_ net446 _06376_ vssd1 vssd1 vccd1 vccd1 _06377_ sky130_fd_sc_hd__and3b_1
XANTENNA__08095__A2 net1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10977__A2 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12504_ _07001_ _07011_ vssd1 vssd1 vccd1 vccd1 _07013_ sky130_fd_sc_hd__nand2_1
X_16272_ clknet_leaf_60_clk _02482_ net1138 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.toreg\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13484_ net3173 _02963_ net124 vssd1 vssd1 vccd1 vccd1 _02497_ sky130_fd_sc_hd__mux2_1
XANTENNA__07842__A2 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10696_ net438 _06311_ vssd1 vssd1 vccd1 vccd1 _06312_ sky130_fd_sc_hd__and2_1
XANTENNA__13376__A0 top.CPU.control_unit.instruction\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_9_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15223_ net1557 _01433_ net1184 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_172_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12435_ net1339 top.I2C.output_state\[9\] top.I2C.output_state\[23\] vssd1 vssd1
+ vccd1 vccd1 _06954_ sky130_fd_sc_hd__a21o_1
XFILLER_126_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14730__900 clknet_leaf_151_clk vssd1 vssd1 vccd1 vccd1 net2369 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13400__A net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15154_ clknet_leaf_42_clk _01364_ net1118 vssd1 vssd1 vccd1 vccd1 top.I2C.data_out\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_39_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12366_ top.I2C.output_state\[14\] top.I2C.output_state\[7\] top.I2C.output_state\[26\]
+ top.I2C.output_state\[20\] vssd1 vssd1 vccd1 vccd1 _06907_ sky130_fd_sc_hd__or4_1
XFILLER_148_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08252__C1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_136_Right_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11317_ net3527 net289 net357 net144 vssd1 vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__a22o_1
X_15085_ clknet_leaf_64_clk _00041_ net1145 vssd1 vssd1 vccd1 vccd1 top.I2C.byte_manager_state\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_91_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12297_ net2581 _06887_ vssd1 vssd1 vccd1 vccd1 _06890_ sky130_fd_sc_hd__nand2_1
XANTENNA__11558__C net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13937__107 clknet_leaf_180_clk vssd1 vssd1 vccd1 vccd1 net1576 sky130_fd_sc_hd__inv_2
X_11248_ net513 _06174_ net540 vssd1 vssd1 vccd1 vccd1 _06679_ sky130_fd_sc_hd__or3_1
XFILLER_79_130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09752__C1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11179_ net133 net3577 net299 vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__mux2_1
XFILLER_121_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14939__Q top.CPU.alu.program_counter\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15987_ net2321 _02197_ net1197 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[787\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09504__C1 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14938_ clknet_leaf_75_clk _01184_ net1159 vssd1 vssd1 vccd1 vccd1 top.CPU.alu.program_counter\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10665__A1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09979__B _05616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11862__B1 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10758__X _06371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11590__A net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08390_ net934 _04028_ vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__or2_1
XANTENNA__11614__A0 _06212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16539_ clknet_leaf_99_clk _02701_ net1256 vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10968__A2 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09995__A _04698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09011_ net1283 _04646_ _04649_ net617 vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__a211o_1
XFILLER_12_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14473__643 clknet_leaf_154_clk vssd1 vssd1 vccd1 vccd1 net2112 sky130_fd_sc_hd__inv_2
XANTENNA__10934__A net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13310__A _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold101 top.CPU.registers.data\[814\] vssd1 vssd1 vccd1 vccd1 net2658 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09130__S1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold112 top.SPI.parameters\[1\] vssd1 vssd1 vccd1 vccd1 net2669 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 net113 vssd1 vssd1 vccd1 vccd1 net2680 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10653__B net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11393__A2 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold134 top.CPU.registers.data\[908\] vssd1 vssd1 vccd1 vccd1 net2691 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_103_Right_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold145 top.SPI.parameters\[2\] vssd1 vssd1 vccd1 vccd1 net2702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 top.SPI.parameters\[9\] vssd1 vssd1 vccd1 vccd1 net2713 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 top.CPU.registers.data\[318\] vssd1 vssd1 vccd1 vccd1 net2724 sky130_fd_sc_hd__dlygate4sd3_1
X_14514__684 clknet_leaf_201_clk vssd1 vssd1 vccd1 vccd1 net2153 sky130_fd_sc_hd__inv_2
Xhold178 _01200_ vssd1 vssd1 vccd1 vccd1 net2735 sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ net386 _05123_ vssd1 vssd1 vccd1 vccd1 _05552_ sky130_fd_sc_hd__and2_1
Xfanout603 _05689_ vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__clkbuf_4
Xhold189 top.SPI.paroutput\[15\] vssd1 vssd1 vccd1 vccd1 net2746 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout614 net615 vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__buf_4
Xfanout625 net626 vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__buf_4
XANTENNA__13456__S net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09743__C1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout636 net639 vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__clkbuf_8
Xfanout647 net650 vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__clkbuf_4
X_09844_ top.CPU.registers.data\[858\] net1306 net1027 top.CPU.registers.data\[890\]
+ net945 vssd1 vssd1 vccd1 vccd1 _05483_ sky130_fd_sc_hd__a221o_1
XANTENNA__08410__Y _04049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1103_A net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout669 _00000_ vssd1 vssd1 vccd1 vccd1 net669 sky130_fd_sc_hd__buf_2
XFILLER_58_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_146_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13846__16 clknet_leaf_76_clk vssd1 vssd1 vccd1 vccd1 net1485 sky130_fd_sc_hd__inv_2
XFILLER_37_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09775_ net679 _05412_ _05413_ vssd1 vssd1 vccd1 vccd1 _05414_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout563_A net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout184_X net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10105__A0 _05332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08726_ top.CPU.registers.data_out_r2_prev\[13\] net689 vssd1 vssd1 vccd1 vccd1 _04365_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_107_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09510__A2 net1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11853__B1 net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08657_ top.CPU.registers.data_out_r2_prev\[14\] net689 vssd1 vssd1 vccd1 vccd1 _04296_
+ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout351_X net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout730_A net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout828_A net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07608_ _03107_ net1397 net1400 vssd1 vssd1 vccd1 vccd1 _03247_ sky130_fd_sc_hd__a21oi_1
XFILLER_41_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08588_ top.CPU.registers.data_out_r2_prev\[15\] net689 vssd1 vssd1 vccd1 vccd1 _04227_
+ sky130_fd_sc_hd__nand2_1
XFILLER_53_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07539_ net1408 top.CPU.control_unit.instruction\[6\] net1278 vssd1 vssd1 vccd1 vccd1
+ _03178_ sky130_fd_sc_hd__or3_1
XANTENNA__11605__B1 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07809__C1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout616_X net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10959__A2 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11005__A net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10550_ net602 _06171_ _06172_ vssd1 vssd1 vccd1 vccd1 _06173_ sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_33_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13358__A0 net1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11620__A3 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12558__D_N _05958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09209_ net618 _04845_ _04846_ _04847_ vssd1 vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__a31o_1
X_10481_ net527 _06106_ vssd1 vssd1 vccd1 vccd1 _06107_ sky130_fd_sc_hd__nor2_1
XFILLER_136_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13220__A top.I2C.output_state\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12220_ _06746_ net234 net168 net2736 vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__a22o_1
XANTENNA__12030__A0 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08234__C1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout985_X net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11384__A2 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12151_ net3934 net172 _06843_ _06655_ vssd1 vssd1 vccd1 vccd1 _01487_ sky130_fd_sc_hd__a22o_1
XFILLER_118_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11102_ net1406 net577 net529 net136 vssd1 vssd1 vccd1 vccd1 _06609_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_34_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12082_ net3946 net650 _06809_ vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__o21a_1
Xhold690 top.CPU.registers.data\[20\] vssd1 vssd1 vccd1 vccd1 net3247 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_34_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12333__A1 _04792_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13530__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09734__C1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11033_ net1401 net479 net534 vssd1 vssd1 vccd1 vccd1 _06576_ sky130_fd_sc_hd__nand3_1
X_15910_ net2244 _02120_ net1072 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[710\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10344__A0 _03613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12270__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08001__A2 net1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11687__A3 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15841_ net2175 _02051_ net1231 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[641\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12097__B1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12984_ _07415_ top.I2C.bit_timer_state\[0\] _07413_ vssd1 vssd1 vccd1 vccd1 _01201_
+ sky130_fd_sc_hd__and3b_1
XFILLER_18_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15772_ net2106 _01982_ net1236 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[572\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_91_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1390 top.CPU.registers.data\[83\] vssd1 vssd1 vccd1 vccd1 net3947 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09501__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10647__B2 _05672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11844__B1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11935_ net520 _06473_ net351 _06773_ vssd1 vssd1 vccd1 vccd1 _01633_ sky130_fd_sc_hd__a31o_1
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09799__B net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11614__S net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13860__30 clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 net1499 sky130_fd_sc_hd__inv_2
XFILLER_60_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08195__S net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11866_ _05771_ net3481 net190 vssd1 vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__mux2_1
X_13605_ top.CPU.alu.program_counter\[22\] _06008_ net1348 vssd1 vssd1 vccd1 vccd1
+ _03030_ sky130_fd_sc_hd__mux2_1
X_10817_ net600 _06426_ vssd1 vssd1 vccd1 vccd1 _06427_ sky130_fd_sc_hd__nor2_1
X_11797_ _06473_ _06643_ net239 _06763_ vssd1 vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__a31o_1
X_14160__330 clknet_leaf_198_clk vssd1 vssd1 vccd1 vccd1 net1799 sky130_fd_sc_hd__inv_2
XFILLER_41_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xteam_08_1414 vssd1 vssd1 vccd1 vccd1 team_08_1414/HI ADR_O[30] sky130_fd_sc_hd__conb_1
X_16324_ clknet_leaf_67_clk _02533_ net1168 vssd1 vssd1 vccd1 vccd1 top.CPU.addressnew\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_159_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13536_ top.CPU.data_out\[26\] net590 net339 _02988_ vssd1 vssd1 vccd1 vccd1 _02524_
+ sky130_fd_sc_hd__o22a_1
X_10748_ _05626_ _05628_ net305 vssd1 vssd1 vccd1 vccd1 _06361_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08923__S net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11072__B2 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14457__627 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 net2096 sky130_fd_sc_hd__inv_2
Xteam_08_1425 vssd1 vssd1 vccd1 vccd1 team_08_1425/HI gpio_oeb[11] sky130_fd_sc_hd__conb_1
Xteam_08_1436 vssd1 vssd1 vccd1 vccd1 team_08_1436/HI gpio_out[21] sky130_fd_sc_hd__conb_1
Xteam_08_1447 vssd1 vssd1 vccd1 vccd1 team_08_1447/HI gpio_out[32] sky130_fd_sc_hd__conb_1
XFILLER_158_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xteam_08_1458 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] team_08_1458/LO sky130_fd_sc_hd__conb_1
XFILLER_145_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16255_ clknet_leaf_61_clk _02465_ net1160 vssd1 vssd1 vccd1 vccd1 top.CPU.alu.immediate\[31\]
+ sky130_fd_sc_hd__dfrtp_4
Xteam_08_1469 vssd1 vssd1 vccd1 vccd1 gpio_out[12] team_08_1469/LO sky130_fd_sc_hd__conb_1
X_13467_ net1396 net872 _02913_ net418 vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__a31o_1
XANTENNA__09017__A1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10679_ _06261_ _06294_ net305 vssd1 vssd1 vccd1 vccd1 _06295_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_93_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16368__RESET_B net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14201__371 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 net1840 sky130_fd_sc_hd__inv_2
X_15206_ net1540 _01416_ net1082 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_173_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12418_ _06920_ _06937_ _06939_ vssd1 vssd1 vccd1 vccd1 _06944_ sky130_fd_sc_hd__or3_1
XFILLER_127_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16186_ net2520 _02396_ net1243 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[986\]
+ sky130_fd_sc_hd__dfrtp_1
X_13398_ top.mmio.mem_data_i\[25\] net593 net1346 vssd1 vssd1 vccd1 vccd1 _02916_
+ sky130_fd_sc_hd__a21o_1
XFILLER_154_672 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12572__A1 top.CPU.done vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08776__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15137_ clknet_leaf_47_clk _01347_ net1130 vssd1 vssd1 vccd1 vccd1 top.I2C.data_out\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_12349_ net1340 top.I2C.output_state\[15\] net2968 vssd1 vssd1 vccd1 vccd1 _06897_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__11288__C _06471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_34_Left_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15068_ clknet_leaf_55_clk _00016_ net1134 vssd1 vssd1 vccd1 vccd1 top.I2C.output_state\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11127__A2 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12324__A1 _04188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07890_ top.CPU.registers.data\[476\] net1338 net870 top.CPU.registers.data\[508\]
+ net778 vssd1 vssd1 vccd1 vccd1 _03529_ sky130_fd_sc_hd__a221o_1
XFILLER_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11678__A3 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10886__A1 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07751__A1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09560_ top.CPU.registers.data\[544\] top.CPU.registers.data\[512\] net973 vssd1
+ vssd1 vccd1 vccd1 _05199_ sky130_fd_sc_hd__mux2_1
XFILLER_49_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08511_ net770 _04148_ _04149_ net694 vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__a31o_1
X_09491_ net947 _05129_ vssd1 vssd1 vccd1 vccd1 _05130_ sky130_fd_sc_hd__or2_1
XFILLER_82_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11835__B1 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_43_Left_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08700__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08442_ net709 _04079_ _04080_ _04078_ vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_102_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08373_ top.CPU.registers.data\[306\] top.CPU.registers.data\[274\] net818 vssd1
+ vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__mux2_1
XFILLER_149_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16616__A net1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout144_A _06290_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11063__B2 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11602__A3 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout311_A net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout409_A _05023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09559__A2 net1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08767__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16038__RESET_B net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11366__A2 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_52_Left_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1220_A net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1318_A net1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07973__A top.CPU.alu.program_counter\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09517__X _05156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout400 net401 vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__buf_2
XANTENNA_fanout680_A net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout411 net412 vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__clkbuf_4
Xfanout1409 top.CPU.control_unit.instruction\[4\] vssd1 vssd1 vccd1 vccd1 net1409
+ sky130_fd_sc_hd__buf_2
XANTENNA__12315__A1 _05361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout422 net423 vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__buf_6
XANTENNA_fanout778_A net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09716__C1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07692__B _03262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout433 _06602_ vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__clkbuf_8
XFILLER_101_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout444 net445 vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__buf_4
Xfanout455 _03330_ vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__clkbuf_4
XFILLER_113_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_126_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout466 net467 vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09192__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09827_ _05465_ vssd1 vssd1 vccd1 vccd1 _05466_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_6_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout477 _03193_ vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_161_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout488 net491 vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_161_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout566_X net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout499 net500 vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__buf_4
XANTENNA__07742__A1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout945_A net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09758_ top.CPU.registers.data_out_r1_prev\[27\] net875 net637 _05396_ _05394_ vssd1
+ vssd1 vccd1 vccd1 _05397_ sky130_fd_sc_hd__o221ai_4
XFILLER_73_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13815__B2 top.CPU.data_out\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09252__X _04891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08709_ top.CPU.registers.data\[237\] net1386 net807 top.CPU.registers.data\[205\]
+ net762 vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_61_Left_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11826__B1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09689_ net710 _05325_ _05326_ _05327_ vssd1 vssd1 vccd1 vccd1 _05328_ sky130_fd_sc_hd__a31o_1
XFILLER_42_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10839__A net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11434__S net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11720_ _06561_ net206 net423 net3042 vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__a22o_1
X_14144__314 clknet_leaf_112_clk vssd1 vssd1 vccd1 vccd1 net1783 sky130_fd_sc_hd__inv_2
XFILLER_154_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11651_ _06272_ net198 net424 net3323 vssd1 vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout900_X net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09247__A1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10602_ _05667_ _05827_ _05829_ _05671_ _06140_ vssd1 vssd1 vccd1 vccd1 _06222_ sky130_fd_sc_hd__o221a_1
XANTENNA__13502__X _02971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09839__S net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11054__B2 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09798__A2 net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11582_ net3010 net247 _06747_ net483 vssd1 vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__a22o_1
XFILLER_11_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13321_ top.I2C.data_out\[4\] net554 _02859_ top.mmio.mem_data_i\[4\] vssd1 vssd1
+ vccd1 vccd1 _02860_ sky130_fd_sc_hd__a22o_1
X_10533_ _04330_ _05569_ net445 vssd1 vssd1 vccd1 vccd1 _06156_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10801__A1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12265__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16040_ net2374 _02250_ net1099 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[840\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_70_Left_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13252_ net3917 _02805_ _02810_ _02803_ vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__a22o_1
X_10464_ _05998_ _06089_ net392 vssd1 vssd1 vccd1 vccd1 _06090_ sky130_fd_sc_hd__mux2_1
XFILLER_164_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11357__A2 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12203_ _06543_ _06868_ _06796_ vssd1 vssd1 vccd1 vccd1 _06869_ sky130_fd_sc_hd__or3b_1
XFILLER_109_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13183_ _02760_ _02761_ _02763_ top.I2C.within_byte_counter_writing\[2\] vssd1 vssd1
+ vccd1 vccd1 _02764_ sky130_fd_sc_hd__o211a_1
XFILLER_124_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10395_ net408 _06023_ vssd1 vssd1 vccd1 vccd1 _06024_ sky130_fd_sc_hd__nor2_1
XFILLER_151_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09574__S net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12134_ top.CPU.registers.data\[85\] net653 net244 vssd1 vssd1 vccd1 vccd1 _06835_
+ sky130_fd_sc_hd__o21a_1
XFILLER_151_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11109__A2 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07981__A1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11609__S net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09707__C1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12065_ net3905 net655 _06801_ vssd1 vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__o21a_1
X_11016_ net3812 net216 _06564_ net311 vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__a22o_1
XFILLER_65_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15824_ net2158 _02034_ net1154 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[624\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13806__B2 top.CPU.data_out\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07822__S net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12967_ top.I2C.bit_timer_counter\[1\] top.I2C.bit_timer_counter\[0\] _07401_ net1341
+ vssd1 vssd1 vccd1 vccd1 _07404_ sky130_fd_sc_hd__a31o_1
X_15755_ net2089 _01965_ net1065 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[555\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11918_ net3284 net187 net345 _06193_ vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__a22o_1
XANTENNA__11293__B2 _05808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12898_ _07341_ _07342_ vssd1 vssd1 vccd1 vccd1 _07343_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08219__A _03822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15686_ net2020 _01896_ net1073 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[486\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11832__A3 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11849_ net461 _06681_ net236 net153 net2689 vssd1 vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__a32o_1
XFILLER_159_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16549__RESET_B net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11045__B2 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12683__B _04919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_109_Left_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08997__B1 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11596__A2 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16307_ clknet_leaf_95_clk _02516_ net1262 vssd1 vssd1 vccd1 vccd1 top.CPU.data_out\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_173_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13519_ _04048_ net584 vssd1 vssd1 vccd1 vccd1 _02980_ sky130_fd_sc_hd__and2_1
XFILLER_119_639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08461__A2 net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload10 clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clkload10/Y sky130_fd_sc_hd__inv_8
Xclkload21 clknet_leaf_197_clk vssd1 vssd1 vccd1 vccd1 clkload21/Y sky130_fd_sc_hd__clkinv_16
XANTENNA__10915__C net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16238_ clknet_leaf_61_clk _02448_ net1160 vssd1 vssd1 vccd1 vccd1 top.CPU.control_unit.instruction\[14\]
+ sky130_fd_sc_hd__dfrtp_4
Xclkload32 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 clkload32/Y sky130_fd_sc_hd__clkinv_8
Xclkload43 clknet_leaf_187_clk vssd1 vssd1 vccd1 vccd1 clkload43/Y sky130_fd_sc_hd__clkinv_16
XFILLER_173_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload54 clknet_leaf_173_clk vssd1 vssd1 vccd1 vccd1 clkload54/Y sky130_fd_sc_hd__inv_4
XANTENNA__11348__A2 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload65 clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 clkload65/Y sky130_fd_sc_hd__inv_6
Xclkload76 clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 clkload76/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__10771__X _06383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16169_ net2503 _02379_ net1055 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[969\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload87 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 clkload87/Y sky130_fd_sc_hd__bufinv_16
Xclkload98 clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 clkload98/Y sky130_fd_sc_hd__inv_8
XANTENNA__11899__A3 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08991_ top.CPU.registers.data\[969\] net1309 net840 top.CPU.registers.data\[1001\]
+ net761 vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__a221o_1
XFILLER_173_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07942_ _03580_ vssd1 vssd1 vccd1 vccd1 _03581_ sky130_fd_sc_hd__inv_2
XFILLER_114_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14585__755 clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 net2224 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_118_Left_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_143_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07873_ top.CPU.registers.data\[572\] top.CPU.registers.data\[540\] net833 vssd1
+ vssd1 vccd1 vccd1 _03512_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07724__A1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09612_ top.CPU.registers.data\[576\] net1315 net844 top.CPU.registers.data\[608\]
+ net741 vssd1 vssd1 vccd1 vccd1 _05251_ sky130_fd_sc_hd__a221o_1
XANTENNA__08921__B1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07732__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14626__796 clknet_leaf_143_clk vssd1 vssd1 vccd1 vccd1 net2265 sky130_fd_sc_hd__inv_2
XANTENNA__15084__RESET_B net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09543_ top.CPU.registers.data\[449\] net1337 net866 top.CPU.registers.data\[481\]
+ net779 vssd1 vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout261_A net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout359_A _06704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11284__A1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09474_ net748 _05112_ vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__or2_1
XFILLER_64_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11823__A3 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08425_ top.CPU.registers.data\[81\] net1326 net857 top.CPU.registers.data\[113\]
+ net774 vssd1 vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__a221o_1
XANTENNA__09229__A1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1170_A net1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout147_X net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout526_A net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13322__X _02861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1268_A net1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11036__B2 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08356_ net744 _03994_ _03993_ vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13689__B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08563__S net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload4 clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clkload4/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_109_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08988__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11587__A2 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08287_ top.CPU.registers.data\[307\] top.CPU.registers.data\[275\] net825 vssd1
+ vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_119_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout314_X net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout895_A net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11339__A2 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07974__Y _03613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10180_ net305 _05700_ _05701_ _05815_ vssd1 vssd1 vccd1 vccd1 _05816_ sky130_fd_sc_hd__o31a_1
XFILLER_133_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout683_X net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1206 net1209 vssd1 vssd1 vccd1 vccd1 net1206 sky130_fd_sc_hd__clkbuf_4
XFILLER_121_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1217 net1218 vssd1 vssd1 vccd1 vccd1 net1217 sky130_fd_sc_hd__buf_2
XANTENNA__12114__A net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1228 net1229 vssd1 vssd1 vccd1 vccd1 net1228 sky130_fd_sc_hd__clkbuf_4
Xfanout230 _06772_ vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__clkbuf_4
Xfanout241 net242 vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__buf_4
Xfanout1239 net1240 vssd1 vssd1 vccd1 vccd1 net1239 sky130_fd_sc_hd__buf_2
Xfanout252 _06733_ vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__buf_4
Xfanout263 net264 vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__buf_4
XFILLER_87_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout850_X net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout274 _06714_ vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__buf_4
XFILLER_47_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout285 _06712_ vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__buf_6
XANTENNA_fanout948_X net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13644__S net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08912__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout296 _06662_ vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__clkbuf_4
XFILLER_101_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12821_ top.CPU.alu.program_counter\[17\] _07273_ net1359 vssd1 vssd1 vccd1 vccd1
+ _01180_ sky130_fd_sc_hd__mux2_1
XANTENNA__09012__S0 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10569__A _06190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12752_ net125 _07210_ vssd1 vssd1 vccd1 vccd1 _07211_ sky130_fd_sc_hd__or2_1
X_15540_ net1874 _01750_ net1073 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[340\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11814__A3 net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11703_ _06535_ net200 net421 net3187 vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__a22o_1
X_15471_ net1805 _01681_ net1094 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[271\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10856__X _06464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12683_ top.CPU.alu.program_counter\[5\] _04919_ vssd1 vssd1 vccd1 vccd1 _07148_
+ sky130_fd_sc_hd__or2_1
XANTENNA__12784__A top.CPU.alu.program_counter\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11634_ _05880_ net204 net426 net3506 vssd1 vssd1 vccd1 vccd1 _01917_ sky130_fd_sc_hd__a22o_1
XANTENNA__12224__B1 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11027__B2 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08979__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11578__A2 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11565_ _06676_ net258 net247 net2705 vssd1 vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__a22o_1
XANTENNA__08045__Y _03684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13304_ _06930_ _06936_ _02846_ vssd1 vssd1 vccd1 vccd1 _02847_ sky130_fd_sc_hd__and3_2
X_10516_ net415 _06139_ vssd1 vssd1 vccd1 vccd1 _06140_ sky130_fd_sc_hd__or2_2
X_11496_ net562 net480 _06628_ net254 net2850 vssd1 vssd1 vccd1 vccd1 _02028_ sky130_fd_sc_hd__a32o_1
X_13235_ _02789_ _02793_ vssd1 vssd1 vccd1 vccd1 _02801_ sky130_fd_sc_hd__nor2_1
X_16023_ net2357 _02233_ net1180 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[823\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_143_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10591__X _06212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10447_ _03989_ net504 vssd1 vssd1 vccd1 vccd1 _06074_ sky130_fd_sc_hd__nor2_1
X_14272__442 clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 net1911 sky130_fd_sc_hd__inv_2
XFILLER_156_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13166_ _02752_ _02751_ top.I2C.within_byte_counter_reading\[0\] vssd1 vssd1 vccd1
+ vccd1 _01334_ sky130_fd_sc_hd__mux2_1
X_10378_ _05993_ _05994_ _06007_ _05992_ vssd1 vssd1 vccd1 vccd1 _06008_ sky130_fd_sc_hd__a211o_1
X_14569__739 clknet_leaf_155_clk vssd1 vssd1 vccd1 vccd1 net2208 sky130_fd_sc_hd__inv_2
XFILLER_3_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07954__A1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11750__A2 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12117_ net3916 net657 _06826_ vssd1 vssd1 vccd1 vccd1 _01504_ sky130_fd_sc_hd__o21a_1
X_13097_ _06946_ _07426_ vssd1 vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__and2_1
XFILLER_111_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14313__483 clknet_leaf_157_clk vssd1 vssd1 vccd1 vccd1 net1952 sky130_fd_sc_hd__inv_2
X_12048_ _06595_ _06779_ net150 net3256 vssd1 vssd1 vccd1 vccd1 _01540_ sky130_fd_sc_hd__a22o_1
XANTENNA__11502__A2 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08648__S net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14947__Q top.CPU.alu.program_counter\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15807_ net2141 _02017_ net1224 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[607\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_93_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_66_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08667__C1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15738_ net2072 _01948_ net1250 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[538\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11588__A2_N _06726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13007__A2 _07429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15669_ net2003 _01879_ net1215 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[469\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08210_ top.CPU.registers.data\[343\] net1295 net1017 top.CPU.registers.data\[375\]
+ net937 vssd1 vssd1 vccd1 vccd1 _03849_ sky130_fd_sc_hd__a221o_1
XANTENNA__11802__S net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09190_ top.CPU.alu.program_counter\[6\] _04828_ net1034 vssd1 vssd1 vccd1 vccd1
+ _04829_ sky130_fd_sc_hd__mux2_2
XANTENNA__12215__B1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07890__B1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11569__A2 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08141_ top.CPU.registers.data\[469\] net1300 net1021 top.CPU.registers.data\[501\]
+ net917 vssd1 vssd1 vccd1 vccd1 _03780_ sky130_fd_sc_hd__a221o_1
XFILLER_159_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload110 clknet_leaf_156_clk vssd1 vssd1 vccd1 vccd1 clkload110/Y sky130_fd_sc_hd__clkinv_8
X_08072_ _03707_ _03708_ _03709_ _03710_ net674 vssd1 vssd1 vccd1 vccd1 _03711_ sky130_fd_sc_hd__a221o_1
XFILLER_146_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14859__1029 clknet_leaf_137_clk vssd1 vssd1 vccd1 vccd1 net2498 sky130_fd_sc_hd__inv_2
Xclkload121 clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 clkload121/Y sky130_fd_sc_hd__clkinv_8
Xclkload132 clknet_leaf_137_clk vssd1 vssd1 vccd1 vccd1 clkload132/Y sky130_fd_sc_hd__inv_12
XFILLER_20_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload143 clknet_leaf_151_clk vssd1 vssd1 vccd1 vccd1 clkload143/Y sky130_fd_sc_hd__clkinv_8
XFILLER_174_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload154 clknet_leaf_136_clk vssd1 vssd1 vccd1 vccd1 clkload154/Y sky130_fd_sc_hd__inv_16
XFILLER_161_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10942__A _06472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload165 clknet_leaf_125_clk vssd1 vssd1 vccd1 vccd1 clkload165/Y sky130_fd_sc_hd__inv_4
Xclkload176 clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 clkload176/Y sky130_fd_sc_hd__inv_8
Xclkload187 clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 clkload187/Y sky130_fd_sc_hd__clkinv_4
XFILLER_143_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08198__A1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_126_Left_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11741__A2 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08974_ top.CPU.registers.data\[233\] net1386 net805 top.CPU.registers.data\[201\]
+ net761 vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__a221o_1
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1016_A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09147__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold16 top.CPU.registers.data_out_r2_prev\[8\] vssd1 vssd1 vccd1 vccd1 net2573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 top.CPU.registers.data_out_r2_prev\[23\] vssd1 vssd1 vccd1 vccd1 net2584 sky130_fd_sc_hd__dlygate4sd3_1
X_07925_ net948 _03562_ _03563_ net958 vssd1 vssd1 vccd1 vccd1 _03564_ sky130_fd_sc_hd__o211a_1
Xhold38 _00029_ vssd1 vssd1 vccd1 vccd1 net2595 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 top.CPU.registers.data_out_r2_prev\[14\] vssd1 vssd1 vccd1 vccd1 net2606 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout476_A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07856_ top.CPU.registers.data\[829\] top.CPU.registers.data\[797\] net980 vssd1
+ vssd1 vccd1 vccd1 _03495_ sky130_fd_sc_hd__mux2_1
XANTENNA__10701__B1 _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07787_ _03421_ _03424_ _03425_ vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout264_X net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12049__A3 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout643_A net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09526_ net803 _05163_ _05164_ net699 vssd1 vssd1 vccd1 vccd1 _05165_ sky130_fd_sc_hd__a31o_1
XFILLER_43_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11257__B2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_135_Left_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09457_ top.CPU.registers.data\[226\] net1393 net823 top.CPU.registers.data\[194\]
+ net773 vssd1 vssd1 vccd1 vccd1 _05096_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout810_A net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout431_X net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout529_X net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout908_A net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08408_ net625 _04044_ _04045_ _04046_ vssd1 vssd1 vccd1 vccd1 _04047_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_156_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09388_ top.CPU.registers.data\[35\] top.CPU.registers.data\[3\] net828 vssd1 vssd1
+ vccd1 vccd1 _05027_ sky130_fd_sc_hd__mux2_1
XANTENNA__07881__B1 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_173_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08339_ net938 _03968_ _03969_ _03977_ net606 vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__a311o_1
XANTENNA__08425__A2 net1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09083__C1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12221__A3 _06796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11013__A net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07633__B1 net1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11350_ net3748 net285 net277 _06233_ vssd1 vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_134_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14256__426 clknet_leaf_200_clk vssd1 vssd1 vccd1 vccd1 net1895 sky130_fd_sc_hd__inv_2
XANTENNA__13639__S net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10301_ _03167_ _05933_ vssd1 vssd1 vccd1 vccd1 _05934_ sky130_fd_sc_hd__nor2_1
XANTENNA__11980__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11281_ net521 _06570_ vssd1 vssd1 vccd1 vccd1 _06698_ sky130_fd_sc_hd__nor2_1
XFILLER_153_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13020_ net2769 _07435_ net896 vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__mux2_1
X_10232_ net402 _05866_ vssd1 vssd1 vccd1 vccd1 _05867_ sky130_fd_sc_hd__or2_1
XANTENNA__09418__A net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14000__170 clknet_leaf_200_clk vssd1 vssd1 vccd1 vccd1 net1639 sky130_fd_sc_hd__inv_2
XANTENNA__11193__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11732__A2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10163_ _05651_ _05657_ net384 vssd1 vssd1 vccd1 vccd1 _05800_ sky130_fd_sc_hd__mux2_1
Xfanout1003 _03334_ vssd1 vssd1 vccd1 vccd1 net1003 sky130_fd_sc_hd__buf_4
Xfanout1014 net1015 vssd1 vssd1 vccd1 vccd1 net1014 sky130_fd_sc_hd__clkbuf_4
Xfanout1025 net1026 vssd1 vssd1 vccd1 vccd1 net1025 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1036 net1037 vssd1 vssd1 vccd1 vccd1 net1036 sky130_fd_sc_hd__clkbuf_8
XANTENNA_input37_A gpio_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1047 _03151_ vssd1 vssd1 vccd1 vccd1 net1047 sky130_fd_sc_hd__buf_2
X_10094_ _05726_ _05731_ net389 vssd1 vssd1 vccd1 vccd1 _05732_ sky130_fd_sc_hd__mux2_1
X_14971_ clknet_leaf_95_clk _01216_ net1260 vssd1 vssd1 vccd1 vccd1 top.SPI.paroutput\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09689__A1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1058 net1059 vssd1 vssd1 vccd1 vccd1 net1058 sky130_fd_sc_hd__clkbuf_4
Xfanout1069 net1075 vssd1 vssd1 vccd1 vccd1 net1069 sky130_fd_sc_hd__clkbuf_4
XFILLER_87_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10299__A2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11496__A1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11970__X _06777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12804_ _07254_ _07256_ vssd1 vssd1 vccd1 vccd1 _07258_ sky130_fd_sc_hd__nor2_1
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08649__C1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13784_ net12 net1051 net886 net3788 vssd1 vssd1 vccd1 vccd1 _02665_ sky130_fd_sc_hd__a22o_1
X_10996_ net515 net439 _06231_ net544 vssd1 vssd1 vccd1 vccd1 _06552_ sky130_fd_sc_hd__and4_1
XFILLER_163_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08113__A1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15523_ net1857 _01733_ net1207 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[323\]
+ sky130_fd_sc_hd__dfrtp_1
X_12735_ top.CPU.alu.program_counter\[10\] _04598_ vssd1 vssd1 vccd1 vccd1 _07195_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_26_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09861__A1 _05499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11622__S net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12666_ _07123_ _07127_ _07122_ vssd1 vssd1 vccd1 vccd1 _07133_ sky130_fd_sc_hd__a21o_1
X_15454_ net1788 _01664_ net1238 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[254\]
+ sky130_fd_sc_hd__dfrtp_1
X_11617_ net145 net3696 net212 vssd1 vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__mux2_1
XANTENNA__09074__C1 net1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12597_ top.SPI.count\[1\] _03142_ _03143_ top.SPI.count\[0\] vssd1 vssd1 vccd1 vccd1
+ _07098_ sky130_fd_sc_hd__o22a_1
X_15385_ net1719 _01595_ net1238 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[185\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_129_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12212__A3 _06796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11548_ _03181_ net461 net541 _06603_ vssd1 vssd1 vccd1 vccd1 _06739_ sky130_fd_sc_hd__or4_1
Xwire450 _04427_ vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__clkbuf_4
XFILLER_144_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold508 _01213_ vssd1 vssd1 vccd1 vccd1 net3065 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11971__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold519 top.CPU.registers.data\[360\] vssd1 vssd1 vccd1 vccd1 net3076 sky130_fd_sc_hd__dlygate4sd3_1
X_11479_ _06609_ net260 net256 net3146 vssd1 vssd1 vccd1 vccd1 _02045_ sky130_fd_sc_hd__a22o_1
XANTENNA__10762__A net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13218_ top.I2C.which_data_address\[2\] _02775_ vssd1 vssd1 vccd1 vccd1 _02791_ sky130_fd_sc_hd__nor2_1
XANTENNA__09377__B1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16006_ net2340 _02216_ net1080 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[806\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_143_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11723__A2 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13149_ _03118_ _07126_ vssd1 vssd1 vccd1 vccd1 _02741_ sky130_fd_sc_hd__nor2_1
XFILLER_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11296__C net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10931__B1 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1208 top.CPU.registers.data\[611\] vssd1 vssd1 vccd1 vccd1 net3765 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1219 top.CPU.registers.data\[581\] vssd1 vssd1 vccd1 vccd1 net3776 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07710_ top.CPU.control_unit.instruction\[24\] _03331_ vssd1 vssd1 vccd1 vccd1 _03349_
+ sky130_fd_sc_hd__or2_2
XANTENNA__11487__A1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08690_ _04294_ _04326_ vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__or2_1
X_07641_ _03161_ _03278_ _03279_ vssd1 vssd1 vccd1 vccd1 _03280_ sky130_fd_sc_hd__or3_1
XFILLER_26_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07572_ net776 _03207_ net726 _03210_ vssd1 vssd1 vccd1 vccd1 _03211_ sky130_fd_sc_hd__a211o_1
XFILLER_81_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11239__B2 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14697__867 clknet_leaf_155_clk vssd1 vssd1 vccd1 vccd1 net2336 sky130_fd_sc_hd__inv_2
X_09311_ net607 _04947_ _04949_ net627 vssd1 vssd1 vccd1 vccd1 _04950_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_24_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08655__A2 _04291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_807 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09242_ net702 _04876_ _04877_ net640 vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__a31o_1
XANTENNA__10462__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09002__S net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09173_ net704 _04810_ _04811_ _04808_ vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout224_A _05762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08124_ top.CPU.registers.data_out_r2_prev\[21\] net687 _03760_ _03762_ vssd1 vssd1
+ vccd1 vccd1 _03763_ sky130_fd_sc_hd__o22a_1
XANTENNA__07615__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10214__A2 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08841__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_151_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12871__B _03823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08055_ top.CPU.registers.data\[756\] net1379 net979 top.CPU.registers.data\[724\]
+ net905 vssd1 vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1133_A net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput39 net39 vssd1 vssd1 vccd1 vccd1 ADR_O[0] sky130_fd_sc_hd__buf_2
XANTENNA__10391__B _06019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07918__A1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11714__A2 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08040__B1 net1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1300_A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10922__B1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08957_ net1047 _04595_ vssd1 vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__and2_2
XANTENNA__13467__A2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout858_A _03203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout479_X net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11478__A1 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07908_ top.CPU.registers.data\[188\] net1025 net924 vssd1 vssd1 vccd1 vccd1 _03547_
+ sky130_fd_sc_hd__a21o_1
X_08888_ net702 _04504_ _04507_ _04522_ _04526_ vssd1 vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__o32a_1
XANTENNA__08879__C1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14641__811 clknet_leaf_188_clk vssd1 vssd1 vccd1 vccd1 net2280 sky130_fd_sc_hd__inv_2
XANTENNA__08343__A1 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07839_ top.CPU.registers.data\[61\] net1007 net931 vssd1 vssd1 vccd1 vccd1 _03478_
+ sky130_fd_sc_hd__a21o_1
XFILLER_112_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout646_X net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1290_X net1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1388_X net1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10850_ _06456_ _06457_ net394 vssd1 vssd1 vccd1 vccd1 _06458_ sky130_fd_sc_hd__a21oi_1
XFILLER_112_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09509_ top.CPU.registers.data\[225\] net1384 net998 top.CPU.registers.data\[193\]
+ net923 vssd1 vssd1 vccd1 vccd1 _05148_ sky130_fd_sc_hd__a221o_1
XFILLER_112_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10781_ net529 _06392_ vssd1 vssd1 vccd1 vccd1 _06393_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout813_X net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12520_ _07026_ _07027_ _07028_ vssd1 vssd1 vccd1 vccd1 _07029_ sky130_fd_sc_hd__or3_1
XANTENNA__08317__A _03955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_117_Right_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12451_ net1341 top.I2C.output_state\[19\] net2973 vssd1 vssd1 vccd1 vccd1 _06961_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_138_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11402_ _06531_ net281 net269 net2815 vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__a22o_1
XFILLER_172_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15170_ net1507 _01380_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r1_prev\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_12382_ top.CPU.handler.readout _03126_ top.CPU.addressnew\[17\] top.CPU.addressnew\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06920_ sky130_fd_sc_hd__or4b_1
XANTENNA__08803__C1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13369__S net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11333_ net3804 net285 net277 _05811_ vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__a22o_1
XFILLER_125_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09359__B1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11264_ net471 _06688_ vssd1 vssd1 vccd1 vccd1 _06689_ sky130_fd_sc_hd__nor2_1
XANTENNA__11397__B net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13003_ _07426_ _07428_ vssd1 vssd1 vccd1 vccd1 _07430_ sky130_fd_sc_hd__nand2_1
XFILLER_134_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11705__A2 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10215_ _03649_ _05300_ _05366_ _05503_ _05365_ vssd1 vssd1 vccd1 vccd1 _05850_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_37_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11195_ net3426 net297 _06655_ net323 vssd1 vssd1 vccd1 vccd1 _02255_ sky130_fd_sc_hd__a22o_1
XANTENNA__09582__S net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10146_ _05778_ _05782_ net401 vssd1 vssd1 vccd1 vccd1 _05783_ sky130_fd_sc_hd__mux2_1
XFILLER_67_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07790__C1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11617__S net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14954_ clknet_leaf_53_clk net2735 net1135 vssd1 vssd1 vccd1 vccd1 top.I2C.bit_timer_counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10077_ _04765_ net373 vssd1 vssd1 vccd1 vccd1 _05715_ sky130_fd_sc_hd__nor2_1
XFILLER_75_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12130__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14384__554 clknet_leaf_200_clk vssd1 vssd1 vccd1 vccd1 net2023 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_50_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_195_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_195_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12021__B _06781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14858__1028 clknet_leaf_145_clk vssd1 vssd1 vccd1 vccd1 net2497 sky130_fd_sc_hd__inv_2
XANTENNA_clkload2_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16624_ top.SPI.wrx vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12956__B top.CPU.alu.program_counter\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14425__595 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 net2064 sky130_fd_sc_hd__inv_2
X_13767_ net24 net1051 net886 net3929 vssd1 vssd1 vccd1 vccd1 _02648_ sky130_fd_sc_hd__a22o_1
XANTENNA__09295__C1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10979_ net518 net440 net132 net546 vssd1 vssd1 vccd1 vccd1 _06542_ sky130_fd_sc_hd__and4_1
XFILLER_15_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15506_ net1840 _01716_ net1102 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[306\]
+ sky130_fd_sc_hd__dfrtp_1
X_12718_ _07167_ _07179_ vssd1 vssd1 vccd1 vccd1 _07180_ sky130_fd_sc_hd__or2_1
XANTENNA__07845__B1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16486_ clknet_leaf_41_clk _02648_ net1116 vssd1 vssd1 vccd1 vccd1 top.mmio.mem_data_i\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13698_ net3450 _03052_ vssd1 vssd1 vccd1 vccd1 _02621_ sky130_fd_sc_hd__xor2_1
XFILLER_129_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15437_ net1771 _01647_ net1057 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[237\]
+ sky130_fd_sc_hd__dfrtp_1
X_12649_ net1411 net1341 net2926 vssd1 vssd1 vccd1 vccd1 _00016_ sky130_fd_sc_hd__and3_1
XANTENNA__09598__B1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12197__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15368_ net1702 _01578_ net1087 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[168\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_157_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09062__A2 net1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold305 top.CPU.registers.data\[321\] vssd1 vssd1 vccd1 vccd1 net2862 sky130_fd_sc_hd__dlygate4sd3_1
Xhold316 top.I2C.data_out\[29\] vssd1 vssd1 vccd1 vccd1 net2873 sky130_fd_sc_hd__dlygate4sd3_1
X_15299_ net1633 _01509_ net1212 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[99\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_57_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold327 top.CPU.fetch.current_ra\[15\] vssd1 vssd1 vccd1 vccd1 net2884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 top.CPU.registers.data\[293\] vssd1 vssd1 vccd1 vccd1 net2895 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold349 top.CPU.registers.data\[296\] vssd1 vssd1 vccd1 vccd1 net2906 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09860_ top.CPU.control_unit.instruction\[26\] net1046 net899 vssd1 vssd1 vccd1 vccd1
+ _05499_ sky130_fd_sc_hd__o21a_2
Xfanout807 net813 vssd1 vssd1 vccd1 vccd1 net807 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11100__B net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12911__S net1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08897__A top.CPU.alu.program_counter\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout818 net822 vssd1 vssd1 vccd1 vccd1 net818 sky130_fd_sc_hd__buf_4
XANTENNA__10904__B1 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout829 net831 vssd1 vssd1 vccd1 vccd1 net829 sky130_fd_sc_hd__clkbuf_4
X_13992__162 clknet_leaf_126_clk vssd1 vssd1 vccd1 vccd1 net1631 sky130_fd_sc_hd__inv_2
XANTENNA__09770__B1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11594__Y _06753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08811_ top.CPU.registers.data\[556\] top.CPU.registers.data\[524\] net978 vssd1
+ vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__mux2_1
XFILLER_97_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09791_ _05428_ _05429_ net455 vssd1 vssd1 vccd1 vccd1 _05430_ sky130_fd_sc_hd__mux2_1
XFILLER_100_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10380__A1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1005 top.CPU.registers.data\[832\] vssd1 vssd1 vccd1 vccd1 net3562 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1016 top.CPU.registers.data\[1020\] vssd1 vssd1 vccd1 vccd1 net3573 sky130_fd_sc_hd__dlygate4sd3_1
X_08742_ top.CPU.registers.data\[941\] top.CPU.registers.data\[909\] top.CPU.registers.data\[813\]
+ top.CPU.registers.data\[781\] net968 net1280 vssd1 vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__mux4_1
Xhold1027 top.CPU.registers.data\[726\] vssd1 vssd1 vccd1 vccd1 net3584 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1038 top.CPU.registers.data\[873\] vssd1 vssd1 vccd1 vccd1 net3595 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 net64 vssd1 vssd1 vccd1 vccd1 net3606 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12121__A2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08673_ net1285 _04310_ _04311_ vssd1 vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_186_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_186_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout174_A _06825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08876__A2 net1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16619__A net1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07624_ top.CPU.control_unit.instruction\[14\] net1400 vssd1 vssd1 vccd1 vccd1 _03263_
+ sky130_fd_sc_hd__or2_2
XFILLER_38_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07740__S net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13082__A0 top.CPU.data_out\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13314__Y _02855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07555_ _03184_ _03192_ vssd1 vssd1 vccd1 vccd1 _03194_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout341_A net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout439_A _05697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07486_ top.CPU.handler.writeout vssd1 vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_153_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09225_ top.CPU.registers.data\[261\] net1309 net841 top.CPU.registers.data\[293\]
+ net690 vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__a221o_1
XFILLER_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09038__C1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout606_A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1250_A net1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout227_X net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12188__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09156_ _04794_ vssd1 vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__inv_2
XANTENNA__12042__D1 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11396__B1 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08107_ net637 _03742_ _03745_ vssd1 vssd1 vccd1 vccd1 _03746_ sky130_fd_sc_hd__or3_1
X_09087_ _03342_ _04725_ _04712_ vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__a21oi_4
XANTENNA__08261__B1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_110_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_110_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1136_X net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08038_ top.CPU.registers.data\[916\] net1319 net850 top.CPU.registers.data\[948\]
+ net722 vssd1 vssd1 vccd1 vccd1 _03677_ sky130_fd_sc_hd__a221o_1
XFILLER_123_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold850 top.CPU.registers.data\[552\] vssd1 vssd1 vccd1 vccd1 net3407 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11148__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09436__S0 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout975_A net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold861 top.CPU.registers.data\[157\] vssd1 vssd1 vccd1 vccd1 net3418 sky130_fd_sc_hd__dlygate4sd3_1
Xhold872 top.CPU.registers.data\[333\] vssd1 vssd1 vccd1 vccd1 net3429 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10552__D net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12821__S net1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold883 top.CPU.registers.data\[337\] vssd1 vssd1 vccd1 vccd1 net3440 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_168_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09210__C1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1303_X net1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold894 top.CPU.registers.data\[825\] vssd1 vssd1 vccd1 vccd1 net3451 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_168_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10000_ _05637_ _05638_ net383 vssd1 vssd1 vccd1 vccd1 _05639_ sky130_fd_sc_hd__mux2_1
XFILLER_89_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14071__241 clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 net1710 sky130_fd_sc_hd__inv_2
X_09989_ _04891_ net377 vssd1 vssd1 vccd1 vccd1 _05628_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout763_X net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14368__538 clknet_leaf_112_clk vssd1 vssd1 vccd1 vccd1 net2007 sky130_fd_sc_hd__inv_2
XFILLER_103_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_129_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12112__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_177_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_177_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout930_X net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11951_ _06495_ net345 net230 net2988 vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__a22o_1
XANTENNA__08867__A2 net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14112__282 clknet_leaf_112_clk vssd1 vssd1 vccd1 vccd1 net1751 sky130_fd_sc_hd__inv_2
XANTENNA__13652__S net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14409__579 clknet_leaf_156_clk vssd1 vssd1 vccd1 vccd1 net2048 sky130_fd_sc_hd__inv_2
X_10902_ net487 net465 _06494_ net222 net3144 vssd1 vssd1 vccd1 vccd1 _02387_ sky130_fd_sc_hd__a32o_1
X_11882_ net143 net3016 net188 vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__mux2_1
XANTENNA__12776__B _04325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09431__A net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13621_ top.CPU.alu.program_counter\[29\] _05806_ net1351 vssd1 vssd1 vccd1 vccd1
+ _03039_ sky130_fd_sc_hd__mux2_1
XANTENNA__13073__A0 top.CPU.data_out\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10833_ net394 _06362_ _06440_ _06441_ net409 vssd1 vssd1 vccd1 vccd1 _06442_ sky130_fd_sc_hd__a221o_1
XANTENNA__12268__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13612__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11025__X _06570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16340_ clknet_leaf_68_clk _02549_ net1167 vssd1 vssd1 vccd1 vccd1 top.CPU.addressnew\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13552_ top.CPU.addressnew\[1\] _02997_ net580 vssd1 vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__mux2_1
X_10764_ _05057_ _05271_ _04990_ vssd1 vssd1 vccd1 vccd1 _06376_ sky130_fd_sc_hd__a21o_1
XANTENNA__09292__A2 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12503_ _04828_ _04855_ _07001_ vssd1 vssd1 vccd1 vccd1 _07012_ sky130_fd_sc_hd__nand3b_1
XFILLER_158_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16271_ clknet_leaf_60_clk _02481_ net1138 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.toreg\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13483_ _03107_ net1397 _03200_ _02935_ vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__o31a_1
X_10695_ top.CPU.fetch.current_ra\[8\] net1040 net633 top.CPU.handler.toreg\[8\] _06310_
+ vssd1 vssd1 vccd1 vccd1 _06311_ sky130_fd_sc_hd__a221o_4
XANTENNA__12179__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12434_ net898 _06953_ vssd1 vssd1 vccd1 vccd1 _00056_ sky130_fd_sc_hd__nor2_1
XFILLER_145_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15222_ net1556 _01432_ net1230 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_173_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11387__B1 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11926__A2 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12365_ net898 _06906_ vssd1 vssd1 vccd1 vccd1 _00052_ sky130_fd_sc_hd__nor2_1
X_15153_ clknet_leaf_42_clk _01363_ net1118 vssd1 vssd1 vccd1 vccd1 top.I2C.data_out\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_126_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_101_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_101_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11316_ net3743 net289 net357 net145 vssd1 vssd1 vccd1 vccd1 _02188_ sky130_fd_sc_hd__a22o_1
X_15084_ clknet_leaf_57_clk _00014_ net1145 vssd1 vssd1 vccd1 vccd1 top.I2C.byte_manager_done
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_153_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12296_ net2623 _04531_ net1067 vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__mux2_1
X_14810__980 clknet_leaf_165_clk vssd1 vssd1 vccd1 vccd1 net2449 sky130_fd_sc_hd__inv_2
XANTENNA__11139__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13976__146 clknet_leaf_167_clk vssd1 vssd1 vccd1 vccd1 net1615 sky130_fd_sc_hd__inv_2
XANTENNA__11558__D net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11247_ net486 net462 _06678_ net294 net2991 vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__a32o_1
XANTENNA__12887__B1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09201__C1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11178_ _05962_ net3741 net298 vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__mux2_1
XFILLER_80_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07763__C1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10129_ _05614_ _05766_ _05765_ _05699_ vssd1 vssd1 vccd1 vccd1 _05767_ sky130_fd_sc_hd__a211o_1
XANTENNA__14932__RESET_B net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15986_ net2320 _02196_ net1103 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[786\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08307__A1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12103__A2 _06770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14937_ clknet_leaf_74_clk _01183_ net1159 vssd1 vssd1 vccd1 vccd1 top.CPU.alu.program_counter\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_48_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_168_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_168_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_63_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13819_ net2749 net334 net327 top.CPU.data_out\[21\] vssd1 vssd1 vccd1 vccd1 _02699_
+ sky130_fd_sc_hd__a22o_1
XFILLER_51_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16538_ clknet_leaf_99_clk _02700_ net1257 vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07818__B1 top.CPU.control_unit.instruction\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_149_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16469_ clknet_leaf_88_clk _02631_ net1272 vssd1 vssd1 vccd1 vccd1 top.SPI.timem\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15791__RESET_B net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09010_ _04647_ _04648_ net1366 vssd1 vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__o21a_1
XFILLER_136_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11589__Y _06748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08391__S net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09035__A2 net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11378__B1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10934__B net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11917__A2 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09059__Y _04698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold102 top.CPU.addressnew\[31\] vssd1 vssd1 vccd1 vccd1 net2659 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 _01207_ vssd1 vssd1 vccd1 vccd1 net2670 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10050__B1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold124 top.CPU.registers.data\[307\] vssd1 vssd1 vccd1 vccd1 net2681 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07597__A2 net1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold135 top.CPU.registers.data\[289\] vssd1 vssd1 vccd1 vccd1 net2692 sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 _01208_ vssd1 vssd1 vccd1 vccd1 net2703 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 top.CPU.registers.data\[519\] vssd1 vssd1 vccd1 vccd1 net2714 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 top.CPU.registers.data\[561\] vssd1 vssd1 vccd1 vccd1 net2725 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09912_ _05127_ _05550_ vssd1 vssd1 vccd1 vccd1 _05551_ sky130_fd_sc_hd__and2_1
Xhold179 top.CPU.registers.data\[41\] vssd1 vssd1 vccd1 vccd1 net2736 sky130_fd_sc_hd__dlygate4sd3_1
X_14055__225 clknet_leaf_184_clk vssd1 vssd1 vccd1 vccd1 net1694 sky130_fd_sc_hd__inv_2
XANTENNA__10950__A net1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout604 net605 vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__buf_4
Xfanout615 net616 vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__buf_4
XANTENNA__08546__A1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout626 net630 vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__buf_4
X_09843_ top.CPU.registers.data_out_r2_prev\[26\] net688 net621 _05475_ _05481_ vssd1
+ vssd1 vccd1 vccd1 _05482_ sky130_fd_sc_hd__o2111a_1
Xfanout637 net639 vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10353__A1 _03315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout648 net650 vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__buf_2
XANTENNA_fanout291_A net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout659 net660 vssd1 vssd1 vccd1 vccd1 net659 sky130_fd_sc_hd__buf_4
XANTENNA__11550__B1 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07754__C1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout389_A net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_146_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09774_ top.CPU.registers.data\[603\] net1297 net1019 top.CPU.registers.data\[635\]
+ net939 vssd1 vssd1 vccd1 vccd1 _05413_ sky130_fd_sc_hd__a221o_1
XFILLER_37_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_163_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08725_ net878 _04361_ _04332_ vssd1 vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_107_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_159_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_159_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12877__A _07322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10949__X _06524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08849__A2 net1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_174_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13472__S net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout556_A _02847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout177_X net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1298_A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08656_ net878 _04291_ _04293_ vssd1 vssd1 vccd1 vccd1 _04295_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_124_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11853__A1 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_54_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07607_ top.CPU.control_unit.instruction\[4\] top.CPU.control_unit.instruction\[6\]
+ net1278 vssd1 vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__or3_2
XANTENNA__09251__A _04889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08587_ net878 _04222_ _04224_ vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__o21a_1
XANTENNA__09259__C1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout723_A net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout344_X net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07538_ _03104_ _03105_ net1279 vssd1 vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__and3_1
XANTENNA__10408__A2 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_189_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14753__923 clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 net2392 sky130_fd_sc_hd__inv_2
XANTENNA__10813__C1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout511_X net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07469_ net1391 vssd1 vssd1 vccd1 vccd1 _03109_ sky130_fd_sc_hd__inv_2
XFILLER_168_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_69_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout609_X net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09208_ net625 _04843_ _04844_ net610 vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__a31o_1
X_10480_ _03167_ net551 net501 _06105_ vssd1 vssd1 vccd1 vccd1 _06106_ sky130_fd_sc_hd__or4b_1
XFILLER_136_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10844__B _05266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11369__B1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_112_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11908__A2 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09139_ top.CPU.registers.data_out_r2_prev\[7\] net687 net621 _04770_ _04777_ vssd1
+ vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__o2111a_1
XFILLER_135_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08234__B1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11021__A net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08785__A1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07588__A2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14857__1027 clknet_leaf_155_clk vssd1 vssd1 vccd1 vccd1 net2496 sky130_fd_sc_hd__inv_2
X_12150_ top.CPU.registers.data\[77\] net646 net244 vssd1 vssd1 vccd1 vccd1 _06843_
+ sky130_fd_sc_hd__o21a_1
XFILLER_163_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout880_X net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11101_ net3589 net304 _06608_ net321 vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout978_X net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13647__S net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12869__A0 top.CPU.alu.program_counter\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12081_ net563 net361 _06620_ net179 top.CPU.registers.data\[112\] vssd1 vssd1 vccd1
+ vccd1 _06809_ sky130_fd_sc_hd__a32o_1
XFILLER_1_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10860__A net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold680 top.CPU.registers.data\[366\] vssd1 vssd1 vccd1 vccd1 net3237 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_127_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold691 top.CPU.registers.data\[277\] vssd1 vssd1 vccd1 vccd1 net3248 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08537__A1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11032_ _03180_ _03182_ vssd1 vssd1 vccd1 vccd1 _06575_ sky130_fd_sc_hd__or2_4
XFILLER_2_889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10344__A1 _03822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07745__C1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16320__Q top.CPU.data_out\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15840_ net2174 _02050_ net1090 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[640\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07760__A2 net1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15771_ net2105 _01981_ net1216 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[571\]
+ sky130_fd_sc_hd__dfrtp_1
X_12983_ top.I2C.bit_timer_counter\[3\] _07407_ _07414_ vssd1 vssd1 vccd1 vccd1 _07415_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09498__C1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1380 _01333_ vssd1 vssd1 vccd1 vccd1 net3937 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1391 top.CPU.registers.data\[109\] vssd1 vssd1 vccd1 vccd1 net3948 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11844__A1 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11934_ top.CPU.registers.data\[223\] net232 vssd1 vssd1 vccd1 vccd1 _06773_ sky130_fd_sc_hd__and2_1
XFILLER_60_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11865_ _06703_ net241 net190 net2905 vssd1 vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__a22o_1
XFILLER_60_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13604_ net3253 _03029_ net583 vssd1 vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__mux2_1
X_10816_ _06418_ _06419_ _06421_ _06425_ vssd1 vssd1 vccd1 vccd1 _06426_ sky130_fd_sc_hd__o211a_2
X_11796_ top.CPU.registers.data\[351\] net158 vssd1 vssd1 vccd1 vccd1 _06763_ sky130_fd_sc_hd__and2_1
XFILLER_159_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16323_ clknet_leaf_66_clk _02532_ net1165 vssd1 vssd1 vccd1 vccd1 top.CPU.addressnew\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13535_ _05498_ net585 vssd1 vssd1 vccd1 vccd1 _02988_ sky130_fd_sc_hd__and2_1
XANTENNA__11072__A2 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08473__B1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14496__666 clknet_leaf_126_clk vssd1 vssd1 vccd1 vccd1 net2135 sky130_fd_sc_hd__inv_2
Xteam_08_1415 vssd1 vssd1 vccd1 vccd1 team_08_1415/HI ADR_O[31] sky130_fd_sc_hd__conb_1
X_10747_ net389 _06279_ vssd1 vssd1 vccd1 vccd1 _06360_ sky130_fd_sc_hd__nor2_1
XFILLER_159_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xteam_08_1426 vssd1 vssd1 vccd1 vccd1 team_08_1426/HI gpio_oeb[12] sky130_fd_sc_hd__conb_1
XANTENNA__09670__C1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_08_1437 vssd1 vssd1 vccd1 vccd1 team_08_1437/HI gpio_out[22] sky130_fd_sc_hd__conb_1
Xteam_08_1448 vssd1 vssd1 vccd1 vccd1 team_08_1448/HI gpio_out[33] sky130_fd_sc_hd__conb_1
X_16254_ clknet_leaf_60_clk _02464_ net1138 vssd1 vssd1 vccd1 vccd1 top.CPU.control_unit.instruction\[30\]
+ sky130_fd_sc_hd__dfrtp_2
Xteam_08_1459 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] team_08_1459/LO sky130_fd_sc_hd__conb_1
X_10678_ _04634_ net372 _05714_ vssd1 vssd1 vccd1 vccd1 _06294_ sky130_fd_sc_hd__o21ba_1
X_13466_ top.CPU.handler.toreg\[22\] _02954_ net120 vssd1 vssd1 vccd1 vccd1 _02488_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_93_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15205_ net1539 _01415_ net1065 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_12417_ top.CPU.addressnew\[0\] top.CPU.addressnew\[1\] top.CPU.addressnew\[13\]
+ top.CPU.addressnew\[12\] vssd1 vssd1 vccd1 vccd1 _06943_ sky130_fd_sc_hd__or4b_1
XFILLER_154_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16185_ net2519 _02395_ net1243 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[985\]
+ sky130_fd_sc_hd__dfrtp_1
X_13397_ top.CPU.control_unit.instruction\[24\] _02915_ net671 vssd1 vssd1 vccd1 vccd1
+ _02458_ sky130_fd_sc_hd__mux2_1
XFILLER_127_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07579__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14039__209 clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 net1678 sky130_fd_sc_hd__inv_2
XANTENNA__12572__A2 _06462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15136_ clknet_leaf_46_clk _01346_ net1137 vssd1 vssd1 vccd1 vccd1 top.I2C.data_out\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_154_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12348_ net898 _06896_ vssd1 vssd1 vccd1 vccd1 _00066_ sky130_fd_sc_hd__nor2_1
XANTENNA__10583__A1 _05667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11288__D net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10583__B2 _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11780__B1 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07984__C1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15067_ clknet_leaf_55_clk _00046_ net1134 vssd1 vssd1 vccd1 vccd1 top.I2C.output_state\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_12279_ _05397_ _06887_ _06888_ vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__o21ai_1
XFILLER_4_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11532__B1 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10886__A2 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15969_ net2303 _02179_ net1250 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[769\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10099__A0 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12697__A net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08894__B _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11805__S net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08510_ top.CPU.registers.data\[912\] net1322 net853 top.CPU.registers.data\[944\]
+ net721 vssd1 vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_69_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09490_ top.CPU.registers.data\[33\] top.CPU.registers.data\[1\] net998 vssd1 vssd1
+ vccd1 vccd1 _05129_ sky130_fd_sc_hd__mux2_1
XANTENNA__08386__S net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08441_ top.CPU.registers.data\[977\] net1326 net857 top.CPU.registers.data\[1009\]
+ net725 vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__a221o_1
X_14440__610 clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 net2079 sky130_fd_sc_hd__inv_2
XFILLER_23_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14737__907 clknet_leaf_190_clk vssd1 vssd1 vccd1 vccd1 net2376 sky130_fd_sc_hd__inv_2
XFILLER_51_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13588__A1 _06147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08372_ top.CPU.registers.data\[82\] net1320 net851 top.CPU.registers.data\[114\]
+ net769 vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__a221o_1
XANTENNA__11599__A0 _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12260__A1 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11063__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout137_A _05771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10271__B1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08216__A0 _03854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12582__D _06918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout304_A _06604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13906__76 clknet_leaf_192_clk vssd1 vssd1 vccd1 vccd1 net1545 sky130_fd_sc_hd__inv_2
XANTENNA__11771__B1 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07973__B net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08519__A1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout401 net405 vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__buf_2
Xfanout412 _04958_ vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07990__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout423 _06758_ vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__clkbuf_8
XFILLER_48_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout434 _06602_ vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__clkbuf_4
Xfanout445 _05521_ vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__buf_4
XFILLER_141_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout673_A net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11523__B1 _06734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout294_X net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout456 net463 vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09826_ net780 _05450_ _05451_ _05464_ vssd1 vssd1 vccd1 vccd1 _05465_ sky130_fd_sc_hd__a31o_2
Xfanout467 _03194_ vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout478 net479 vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1001_X net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout489 net490 vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12079__A1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13276__B1 top.CPU.control_unit.instruction\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09757_ net696 _05382_ _05385_ _05395_ _05379_ vssd1 vssd1 vccd1 vccd1 _05396_ sky130_fd_sc_hd__o32a_1
XANTENNA_fanout840_A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout461_X net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout938_A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10629__A2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08708_ top.CPU.registers.data\[173\] top.CPU.registers.data\[141\] net807 vssd1
+ vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__mux2_1
XFILLER_104_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09688_ net698 _05323_ _05324_ net638 vssd1 vssd1 vccd1 vccd1 _05327_ sky130_fd_sc_hd__a31o_1
XANTENNA__08152__C1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10839__B _06447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08639_ net792 _04276_ _04277_ net720 vssd1 vssd1 vccd1 vccd1 _04278_ sky130_fd_sc_hd__o211a_1
X_14183__353 clknet_leaf_183_clk vssd1 vssd1 vccd1 vccd1 net1822 sky130_fd_sc_hd__inv_2
XANTENNA_fanout1370_X net1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout726_X net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11650_ _06255_ net196 net424 net3818 vssd1 vssd1 vccd1 vccd1 _01901_ sky130_fd_sc_hd__a22o_1
XFILLER_168_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10601_ net406 _06041_ vssd1 vssd1 vccd1 vccd1 _06221_ sky130_fd_sc_hd__nand2_1
XANTENNA__08455__B1 _04092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11581_ _06562_ _06731_ vssd1 vssd1 vccd1 vccd1 _06747_ sky130_fd_sc_hd__nor2_1
XANTENNA__12251__A1 _06056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11054__A2 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14224__394 clknet_leaf_198_clk vssd1 vssd1 vccd1 vccd1 net1863 sky130_fd_sc_hd__inv_2
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13320_ _03130_ net598 net592 vssd1 vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__and3_1
X_10532_ _04330_ _06153_ _04327_ vssd1 vssd1 vccd1 vccd1 _06155_ sky130_fd_sc_hd__o21ai_1
XFILLER_80_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10801__A2 _06410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10463_ _06039_ _06088_ net307 vssd1 vssd1 vccd1 vccd1 _06089_ sky130_fd_sc_hd__mux2_1
X_13251_ top.I2C.data_out\[10\] net891 _02780_ vssd1 vssd1 vccd1 vccd1 _02810_ sky130_fd_sc_hd__mux2_1
XFILLER_136_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_73 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09404__C1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12202_ top.CPU.registers.data\[50\] net648 vssd1 vssd1 vccd1 vccd1 _06868_ sky130_fd_sc_hd__nor2_1
X_13182_ top.I2C.within_byte_counter_writing\[0\] top.I2C.which_data_address\[2\]
+ _02762_ top.I2C.within_byte_counter_writing\[1\] vssd1 vssd1 vccd1 vccd1 _02763_
+ sky130_fd_sc_hd__a22o_1
XFILLER_164_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10394_ _05912_ _06022_ net390 vssd1 vssd1 vccd1 vccd1 _06023_ sky130_fd_sc_hd__mux2_1
XFILLER_123_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10565__A1 _04325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11762__B1 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12133_ net3944 net175 _06834_ _06488_ vssd1 vssd1 vccd1 vccd1 _01496_ sky130_fd_sc_hd__a22o_1
XFILLER_123_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13503__A1 top.CPU.data_out\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09707__B1 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13503__B2 _02971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12064_ net568 net364 _06611_ net179 top.CPU.registers.data\[121\] vssd1 vssd1 vccd1
+ vccd1 _06801_ sky130_fd_sc_hd__a32o_1
XANTENNA__08605__S1 net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07718__C1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11015_ net514 _06374_ net542 vssd1 vssd1 vccd1 vccd1 _06564_ sky130_fd_sc_hd__and3_1
XANTENNA__09183__A1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13920__90 clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 net1559 sky130_fd_sc_hd__inv_2
Xfanout990 net994 vssd1 vssd1 vccd1 vccd1 net990 sky130_fd_sc_hd__buf_4
XFILLER_93_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15823_ net2157 _02033_ net1094 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[623\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_92_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11625__S net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15754_ net2088 _01964_ net1090 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[554\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11817__A1 _06213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12966_ top.I2C.bit_timer_counter\[0\] _07401_ net3992 vssd1 vssd1 vccd1 vccd1 _07403_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_80_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11917_ net3753 net185 net343 _06175_ vssd1 vssd1 vccd1 vccd1 _01649_ sky130_fd_sc_hd__a22o_1
XANTENNA__11293__A2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15685_ net2019 _01895_ net1083 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[485\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12897_ _07326_ _07331_ vssd1 vssd1 vccd1 vccd1 _07342_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_47_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10536__A1_N net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11848_ _06680_ net243 net152 net2676 vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__a22o_1
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11045__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12242__A1 _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11779_ net461 _06622_ net236 net161 net3237 vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__a32o_1
XANTENNA__10239__B1_N net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16306_ clknet_leaf_95_clk _02515_ net1262 vssd1 vssd1 vccd1 vccd1 top.CPU.data_out\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13518_ top.CPU.data_out\[17\] net590 net340 _02979_ vssd1 vssd1 vccd1 vccd1 _02515_
+ sky130_fd_sc_hd__o22a_1
XFILLER_9_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16237_ clknet_leaf_46_clk _02447_ net1137 vssd1 vssd1 vccd1 vccd1 top.CPU.control_unit.instruction\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload11 clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clkload11/Y sky130_fd_sc_hd__inv_12
X_13449_ net890 _02888_ _02937_ _02939_ vssd1 vssd1 vccd1 vccd1 _02946_ sky130_fd_sc_hd__a31o_1
Xclkload22 clknet_leaf_198_clk vssd1 vssd1 vccd1 vccd1 clkload22/Y sky130_fd_sc_hd__inv_16
XFILLER_62_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload33 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 clkload33/Y sky130_fd_sc_hd__clkinv_8
Xclkload44 clknet_leaf_188_clk vssd1 vssd1 vccd1 vccd1 clkload44/Y sky130_fd_sc_hd__inv_6
XANTENNA__08749__A1 net1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload55 clknet_leaf_175_clk vssd1 vssd1 vccd1 vccd1 clkload55/Y sky130_fd_sc_hd__clkinv_8
XFILLER_6_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16168_ net2502 _02378_ net1098 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[968\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload66 clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 clkload66/Y sky130_fd_sc_hd__clkinv_4
Xclkload77 clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 clkload77/Y sky130_fd_sc_hd__clkinv_4
XFILLER_127_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11753__B1 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload88 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 clkload88/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__07957__C1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload99 clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 clkload99/Y sky130_fd_sc_hd__clkinv_8
XFILLER_126_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15119_ net1501 _01332_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r2_prev\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_142_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16099_ net2433 _02309_ net1206 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[899\]
+ sky130_fd_sc_hd__dfrtp_1
X_08990_ top.CPU.registers.data\[937\] top.CPU.registers.data\[905\] net805 vssd1
+ vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__mux2_1
XFILLER_170_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07941_ _03578_ _03579_ vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__and2b_1
XFILLER_87_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11505__B1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07709__C1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09174__A1 _03111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07872_ _03476_ _03509_ vssd1 vssd1 vccd1 vccd1 _03511_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_143_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09611_ _05246_ _05249_ net636 vssd1 vssd1 vccd1 vccd1 _05250_ sky130_fd_sc_hd__a21o_1
XFILLER_18_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11520__A3 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10499__X _06124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14167__337 clknet_leaf_171_clk vssd1 vssd1 vccd1 vccd1 net1806 sky130_fd_sc_hd__inv_2
X_09542_ net802 _05179_ _05180_ net734 vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__o211a_1
XANTENNA__09477__A2 net1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08134__C1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14856__1026 clknet_leaf_126_clk vssd1 vssd1 vccd1 vccd1 net2495 sky130_fd_sc_hd__inv_2
XANTENNA__11284__A2 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09473_ top.CPU.registers.data\[546\] top.CPU.registers.data\[514\] net823 vssd1
+ vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__mux2_1
XFILLER_52_833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_90_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_90_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout254_A _06728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12218__D1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08424_ top.CPU.registers.data\[49\] top.CPU.registers.data\[17\] net825 vssd1 vssd1
+ vccd1 vccd1 _04063_ sky130_fd_sc_hd__mux2_1
X_14208__378 clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 net1847 sky130_fd_sc_hd__inv_2
XANTENNA__11036__A2 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08355_ top.CPU.registers.data\[562\] top.CPU.registers.data\[530\] net818 vssd1
+ vssd1 vccd1 vccd1 _03994_ sky130_fd_sc_hd__mux2_1
XFILLER_11_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08437__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10675__A net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout421_A net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1163_A net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout519_A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload5 clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clkload5/Y sky130_fd_sc_hd__inv_8
X_08286_ _03723_ _03789_ _03924_ vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__or3_1
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11992__B1 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1330_A net1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09675__S net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout790_A net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09401__A2 net1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10547__B2 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11744__B1 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07948__C1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07963__A2 net1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1207 net1209 vssd1 vssd1 vccd1 vccd1 net1207 sky130_fd_sc_hd__clkbuf_2
Xfanout1218 net1233 vssd1 vssd1 vccd1 vccd1 net1218 sky130_fd_sc_hd__buf_2
Xfanout220 _06469_ vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__buf_6
XFILLER_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12114__B net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout231 _06772_ vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__clkbuf_8
Xfanout1229 net1233 vssd1 vssd1 vccd1 vccd1 net1229 sky130_fd_sc_hd__buf_2
XANTENNA__09165__A1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout676_X net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout242 net243 vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__clkbuf_4
Xfanout253 _06733_ vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__buf_2
Xfanout264 net266 vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__buf_6
XFILLER_19_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout275 net279 vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__buf_4
XANTENNA__07715__A2 net1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout286 _06712_ vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07923__S net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout297 _06645_ vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11953__B net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09809_ top.CPU.registers.data\[282\] net1337 net867 top.CPU.registers.data\[314\]
+ net699 vssd1 vssd1 vccd1 vccd1 _05448_ sky130_fd_sc_hd__a221o_1
XFILLER_86_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout843_X net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12820_ _07272_ _07269_ net128 vssd1 vssd1 vccd1 vccd1 _07273_ sky130_fd_sc_hd__mux2_1
XANTENNA__09012__S1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09468__A2 net1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12751_ _07208_ _07209_ vssd1 vssd1 vccd1 vccd1 _07210_ sky130_fd_sc_hd__nor2_1
XFILLER_27_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_81_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_70_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11702_ _06534_ net209 net423 net2950 vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__a22o_1
XFILLER_15_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15470_ net1804 _01680_ net1193 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[270\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08754__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12682_ top.CPU.alu.program_counter\[5\] _04919_ vssd1 vssd1 vccd1 vccd1 _07147_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_139_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12224__A1 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11633_ _05849_ net206 net427 net3093 vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__a22o_1
XANTENNA__11027__A2 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11564_ _06675_ net260 net248 net2824 vssd1 vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__a22o_1
XANTENNA__10786__A1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11983__B1 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13303_ top.CPU.addressnew\[16\] top.CPU.addressnew\[19\] _06921_ _02845_ vssd1 vssd1
+ vccd1 vccd1 _02846_ sky130_fd_sc_hd__and4b_1
XFILLER_156_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10515_ _05665_ _05672_ vssd1 vssd1 vccd1 vccd1 _06139_ sky130_fd_sc_hd__nor2_4
X_11495_ net562 net478 _06627_ net254 net2957 vssd1 vssd1 vccd1 vccd1 _02029_ sky130_fd_sc_hd__a32o_1
XFILLER_171_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_982 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16022_ net2356 _02232_ net1228 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[822\]
+ sky130_fd_sc_hd__dfrtp_1
X_10446_ net408 _05861_ _06072_ _05742_ vssd1 vssd1 vccd1 vccd1 _06073_ sky130_fd_sc_hd__a211o_1
X_13234_ net2816 _02776_ _02800_ vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__mux2_1
XFILLER_124_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11735__B1 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13165_ top.I2C.output_state\[20\] top.I2C.initiate_read_bit _06950_ vssd1 vssd1
+ vccd1 vccd1 _02752_ sky130_fd_sc_hd__and3_1
X_10377_ net224 _06006_ _06004_ vssd1 vssd1 vccd1 vccd1 _06007_ sky130_fd_sc_hd__o21ai_2
XFILLER_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08600__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11750__A3 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12116_ net137 net365 net356 net175 top.CPU.registers.data\[94\] vssd1 vssd1 vccd1
+ vccd1 _06826_ sky130_fd_sc_hd__a32o_1
X_13096_ top.CPU.data_out\[31\] net2778 net558 vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__mux2_1
XANTENNA__13488__A0 top.CPU.data_out\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13897__67 clknet_leaf_159_clk vssd1 vssd1 vccd1 vccd1 net1536 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_88_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12047_ net3851 net149 _06778_ vssd1 vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__mux2_1
XFILLER_78_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12160__B1 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08903__A1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07706__A2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10710__A1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15806_ net2140 _02016_ net1202 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[606\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09459__A2 net1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15737_ net2071 _01947_ net1243 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[537\]
+ sky130_fd_sc_hd__dfrtp_1
X_12949_ top.CPU.alu.program_counter\[30\] _07381_ vssd1 vssd1 vccd1 vccd1 _07389_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__08667__B1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13660__B1 _03126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_72_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08664__S net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15668_ net2002 _01878_ net1112 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[468\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12215__A1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15599_ net1933 _01809_ net1095 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[399\]
+ sky130_fd_sc_hd__dfrtp_1
X_08140_ top.CPU.registers.data\[341\] net1300 net1021 top.CPU.registers.data\[373\]
+ net940 vssd1 vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__a221o_1
XANTENNA__13302__C top.CPU.done vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11974__B1 net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload100 clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 clkload100/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_140_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07642__A1 net1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08071_ top.CPU.registers.data\[308\] net1008 net931 vssd1 vssd1 vccd1 vccd1 _03710_
+ sky130_fd_sc_hd__a21oi_1
Xclkload111 clknet_leaf_157_clk vssd1 vssd1 vccd1 vccd1 clkload111/Y sky130_fd_sc_hd__inv_2
X_14552__722 clknet_leaf_169_clk vssd1 vssd1 vccd1 vccd1 net2191 sky130_fd_sc_hd__inv_2
Xclkload122 clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 clkload122/Y sky130_fd_sc_hd__clkinv_8
XFILLER_134_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload133 clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 clkload133/Y sky130_fd_sc_hd__inv_16
XANTENNA__09495__S net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10731__B1_N _06139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload144 clknet_leaf_152_clk vssd1 vssd1 vccd1 vccd1 clkload144/Y sky130_fd_sc_hd__inv_6
XFILLER_134_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload155 clknet_leaf_138_clk vssd1 vssd1 vccd1 vccd1 clkload155/Y sky130_fd_sc_hd__inv_16
Xclkload166 clknet_leaf_80_clk vssd1 vssd1 vccd1 vccd1 clkload166/Y sky130_fd_sc_hd__inv_8
XFILLER_162_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11726__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload177 clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 clkload177/Y sky130_fd_sc_hd__inv_8
XANTENNA__09395__A1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload188 clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 clkload188/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_114_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13479__B1 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08973_ net783 _04611_ vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__or2_1
XFILLER_103_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold17 top.CPU.registers.data_out_r2_prev\[24\] vssd1 vssd1 vccd1 vccd1 net2574 sky130_fd_sc_hd__dlygate4sd3_1
X_07924_ top.CPU.registers.data\[924\] net1303 net1026 top.CPU.registers.data\[956\]
+ net920 vssd1 vssd1 vccd1 vccd1 _03563_ sky130_fd_sc_hd__a221o_1
Xhold28 top.CPU.registers.data_out_r2_prev\[1\] vssd1 vssd1 vccd1 vccd1 net2585 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08839__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold39 top.CPU.registers.data_out_r1_prev\[4\] vssd1 vssd1 vccd1 vccd1 net2596 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09698__A2 net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1009_A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07855_ top.CPU.registers.data\[989\] net1288 net1007 top.CPU.registers.data\[1021\]
+ net906 vssd1 vssd1 vccd1 vccd1 _03494_ sky130_fd_sc_hd__a221o_1
XFILLER_84_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout469_A net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08370__A2 net1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07786_ top.CPU.registers.data_out_r2_prev\[30\] net688 net958 vssd1 vssd1 vccd1
+ vccd1 _03425_ sky130_fd_sc_hd__o21a_1
XFILLER_45_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09525_ top.CPU.registers.data\[961\] net1335 net868 top.CPU.registers.data\[993\]
+ net732 vssd1 vssd1 vccd1 vccd1 _05164_ sky130_fd_sc_hd__a221o_1
XANTENNA__11257__A2 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1280_A net1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09855__C1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_63_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__13480__S net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout257_X net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout636_A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1378_A net1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09456_ top.CPU.registers.data\[162\] top.CPU.registers.data\[130\] net823 vssd1
+ vssd1 vccd1 vccd1 _05095_ sky130_fd_sc_hd__mux2_1
XFILLER_169_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08407_ net618 _04042_ _04043_ net604 vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_156_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout424_X net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09387_ top.CPU.registers.data\[323\] net1328 net859 top.CPU.registers.data\[355\]
+ net775 vssd1 vssd1 vccd1 vccd1 _05026_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout803_A net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10217__B1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08338_ net677 _03966_ _03967_ net913 vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_173_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09083__B1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11965__B1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08269_ top.CPU.registers.data\[566\] top.CPU.registers.data\[534\] net998 vssd1
+ vssd1 vccd1 vccd1 _03908_ sky130_fd_sc_hd__mux2_1
XFILLER_126_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1333_X net1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14295__465 clknet_leaf_172_clk vssd1 vssd1 vccd1 vccd1 net1934 sky130_fd_sc_hd__inv_2
X_10300_ net602 _05931_ _05932_ vssd1 vssd1 vccd1 vccd1 _05933_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_134_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12509__A2 _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16093__RESET_B net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11280_ net2932 net295 _06697_ net316 vssd1 vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__a22o_1
XFILLER_146_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout793_X net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11717__B1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10231_ _05639_ _05646_ net387 vssd1 vssd1 vccd1 vccd1 _05866_ sky130_fd_sc_hd__mux2_1
XANTENNA__08189__A2 net1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11193__A1 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10162_ _05618_ _05783_ _05794_ _05798_ vssd1 vssd1 vccd1 vccd1 _05799_ sky130_fd_sc_hd__o211a_1
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout960_X net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1004 net1032 vssd1 vssd1 vccd1 vccd1 net1004 sky130_fd_sc_hd__buf_4
XFILLER_126_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1015 net1017 vssd1 vssd1 vccd1 vccd1 net1015 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13655__S net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1026 net1031 vssd1 vssd1 vccd1 vccd1 net1026 sky130_fd_sc_hd__clkbuf_2
X_14970_ clknet_leaf_84_clk _01215_ net1261 vssd1 vssd1 vccd1 vccd1 top.SPI.paroutput\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10093_ _05728_ _05730_ net385 vssd1 vssd1 vccd1 vccd1 _05731_ sky130_fd_sc_hd__mux2_1
Xfanout1037 _03199_ vssd1 vssd1 vccd1 vccd1 net1037 sky130_fd_sc_hd__buf_4
XFILLER_0_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1048 _03150_ vssd1 vssd1 vccd1 vccd1 net1048 sky130_fd_sc_hd__buf_2
XFILLER_120_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1059 net1068 vssd1 vssd1 vccd1 vccd1 net1059 sky130_fd_sc_hd__buf_2
XANTENNA__12142__B1 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11496__A2 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08361__A2 net1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12803_ top.CPU.alu.program_counter\[15\] _04256_ _07237_ _07255_ _07254_ vssd1 vssd1
+ vccd1 vccd1 _07257_ sky130_fd_sc_hd__o221a_1
XFILLER_56_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13783_ net11 net1051 net886 net3633 vssd1 vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_54_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_clk sky130_fd_sc_hd__clkbuf_8
X_10995_ net3239 net216 _06551_ net311 vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__a22o_1
XFILLER_55_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09310__A1 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10456__B1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15522_ net1856 _01732_ net1173 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[322\]
+ sky130_fd_sc_hd__dfrtp_1
X_12734_ top.CPU.alu.program_counter\[10\] _04598_ vssd1 vssd1 vccd1 vccd1 _07194_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_26_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15453_ net1787 _01663_ net1112 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[253\]
+ sky130_fd_sc_hd__dfrtp_1
X_12665_ _07130_ _07131_ vssd1 vssd1 vccd1 vccd1 _07132_ sky130_fd_sc_hd__and2_1
XFILLER_169_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11616_ net142 net3396 net212 vssd1 vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__mux2_1
X_14536__706 clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 net2175 sky130_fd_sc_hd__inv_2
XFILLER_156_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09074__B1 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15384_ net1718 _01594_ net1150 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[184\]
+ sky130_fd_sc_hd__dfrtp_1
X_12596_ _07095_ _07096_ vssd1 vssd1 vccd1 vccd1 _07097_ sky130_fd_sc_hd__nand2_1
XANTENNA__09613__A2 net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11956__B1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11547_ net481 net130 net354 net250 net2933 vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__a32o_1
XANTENNA__11420__A2 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire451 _03682_ vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__clkbuf_2
XFILLER_156_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold509 top.CPU.registers.data\[890\] vssd1 vssd1 vccd1 vccd1 net3066 sky130_fd_sc_hd__dlygate4sd3_1
X_11478_ net492 net477 _06608_ net257 net2998 vssd1 vssd1 vccd1 vccd1 _02046_ sky130_fd_sc_hd__a32o_1
XANTENNA__10762__B net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11708__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09377__A1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16005_ net2339 _02215_ net1062 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[805\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_59_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13217_ net3823 _02779_ _02790_ _02773_ vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_59_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10429_ net659 _06056_ vssd1 vssd1 vccd1 vccd1 _06057_ sky130_fd_sc_hd__and2_2
XFILLER_124_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14855__1025 clknet_leaf_184_clk vssd1 vssd1 vccd1 vccd1 net2494 sky130_fd_sc_hd__inv_2
XANTENNA__07927__A2 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_1006 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13148_ _03106_ _05232_ vssd1 vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__nand2_1
XFILLER_112_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10931__A1 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13079_ top.CPU.data_out\[14\] net3373 net559 vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__mux2_1
XFILLER_25_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1209 top.CPU.registers.data_out_r1_prev\[14\] vssd1 vssd1 vccd1 vccd1 net3766
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08337__C1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14958__Q top.SPI.busy vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11487__A2 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07640_ net1398 _03259_ _03263_ _03248_ vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__a31o_1
XANTENNA__10695__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07571_ top.CPU.registers.data\[735\] net1392 net829 top.CPU.registers.data\[767\]
+ net798 vssd1 vssd1 vccd1 vccd1 _03210_ sky130_fd_sc_hd__o221a_1
XANTENNA__11239__A2 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09837__C1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_45_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_81_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09310_ net957 _04925_ _04948_ vssd1 vssd1 vccd1 vccd1 _04949_ sky130_fd_sc_hd__a21o_1
XFILLER_22_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09241_ net691 _04878_ _04879_ vssd1 vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__and3_1
XFILLER_167_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11114__A net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16533__RESET_B net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09172_ top.CPU.registers.data\[326\] net1317 net847 top.CPU.registers.data\[358\]
+ net767 vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__a221o_1
X_14279__449 clknet_leaf_185_clk vssd1 vssd1 vccd1 vccd1 net1918 sky130_fd_sc_hd__inv_2
XANTENNA__09604__A2 net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08123_ net627 _03761_ net612 vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__a21o_1
XANTENNA__11947__B1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11411__A2 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10953__A net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout217_A net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14023__193 clknet_leaf_184_clk vssd1 vssd1 vccd1 vccd1 net1662 sky130_fd_sc_hd__inv_2
X_08054_ net953 _03687_ _03689_ _03692_ vssd1 vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__a31o_1
XANTENNA__11962__A3 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08576__C1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10922__A1 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08591__A2 net1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08956_ net1041 net1039 vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__nor2_1
XFILLER_103_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08328__C1 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12124__B1 _06749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07907_ top.CPU.registers.data\[28\] net996 _03545_ vssd1 vssd1 vccd1 vccd1 _03546_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__08879__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11478__A2 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08887_ net737 _04524_ _04525_ net690 vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout753_A net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14680__850 clknet_leaf_170_clk vssd1 vssd1 vccd1 vccd1 net2319 sky130_fd_sc_hd__inv_2
X_07838_ top.CPU.control_unit.instruction\[29\] net1046 net899 vssd1 vssd1 vccd1 vccd1
+ _03477_ sky130_fd_sc_hd__o21a_1
XFILLER_71_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout920_A net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07769_ _03153_ _03155_ net1363 vssd1 vssd1 vccd1 vccd1 _03408_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout541_X net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1283_X net1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_36_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout639_X net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13504__A _04497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09508_ top.CPU.registers.data\[65\] net1307 net1030 top.CPU.registers.data\[97\]
+ net947 vssd1 vssd1 vccd1 vccd1 _05147_ sky130_fd_sc_hd__a221o_1
X_14721__891 clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 net2360 sky130_fd_sc_hd__inv_2
X_10780_ net552 net502 net147 vssd1 vssd1 vccd1 vccd1 _06392_ sky130_fd_sc_hd__or3b_1
XANTENNA__09843__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09439_ top.CPU.registers.data\[834\] net1294 net1015 top.CPU.registers.data\[866\]
+ net936 vssd1 vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__a221o_1
XFILLER_12_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11650__A2 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout806_X net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12450_ _06905_ _06908_ _06910_ net1054 net3969 vssd1 vssd1 vccd1 vccd1 _00046_ sky130_fd_sc_hd__a32o_1
XFILLER_8_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11938__B1 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11401_ _06530_ net283 net267 net3201 vssd1 vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__a22o_1
XANTENNA__13510__Y _02975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12381_ top.CPU.handler.readout _03126_ vssd1 vssd1 vccd1 vccd1 _06919_ sky130_fd_sc_hd__nor2_1
XFILLER_126_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11402__A2 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08803__B1 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11332_ net3494 net288 net283 _05772_ vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__a22o_1
XFILLER_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08333__A net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11263_ net514 _06557_ vssd1 vssd1 vccd1 vccd1 _06688_ sky130_fd_sc_hd__or2_1
XFILLER_106_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13002_ _07426_ _07428_ vssd1 vssd1 vccd1 vccd1 _07429_ sky130_fd_sc_hd__and2_2
XANTENNA__08567__C1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07909__A2 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10214_ net3573 net227 net321 _05849_ vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__a22o_1
X_11194_ _06213_ net429 vssd1 vssd1 vccd1 vccd1 _06655_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_37_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10145_ _05781_ vssd1 vssd1 vccd1 vccd1 _05782_ sky130_fd_sc_hd__inv_2
XFILLER_122_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13867__37 clknet_leaf_122_clk vssd1 vssd1 vccd1 vccd1 net1506 sky130_fd_sc_hd__inv_2
XFILLER_43_1031 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12115__B1 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07790__B1 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14953_ clknet_leaf_53_clk _01199_ net1136 vssd1 vssd1 vccd1 vccd1 top.I2C.bit_timer_counter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10076_ _04698_ net380 vssd1 vssd1 vccd1 vccd1 _05714_ sky130_fd_sc_hd__nor2_1
XFILLER_153_83 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10677__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10103__A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16623_ top.I2C.scl_out vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__clkbuf_1
XANTENNA__13615__A0 top.CPU.alu.program_counter\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12729__S net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09819__C1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_27_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08098__A1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13766_ net13 net1051 net886 net3932 vssd1 vssd1 vccd1 vccd1 _02647_ sky130_fd_sc_hd__a22o_1
XANTENNA__09295__B1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10978_ net440 net132 net543 vssd1 vssd1 vccd1 vccd1 _06541_ sky130_fd_sc_hd__and3_1
XFILLER_16_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09834__A2 net1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15505_ net1839 _01715_ net1189 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[305\]
+ sky130_fd_sc_hd__dfrtp_1
X_12717_ _07158_ _07159_ _07168_ _07156_ vssd1 vssd1 vccd1 vccd1 _07179_ sky130_fd_sc_hd__o211a_1
XANTENNA__07845__A1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16485_ clknet_leaf_41_clk _02647_ net1115 vssd1 vssd1 vccd1 vccd1 top.mmio.mem_data_i\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11641__A2 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13697_ _03052_ _03053_ vssd1 vssd1 vccd1 vccd1 _02620_ sky130_fd_sc_hd__nor2_1
XFILLER_31_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15436_ net1770 _01646_ net1070 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[236\]
+ sky130_fd_sc_hd__dfrtp_1
X_12648_ top.I2C.bit_timer_state\[1\] net1339 net2791 vssd1 vssd1 vccd1 vccd1 _00017_
+ sky130_fd_sc_hd__and3_1
XFILLER_30_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11929__B1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_154_Left_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14007__177 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 net1646 sky130_fd_sc_hd__inv_2
X_15367_ net1701 _01577_ net1198 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[167\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_96_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12579_ _03246_ _07051_ _07052_ _03137_ vssd1 vssd1 vccd1 vccd1 _07084_ sky130_fd_sc_hd__a31o_1
XFILLER_7_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15298_ net1632 _01508_ net1175 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[98\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold306 top.CPU.registers.data\[393\] vssd1 vssd1 vccd1 vccd1 net2863 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold317 top.CPU.registers.data\[330\] vssd1 vssd1 vccd1 vccd1 net2874 sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 top.CPU.registers.data\[429\] vssd1 vssd1 vccd1 vccd1 net2885 sky130_fd_sc_hd__dlygate4sd3_1
Xhold339 top.SPI.paroutput\[27\] vssd1 vssd1 vccd1 vccd1 net2896 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16233__Q top.CPU.control_unit.instruction\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_74_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09626__X _05265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08022__A1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11100__C net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout808 net813 vssd1 vssd1 vccd1 vccd1 net808 sky130_fd_sc_hd__clkbuf_4
Xfanout819 net822 vssd1 vssd1 vccd1 vccd1 net819 sky130_fd_sc_hd__buf_2
XANTENNA__10904__A1 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08897__B net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08573__A2 net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11808__S net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08810_ top.CPU.registers.data\[940\] top.CPU.registers.data\[908\] top.CPU.registers.data\[812\]
+ top.CPU.registers.data\[780\] net977 net1282 vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__mux4_1
XFILLER_86_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09790_ top.CPU.control_unit.instruction\[27\] net1046 _03408_ vssd1 vssd1 vccd1
+ vccd1 _05429_ sky130_fd_sc_hd__o21a_2
XANTENNA__12052__X _06795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08389__S net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12106__B1 _03185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14664__834 clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 net2303 sky130_fd_sc_hd__inv_2
XFILLER_97_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10380__A2 _06008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1006 top.CPU.registers.data\[326\] vssd1 vssd1 vccd1 vccd1 net3563 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07781__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_163_Left_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1017 top.CPU.registers.data\[144\] vssd1 vssd1 vccd1 vccd1 net3574 sky130_fd_sc_hd__dlygate4sd3_1
X_08741_ top.CPU.registers.data\[845\] net1371 net968 top.CPU.registers.data\[877\]
+ net1280 vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__o221a_1
XANTENNA__10117__C1 _05754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1028 top.CPU.registers.data\[824\] vssd1 vssd1 vccd1 vccd1 net3585 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1039 top.SPI.paroutput\[30\] vssd1 vssd1 vccd1 vccd1 net3596 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1390 net1395 vssd1 vssd1 vccd1 vccd1 net1390 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08325__A2 net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08672_ top.CPU.registers.data\[846\] net1378 net981 top.CPU.registers.data\[878\]
+ net1282 vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_109_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705__875 clknet_leaf_188_clk vssd1 vssd1 vccd1 vccd1 net2344 sky130_fd_sc_hd__inv_2
XFILLER_53_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07623_ _03104_ net1278 _03154_ vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__or3_4
XFILLER_26_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13881__51 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 net1520 sky130_fd_sc_hd__inv_2
XANTENNA__10948__A net1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_18_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout167_A _06757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07554_ _03184_ _03192_ vssd1 vssd1 vccd1 vccd1 _03193_ sky130_fd_sc_hd__and2_4
X_07485_ top.I2C.byte_manager_done vssd1 vssd1 vccd1 vccd1 _03125_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11632__A2 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_172_Left_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09224_ top.CPU.registers.data\[37\] top.CPU.registers.data\[5\] net806 vssd1 vssd1
+ vccd1 vccd1 _04863_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_170_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13385__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09155_ _04792_ _04793_ net453 vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__mux2_1
XFILLER_21_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout122_X net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout501_A _05696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1243_A net1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08106_ net798 _03743_ _03744_ net728 vssd1 vssd1 vccd1 vccd1 _03745_ sky130_fd_sc_hd__o211a_1
XFILLER_147_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11935__A3 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09086_ _03116_ _04720_ _04723_ _04724_ vssd1 vssd1 vccd1 vccd1 _04725_ sky130_fd_sc_hd__a31o_1
XFILLER_135_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08037_ top.CPU.registers.data\[820\] top.CPU.registers.data\[788\] net817 vssd1
+ vssd1 vccd1 vccd1 _03676_ sky130_fd_sc_hd__mux2_1
XFILLER_162_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1031_X net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold840 top.CPU.registers.data\[940\] vssd1 vssd1 vccd1 vccd1 net3397 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11148__A1 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09436__S1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold851 top.CPU.registers.data\[484\] vssd1 vssd1 vccd1 vccd1 net3408 sky130_fd_sc_hd__dlygate4sd3_1
Xhold862 top.CPU.registers.data\[787\] vssd1 vssd1 vccd1 vccd1 net3419 sky130_fd_sc_hd__dlygate4sd3_1
Xhold873 top.CPU.registers.data\[495\] vssd1 vssd1 vccd1 vccd1 net3430 sky130_fd_sc_hd__dlygate4sd3_1
Xhold884 top.CPU.registers.data\[1018\] vssd1 vssd1 vccd1 vccd1 net3441 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09210__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout491_X net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11699__A2 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout870_A _03203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold895 top.CPU.registers.data\[662\] vssd1 vssd1 vccd1 vccd1 net3452 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_168_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08564__A2 net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout968_A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10622__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09988_ _05625_ _05626_ vssd1 vssd1 vccd1 vccd1 _05627_ sky130_fd_sc_hd__nor2_1
XFILLER_77_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08939_ _04576_ _04577_ net673 vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__o21a_1
XFILLER_29_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_150_Right_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout756_X net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08316__A2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09513__A1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11950_ _06494_ net349 net231 net3240 vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_28_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11320__B2 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10901_ net139 net437 vssd1 vssd1 vccd1 vccd1 _06494_ sky130_fd_sc_hd__and2_1
XFILLER_123_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11961__B net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11871__A2 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout923_X net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11881_ net146 net3489 net189 vssd1 vssd1 vccd1 vccd1 _01682_ sky130_fd_sc_hd__mux2_1
XANTENNA__11453__S net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13620_ net2823 _03038_ net582 vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_142_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10832_ net381 _05620_ _05622_ net386 vssd1 vssd1 vccd1 vccd1 _06441_ sky130_fd_sc_hd__o31a_1
XANTENNA__09277__B1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09816__A2 net1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14854__1024 clknet_leaf_123_clk vssd1 vssd1 vccd1 vccd1 net2493 sky130_fd_sc_hd__inv_2
XFILLER_25_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13551_ top.CPU.alu.program_counter\[1\] _06445_ net1351 vssd1 vssd1 vccd1 vccd1
+ _02997_ sky130_fd_sc_hd__mux2_1
XANTENNA__16318__Q top.CPU.data_out\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10763_ net3909 net225 net312 _06375_ vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__a22o_1
XFILLER_41_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12502_ _04828_ _04855_ vssd1 vssd1 vccd1 vccd1 _07011_ sky130_fd_sc_hd__xnor2_1
XFILLER_157_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16270_ clknet_leaf_60_clk _02480_ net1139 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.toreg\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13482_ net2919 _02962_ net120 vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__mux2_1
X_10694_ net600 _06309_ vssd1 vssd1 vccd1 vccd1 _06310_ sky130_fd_sc_hd__nor2_1
XFILLER_12_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10864__Y _06471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15221_ net1555 _01431_ net1227 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_12433_ net1339 top.I2C.output_state\[10\] net3892 vssd1 vssd1 vccd1 vccd1 _06953_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__10593__A net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15152_ clknet_leaf_42_clk _01362_ net1117 vssd1 vssd1 vccd1 vccd1 top.I2C.data_out\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_12364_ net1339 top.I2C.output_state\[28\] net2944 vssd1 vssd1 vccd1 vccd1 _06906_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_39_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11315_ net3292 net289 net357 net142 vssd1 vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__a22o_1
X_15083_ clknet_leaf_56_clk _00040_ net1145 vssd1 vssd1 vccd1 vccd1 top.I2C.byte_manager_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_141_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11139__A1 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12295_ net3801 _04428_ net1077 vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__mux2_1
X_14351__521 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 net1990 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_91_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08004__A1 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14648__818 clknet_leaf_161_clk vssd1 vssd1 vccd1 vccd1 net2287 sky130_fd_sc_hd__inv_2
X_11246_ net516 _06546_ vssd1 vssd1 vccd1 vccd1 _06678_ sky130_fd_sc_hd__nor2_2
XFILLER_122_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09752__A1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10898__B1 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11177_ net494 _06483_ _06648_ net300 net3100 vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__a32o_1
XFILLER_122_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10128_ _03444_ _05524_ _05613_ net445 vssd1 vssd1 vccd1 vccd1 _05766_ sky130_fd_sc_hd__a31oi_1
X_15985_ net2319 _02195_ net1193 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[785\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10104__Y _05742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14936_ clknet_leaf_74_clk _01182_ net1159 vssd1 vssd1 vccd1 vccd1 top.CPU.alu.program_counter\[19\]
+ sky130_fd_sc_hd__dfrtp_4
X_10059_ _03184_ _03185_ vssd1 vssd1 vccd1 vccd1 _05697_ sky130_fd_sc_hd__nand2b_4
XANTENNA__08712__C1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09622__A net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09964__A_N _05601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11862__A2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13818_ net3121 net335 net328 top.CPU.data_out\[20\] vssd1 vssd1 vccd1 vccd1 _02698_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16196__RESET_B net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13064__A1 top.CPU.data_out\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11590__C net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16537_ clknet_leaf_99_clk _02699_ net1257 vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07818__A1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13749_ _03084_ _03085_ vssd1 vssd1 vccd1 vccd1 _02640_ sky130_fd_sc_hd__nor2_1
XFILLER_92_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16468_ clknet_leaf_86_clk _02630_ net1272 vssd1 vssd1 vccd1 vccd1 top.SPI.timem\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_148_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13367__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15419_ net1753 _01629_ net1213 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[219\]
+ sky130_fd_sc_hd__dfrtp_1
X_16399_ clknet_leaf_62_clk net670 net1161 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.state\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_117_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08243__A1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold103 top.CPU.registers.data\[395\] vssd1 vssd1 vccd1 vccd1 net2660 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10050__A1 _03148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold114 top.CPU.registers.data\[546\] vssd1 vssd1 vccd1 vccd1 net2671 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10790__X _06401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold125 top.CPU.registers.data\[810\] vssd1 vssd1 vccd1 vccd1 net2682 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12922__S net1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold136 top.CPU.registers.data\[800\] vssd1 vssd1 vccd1 vccd1 net2693 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_160_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold147 top.CPU.registers.data\[547\] vssd1 vssd1 vccd1 vccd1 net2704 sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 top.I2C.I2C_state\[24\] vssd1 vssd1 vccd1 vccd1 net2715 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_137_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09911_ _05195_ _05547_ _05549_ vssd1 vssd1 vccd1 vccd1 _05550_ sky130_fd_sc_hd__a21o_1
X_14094__264 clknet_leaf_121_clk vssd1 vssd1 vccd1 vccd1 net1733 sky130_fd_sc_hd__inv_2
Xhold169 top.SPI.parameters\[19\] vssd1 vssd1 vccd1 vccd1 net2726 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10950__B net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout605 _03349_ vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__buf_4
XANTENNA__09743__A1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout616 _03343_ vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__buf_2
XANTENNA__10442__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09842_ net682 _05476_ _05477_ _05480_ net615 vssd1 vssd1 vccd1 vccd1 _05481_ sky130_fd_sc_hd__a311o_1
Xfanout627 net630 vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__buf_4
XFILLER_140_560 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout638 net639 vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__clkbuf_8
XFILLER_101_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout649 net650 vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__buf_4
XANTENNA__07754__B1 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ top.CPU.registers.data\[763\] net1381 net991 top.CPU.registers.data\[731\]
+ net916 vssd1 vssd1 vccd1 vccd1 _05412_ sky130_fd_sc_hd__a221o_1
XFILLER_100_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout284_A _06713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08724_ net878 _04361_ _04332_ vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__o21a_2
XFILLER_37_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_7_0_clk_X clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08847__S net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08703__C1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08655_ net878 _04291_ _04293_ vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__o21ai_4
XFILLER_96_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_87_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout549_A net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07606_ top.CPU.control_unit.instruction\[14\] net1397 vssd1 vssd1 vccd1 vccd1 _03245_
+ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_1_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09259__B1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08586_ net879 _04222_ _04224_ vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__o21ai_4
XFILLER_53_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08148__A _03755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11066__B1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07537_ net1401 net660 vssd1 vssd1 vccd1 vccd1 _03176_ sky130_fd_sc_hd__nand2_1
XFILLER_23_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11605__A2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1360_A net1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout716_A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14792__962 clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 net2431 sky130_fd_sc_hd__inv_2
X_07468_ net1398 vssd1 vssd1 vccd1 vccd1 _03108_ sky130_fd_sc_hd__inv_2
XANTENNA__08482__A1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09207_ top.CPU.registers.data\[742\] net1379 net977 top.CPU.registers.data\[710\]
+ net904 vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__a221o_1
XFILLER_33_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11369__A1 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11302__A net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09138_ net608 _04773_ _04776_ vssd1 vssd1 vccd1 vccd1 _04777_ sky130_fd_sc_hd__or3_1
X_13999__169 clknet_leaf_192_clk vssd1 vssd1 vccd1 vccd1 net1638 sky130_fd_sc_hd__inv_2
X_14335__505 clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 net1974 sky130_fd_sc_hd__inv_2
XANTENNA__12832__S net1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09069_ top.CPU.registers.data\[72\] net1373 net969 top.CPU.registers.data\[104\]
+ net901 vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__o221a_1
XFILLER_163_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11100_ net574 net532 net442 _05848_ vssd1 vssd1 vccd1 vccd1 _06608_ sky130_fd_sc_hd__and4_1
XFILLER_150_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12080_ _06619_ net349 net178 net3070 vssd1 vssd1 vccd1 vccd1 _01523_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout873_X net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold670 top.CPU.registers.data\[573\] vssd1 vssd1 vccd1 vccd1 net3227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold681 top.CPU.registers.data\[934\] vssd1 vssd1 vccd1 vccd1 net3238 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09734__A1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09195__C1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11448__S net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold692 top.CPU.registers.data\[541\] vssd1 vssd1 vccd1 vccd1 net3249 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_34_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11031_ _03180_ _03182_ vssd1 vssd1 vccd1 vccd1 _06574_ sky130_fd_sc_hd__nor2_1
XANTENNA__07745__B1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08942__C1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15770_ net2104 _01980_ net1250 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[570\]
+ sky130_fd_sc_hd__dfrtp_1
X_12982_ top.I2C.bit_timer_counter\[5\] top.I2C.bit_timer_counter\[4\] top.I2C.bit_timer_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 _07414_ sky130_fd_sc_hd__and3_1
XANTENNA__12097__A2 _06770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1370 top.I2C.data_out\[4\] vssd1 vssd1 vccd1 vccd1 net3927 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input12_A DAT_I[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1381 top.CPU.registers.data\[928\] vssd1 vssd1 vccd1 vccd1 net3938 sky130_fd_sc_hd__dlygate4sd3_1
X_11933_ net435 net341 vssd1 vssd1 vccd1 vccd1 _06772_ sky130_fd_sc_hd__nand2_8
Xhold1392 top.CPU.addressnew\[15\] vssd1 vssd1 vccd1 vccd1 net3949 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11183__S net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11864_ net564 _03180_ _03181_ _06751_ vssd1 vssd1 vccd1 vccd1 _06767_ sky130_fd_sc_hd__or4_1
XFILLER_73_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13603_ top.CPU.alu.program_counter\[21\] _06031_ net1348 vssd1 vssd1 vccd1 vccd1
+ _03029_ sky130_fd_sc_hd__mux2_1
XANTENNA__11057__B1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10815_ net370 _06422_ _06424_ vssd1 vssd1 vccd1 vccd1 _06425_ sky130_fd_sc_hd__o21a_1
X_11795_ _06644_ _06751_ vssd1 vssd1 vccd1 vccd1 _06762_ sky130_fd_sc_hd__nor2_2
X_16322_ clknet_leaf_67_clk _02531_ net1168 vssd1 vssd1 vccd1 vccd1 top.CPU.addressnew\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13534_ net4005 net590 net340 _02987_ vssd1 vssd1 vccd1 vccd1 _02523_ sky130_fd_sc_hd__o22a_1
XANTENNA__07897__A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10746_ _05273_ _05543_ _06358_ net370 vssd1 vssd1 vccd1 vccd1 _06359_ sky130_fd_sc_hd__a211o_1
XANTENNA__08473__A1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13943__113 clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 net1582 sky130_fd_sc_hd__inv_2
XANTENNA__09670__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08345__X _03984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xteam_08_1416 vssd1 vssd1 vccd1 vccd1 team_08_1416/HI gpio_oeb[2] sky130_fd_sc_hd__conb_1
Xteam_08_1427 vssd1 vssd1 vccd1 vccd1 team_08_1427/HI gpio_oeb[13] sky130_fd_sc_hd__conb_1
XFILLER_174_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16253_ clknet_leaf_60_clk _02463_ net1139 vssd1 vssd1 vccd1 vccd1 top.CPU.control_unit.instruction\[29\]
+ sky130_fd_sc_hd__dfrtp_2
Xteam_08_1438 vssd1 vssd1 vccd1 vccd1 team_08_1438/HI gpio_out[23] sky130_fd_sc_hd__conb_1
XFILLER_173_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13465_ net1396 net873 _02910_ net418 vssd1 vssd1 vccd1 vccd1 _02954_ sky130_fd_sc_hd__a31o_1
Xteam_08_1449 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] team_08_1449/LO sky130_fd_sc_hd__conb_1
X_10677_ net3623 net225 net311 _06293_ vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__a22o_1
XFILLER_139_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15204_ net1538 _01414_ net1211 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_93_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12416_ top.CPU.addressnew\[7\] top.CPU.addressnew\[19\] top.CPU.addressnew\[18\]
+ top.CPU.addressnew\[4\] vssd1 vssd1 vccd1 vccd1 _06942_ sky130_fd_sc_hd__or4b_1
XFILLER_173_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16184_ net2518 _02394_ net1149 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[984\]
+ sky130_fd_sc_hd__dfrtp_1
X_13396_ net890 _02914_ vssd1 vssd1 vccd1 vccd1 _02915_ sky130_fd_sc_hd__and2_1
XANTENNA__12027__B _06781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14078__248 clknet_leaf_153_clk vssd1 vssd1 vccd1 vccd1 net1717 sky130_fd_sc_hd__inv_2
X_15135_ clknet_leaf_47_clk _01345_ net1130 vssd1 vssd1 vccd1 vccd1 top.I2C.data_out\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_127_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08776__A2 net1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12347_ net1339 top.I2C.output_state\[16\] net3234 vssd1 vssd1 vccd1 vccd1 _06896_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_127_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07984__B1 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15066_ clknet_leaf_52_clk _00045_ net1133 vssd1 vssd1 vccd1 vccd1 top.I2C.output_state\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_142_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12278_ net2674 _06887_ vssd1 vssd1 vccd1 vccd1 _06888_ sky130_fd_sc_hd__nand2_1
XFILLER_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08528__A2 net1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14119__289 clknet_leaf_184_clk vssd1 vssd1 vccd1 vccd1 net1758 sky130_fd_sc_hd__inv_2
X_11229_ net3451 net296 _06669_ net319 vssd1 vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__a22o_1
XANTENNA__08933__C1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16377__RESET_B net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12088__A2 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15968_ net2302 _02178_ net1093 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[768\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10099__A1 _03407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14919_ clknet_leaf_76_clk _01165_ net1155 vssd1 vssd1 vccd1 vccd1 top.CPU.alu.program_counter\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_19_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15899_ net2233 _02109_ net1214 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[699\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11835__A2 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08440_ top.CPU.registers.data\[849\] net1326 net857 top.CPU.registers.data\[881\]
+ net750 vssd1 vssd1 vccd1 vccd1 _04079_ sky130_fd_sc_hd__a221o_1
XANTENNA__08700__A2 net1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_886 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13851__21 clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 net1490 sky130_fd_sc_hd__inv_2
X_14776__946 clknet_leaf_160_clk vssd1 vssd1 vccd1 vccd1 net2415 sky130_fd_sc_hd__inv_2
XANTENNA__11048__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08371_ top.CPU.registers.data\[50\] top.CPU.registers.data\[18\] net818 vssd1 vssd1
+ vccd1 vccd1 _04010_ sky130_fd_sc_hd__mux2_1
XANTENNA__11106__B net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11821__S net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09110__C1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09661__B1 _03650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14520__690 clknet_leaf_167_clk vssd1 vssd1 vccd1 vccd1 net2159 sky130_fd_sc_hd__inv_2
X_14817__987 clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 net2456 sky130_fd_sc_hd__inv_2
XFILLER_31_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11122__A net1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08216__A1 _03823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09413__B1 net1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10023__A1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08767__A2 net1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07975__B1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout402 net405 vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08519__A2 _04155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09177__C1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout499_A net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout413 net415 vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__clkbuf_4
X_14853__1023 clknet_leaf_110_clk vssd1 vssd1 vccd1 vccd1 net2492 sky130_fd_sc_hd__inv_2
XFILLER_160_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10025__X _05664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout424 _06756_ vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__buf_6
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout435 _06467_ vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__buf_8
Xfanout446 _05517_ vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08924__C1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input4_A DAT_I[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout457 net463 vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__buf_4
XANTENNA__09192__A2 net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09825_ net803 _05457_ _05463_ vssd1 vssd1 vccd1 vccd1 _05464_ sky130_fd_sc_hd__and3_1
Xfanout468 net470 vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__buf_4
XFILLER_150_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12888__A top.CPU.alu.program_counter\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout479 net482 vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__buf_4
XANTENNA_fanout287_X net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09756_ net751 _05375_ _05376_ net708 vssd1 vssd1 vccd1 vccd1 _05395_ sky130_fd_sc_hd__a31o_1
XANTENNA__12079__A2 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08707_ _04342_ _04345_ net640 vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__a21o_1
XFILLER_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11826__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09687_ top.CPU.registers.data\[473\] net1336 net869 top.CPU.registers.data\[505\]
+ net732 vssd1 vssd1 vccd1 vccd1 _05326_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout454_X net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08152__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout833_A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08638_ top.CPU.registers.data\[78\] net1320 net851 top.CPU.registers.data\[110\]
+ net769 vssd1 vssd1 vccd1 vccd1 _04277_ sky130_fd_sc_hd__a221o_1
XFILLER_55_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10695__X _06311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08569_ top.CPU.registers.data_out_r1_prev\[15\] net871 _04204_ _04207_ net691 vssd1
+ vssd1 vccd1 vccd1 _04208_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout621_X net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1363_X net1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout719_X net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10600_ net400 _06219_ vssd1 vssd1 vccd1 vccd1 _06220_ sky130_fd_sc_hd__nand2_1
XANTENNA__13512__A _04254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08455__A1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11580_ net493 net477 _06692_ net249 net2633 vssd1 vssd1 vccd1 vccd1 _01961_ sky130_fd_sc_hd__a32o_1
XFILLER_70_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10531_ _04330_ _06153_ vssd1 vssd1 vccd1 vccd1 _06154_ sky130_fd_sc_hd__or2_1
XFILLER_128_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11032__A _03180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13250_ net3903 _02805_ _02809_ _02803_ vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__a22o_1
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10462_ _04021_ net373 _05729_ vssd1 vssd1 vccd1 vccd1 _06088_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09404__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout990_X net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13658__S net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12201_ _06541_ _06796_ _06867_ net169 net2943 vssd1 vssd1 vccd1 vccd1 _01461_ sky130_fd_sc_hd__a32o_1
XFILLER_170_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13181_ top.I2C.within_byte_counter_writing\[0\] top.I2C.which_data_address\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__or2_1
XANTENNA__12415__X _06941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10393_ _05975_ _06021_ net308 vssd1 vssd1 vccd1 vccd1 _06022_ sky130_fd_sc_hd__mux2_1
XFILLER_136_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10565__A2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11762__A1 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12132_ top.CPU.registers.data\[86\] net655 _06749_ vssd1 vssd1 vccd1 vccd1 _06834_
+ sky130_fd_sc_hd__o21a_1
XFILLER_124_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08341__A net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09168__C1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11178__S net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10082__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12063_ net4001 net656 _06800_ vssd1 vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__o21a_1
XFILLER_2_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08915__C1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11014_ net3238 net217 _06563_ net313 vssd1 vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__a22o_1
XFILLER_77_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout980 net985 vssd1 vssd1 vccd1 vccd1 net980 sky130_fd_sc_hd__buf_2
XANTENNA__08930__A2 net1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout991 net994 vssd1 vssd1 vccd1 vccd1 net991 sky130_fd_sc_hd__buf_2
X_15822_ net2156 _02032_ net1106 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[622\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08487__S net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10589__Y _06210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13267__B2 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14463__633 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 net2102 sky130_fd_sc_hd__inv_2
X_15753_ net2087 _01963_ net1060 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[553\]
+ sky130_fd_sc_hd__dfrtp_1
X_12965_ net1342 _07402_ vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__nor2_1
XANTENNA__09340__C1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11916_ net3465 net187 net345 _06151_ vssd1 vssd1 vccd1 vccd1 _01650_ sky130_fd_sc_hd__a22o_1
X_15684_ net2018 _01894_ net1212 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[484\]
+ sky130_fd_sc_hd__dfrtp_1
X_12896_ _07339_ _07340_ vssd1 vssd1 vccd1 vccd1 _07341_ sky130_fd_sc_hd__nand2b_1
XFILLER_127_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14504__674 clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 net2143 sky130_fd_sc_hd__inv_2
X_11847_ net468 _06678_ net237 net153 net2656 vssd1 vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__a32o_1
XFILLER_33_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11778_ _06621_ net199 net160 net3637 vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__a22o_1
XANTENNA__10789__C1 _05664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10765__B net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16305_ clknet_leaf_83_clk _02514_ net1261 vssd1 vssd1 vccd1 vccd1 top.CPU.data_out\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13517_ _04122_ net584 vssd1 vssd1 vccd1 vccd1 _02979_ sky130_fd_sc_hd__and2_1
XFILLER_119_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10729_ _06294_ _06342_ net307 vssd1 vssd1 vccd1 vccd1 _06343_ sky130_fd_sc_hd__mux2_1
X_16236_ clknet_leaf_45_clk _02446_ net1138 vssd1 vssd1 vccd1 vccd1 top.CPU.control_unit.instruction\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13448_ net3629 _02945_ net123 vssd1 vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__mux2_1
Xclkload12 clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clkload12/Y sky130_fd_sc_hd__inv_12
Xclkload23 clknet_leaf_199_clk vssd1 vssd1 vccd1 vccd1 clkload23/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__10005__A1 _04020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload34 clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 clkload34/Y sky130_fd_sc_hd__inv_4
Xclkload45 clknet_leaf_189_clk vssd1 vssd1 vccd1 vccd1 clkload45/Y sky130_fd_sc_hd__inv_12
XANTENNA_clkbuf_leaf_173_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16167_ net2501 _02377_ net1198 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[967\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload56 clknet_leaf_176_clk vssd1 vssd1 vccd1 vccd1 clkload56/Y sky130_fd_sc_hd__clkinv_16
X_13379_ _02830_ _02902_ vssd1 vssd1 vccd1 vccd1 _02903_ sky130_fd_sc_hd__nor2_1
Xclkload67 clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 clkload67/Y sky130_fd_sc_hd__inv_16
XANTENNA__10781__A net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload78 clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 clkload78/Y sky130_fd_sc_hd__inv_6
XFILLER_55_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07957__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15118_ net1500 _01331_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r2_prev\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload89 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 clkload89/Y sky130_fd_sc_hd__inv_6
XANTENNA_clkbuf_leaf_53_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16098_ net2432 _02308_ net1171 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[898\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_142_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16241__Q top.CPU.control_unit.instruction\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07940_ _03544_ _03577_ vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__nand2_2
X_15049_ clknet_leaf_92_clk _01294_ net1268 vssd1 vssd1 vccd1 vccd1 top.SPI.command\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10308__A2 _05939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07709__B1 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_188_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12702__B1 top.CPU.alu.program_counter\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07871_ _03509_ vssd1 vssd1 vccd1 vccd1 _03510_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_143_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09610_ net691 _05247_ _05248_ vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_3_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_68_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08921__A2 net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09541_ top.CPU.registers.data\[65\] net1334 net866 top.CPU.registers.data\[97\]
+ net780 vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_111_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09331__C1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09472_ net707 _05109_ _05110_ _05108_ vssd1 vssd1 vccd1 vccd1 _05111_ sky130_fd_sc_hd__a31o_1
XFILLER_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10492__A1 _03315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08423_ top.CPU.registers.data\[337\] net1326 net857 top.CPU.registers.data\[369\]
+ net774 vssd1 vssd1 vccd1 vccd1 _04062_ sky130_fd_sc_hd__a221o_1
XFILLER_52_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10956__A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout247_A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_126_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08354_ top.CPU.registers.data\[658\] net1320 net851 top.CPU.registers.data\[690\]
+ net720 vssd1 vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__a221o_1
XANTENNA__13430__A1 _02861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08988__A2 net1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload6 clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clkload6/Y sky130_fd_sc_hd__clkinv_8
X_08285_ _03859_ _03922_ vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout414_A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10795__A2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13478__S net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09398__C1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout202_X net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1323_A _03109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11744__A1 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07948__B1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08161__A net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout783_A net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1208 net1209 vssd1 vssd1 vccd1 vccd1 net1208 sky130_fd_sc_hd__clkbuf_4
Xfanout210 net211 vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1111_X net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1219 net1226 vssd1 vssd1 vccd1 vccd1 net1219 sky130_fd_sc_hd__clkbuf_4
Xfanout221 _06469_ vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__clkbuf_4
Xfanout232 _06772_ vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__clkbuf_4
XFILLER_115_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14150__320 clknet_leaf_123_clk vssd1 vssd1 vccd1 vccd1 net1789 sky130_fd_sc_hd__inv_2
Xfanout243 _06750_ vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout950_A net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout571_X net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout254 _06728_ vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10704__C1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14447__617 clknet_leaf_178_clk vssd1 vssd1 vccd1 vccd1 net2086 sky130_fd_sc_hd__inv_2
Xfanout265 net266 vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout669_X net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout276 net279 vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__buf_4
X_09808_ net711 _05446_ vssd1 vssd1 vccd1 vccd1 _05447_ sky130_fd_sc_hd__or2_1
XANTENNA__08912__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout287 net288 vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__clkbuf_8
Xfanout298 _06645_ vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09704__B net1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09739_ top.CPU.registers.data\[91\] net1331 net859 top.CPU.registers.data\[123\]
+ net775 vssd1 vssd1 vccd1 vccd1 _05378_ sky130_fd_sc_hd__a221o_1
XFILLER_131_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout836_X net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11397__D_N net1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09322__C1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12750_ top.CPU.alu.program_counter\[11\] _07191_ vssd1 vssd1 vccd1 vccd1 _07209_
+ sky130_fd_sc_hd__nor2_1
XFILLER_83_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11701_ _06533_ net209 net422 net3791 vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__a22o_1
X_12681_ top.CPU.alu.program_counter\[4\] _03118_ _07145_ _07146_ vssd1 vssd1 vccd1
+ vccd1 _01167_ sky130_fd_sc_hd__a22o_1
XANTENNA__11680__B1 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07884__C1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10866__A _05692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11461__S net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11632_ _05811_ net201 net424 net3619 vssd1 vssd1 vccd1 vccd1 _01919_ sky130_fd_sc_hd__a22o_1
XFILLER_168_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_139_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16326__Q top.CPU.addressnew\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08979__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11563_ net3198 net247 _06742_ net485 vssd1 vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__a22o_1
X_13302_ top.CPU.addressnew\[2\] top.CPU.addressnew\[17\] top.CPU.done top.CPU.addressnew\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02845_ sky130_fd_sc_hd__and4b_1
X_10514_ _05944_ _06137_ net403 vssd1 vssd1 vccd1 vccd1 _06138_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_21_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11494_ _06625_ net258 net254 net3663 vssd1 vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__a22o_1
XANTENNA__09389__C1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16021_ net2355 _02231_ net1217 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[821\]
+ sky130_fd_sc_hd__dfrtp_1
X_13233_ _02787_ _02793_ vssd1 vssd1 vccd1 vccd1 _02800_ sky130_fd_sc_hd__nor2_1
X_10445_ net407 _06071_ vssd1 vssd1 vccd1 vccd1 _06072_ sky130_fd_sc_hd__nor2_1
XFILLER_155_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12292__S net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13164_ _06950_ _03123_ top.I2C.initiate_read_bit vssd1 vssd1 vccd1 vccd1 _02751_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__08600__A1 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10376_ net415 _06005_ vssd1 vssd1 vccd1 vccd1 _06006_ sky130_fd_sc_hd__nor2_1
XFILLER_2_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12115_ net655 _06473_ _06749_ net175 net2924 vssd1 vssd1 vccd1 vccd1 _01505_ sky130_fd_sc_hd__a32o_1
XFILLER_3_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13095_ top.CPU.data_out\[30\] net3409 net559 vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__mux2_1
XANTENNA__13488__A1 _05084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_15_0_clk_X clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12046_ net147 net3477 net151 vssd1 vssd1 vccd1 vccd1 _01542_ sky130_fd_sc_hd__mux2_1
XANTENNA__11499__B1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12160__A1 _06311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08364__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09561__C1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10540__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15805_ net2139 _02015_ net1113 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[605\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_18_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12948_ top.CPU.alu.program_counter\[30\] _07381_ vssd1 vssd1 vccd1 vccd1 _07388_
+ sky130_fd_sc_hd__nor2_1
X_15736_ net2070 _01946_ net1102 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[536\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13660__A1 _03152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11671__B1 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07875__C1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12879_ top.CPU.alu.program_counter\[23\] _07325_ net1359 vssd1 vssd1 vccd1 vccd1
+ _01186_ sky130_fd_sc_hd__mux2_1
X_15667_ net2001 _01877_ net1178 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[467\]
+ sky130_fd_sc_hd__dfrtp_1
X_14852__1022 clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 net2491 sky130_fd_sc_hd__inv_2
X_15598_ net1932 _01808_ net1107 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[398\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07890__A2 net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11423__B1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09776__S net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08070_ top.CPU.registers.data\[276\] net979 vssd1 vssd1 vccd1 vccd1 _03709_ sky130_fd_sc_hd__nand2_1
Xclkload101 clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 clkload101/Y sky130_fd_sc_hd__inv_8
X_14591__761 clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 net2230 sky130_fd_sc_hd__inv_2
Xclkload112 clknet_leaf_158_clk vssd1 vssd1 vccd1 vccd1 clkload112/Y sky130_fd_sc_hd__inv_6
Xclkload123 clknet_leaf_121_clk vssd1 vssd1 vccd1 vccd1 clkload123/Y sky130_fd_sc_hd__clkinv_8
Xclkload134 clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 clkload134/Y sky130_fd_sc_hd__inv_12
X_16219_ net2553 _02429_ net1213 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[1019\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload145 clknet_leaf_163_clk vssd1 vssd1 vccd1 vccd1 clkload145/Y sky130_fd_sc_hd__clkinv_8
XFILLER_161_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload156 clknet_leaf_139_clk vssd1 vssd1 vccd1 vccd1 clkload156/Y sky130_fd_sc_hd__inv_8
Xclkload167 clknet_leaf_81_clk vssd1 vssd1 vccd1 vccd1 clkload167/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__07527__A_N _03152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload178 clknet_leaf_126_clk vssd1 vssd1 vccd1 vccd1 clkload178/Y sky130_fd_sc_hd__inv_4
Xclkload189 clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 clkload189/Y sky130_fd_sc_hd__inv_8
XFILLER_143_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08052__C1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14134__304 clknet_leaf_175_clk vssd1 vssd1 vccd1 vccd1 net1773 sky130_fd_sc_hd__inv_2
X_08972_ top.CPU.registers.data\[169\] top.CPU.registers.data\[137\] net806 vssd1
+ vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__mux2_1
XFILLER_103_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10016__A net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13479__A1 net1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09147__A2 net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07923_ top.CPU.registers.data\[828\] top.CPU.registers.data\[796\] net996 vssd1
+ vssd1 vccd1 vccd1 _03562_ sky130_fd_sc_hd__mux2_1
Xhold18 top.CPU.registers.data_out_r2_prev\[6\] vssd1 vssd1 vccd1 vccd1 net2575 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 top.CPU.registers.data_out_r1_prev\[5\] vssd1 vssd1 vccd1 vccd1 net2586 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_60_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout197_A net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13839__9 clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 net1478 sky130_fd_sc_hd__inv_2
XFILLER_60_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07854_ top.CPU.registers.data\[861\] net1288 net1007 top.CPU.registers.data\[893\]
+ net931 vssd1 vssd1 vccd1 vccd1 _03493_ sky130_fd_sc_hd__a221o_1
XFILLER_72_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07785_ net944 _03422_ _03423_ net614 vssd1 vssd1 vccd1 vccd1 _03424_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout364_A net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09304__C1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09524_ top.CPU.registers.data\[833\] net1335 net868 top.CPU.registers.data\[865\]
+ net757 vssd1 vssd1 vccd1 vccd1 _05163_ sky130_fd_sc_hd__a221o_1
XFILLER_24_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09455_ top.CPU.registers.data\[66\] net1324 net855 top.CPU.registers.data\[98\]
+ net773 vssd1 vssd1 vccd1 vccd1 _05094_ sky130_fd_sc_hd__a221o_1
XANTENNA__10686__A net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout531_A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout152_X net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1273_A net1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout629_A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08406_ top.CPU.registers.data\[466\] net1291 net1012 top.CPU.registers.data\[498\]
+ net908 vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__a221o_1
X_09386_ top.CPU.registers.data\[291\] top.CPU.registers.data\[259\] net828 vssd1
+ vssd1 vccd1 vccd1 _05025_ sky130_fd_sc_hd__mux2_1
XANTENNA__12206__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07881__A2 net1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_49_Left_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11414__B1 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08337_ net955 _03975_ _03972_ net612 vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_173_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout417_X net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08268_ net681 _03905_ _03906_ vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__and3_1
XFILLER_119_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout998_A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08199_ top.CPU.registers.data_out_r2_prev\[23\] net687 net620 _03831_ _03837_ vssd1
+ vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__o2111a_1
XANTENNA_fanout1326_X net1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10230_ net395 _05649_ _05864_ net408 vssd1 vssd1 vccd1 vccd1 _05865_ sky130_fd_sc_hd__a211o_1
XFILLER_105_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout786_X net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11193__A2 _06500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10161_ net550 _05513_ _05796_ _05797_ vssd1 vssd1 vccd1 vccd1 _05798_ sky130_fd_sc_hd__o211a_1
XANTENNA__12840__S net1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1005 net1032 vssd1 vssd1 vccd1 vccd1 net1005 sky130_fd_sc_hd__clkbuf_2
Xfanout1016 net1017 vssd1 vssd1 vccd1 vccd1 net1016 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_58_Left_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13508__Y _02974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1027 net1028 vssd1 vssd1 vccd1 vccd1 net1027 sky130_fd_sc_hd__buf_2
X_10092_ _03684_ net373 _05729_ vssd1 vssd1 vccd1 vccd1 _05730_ sky130_fd_sc_hd__a21o_1
Xfanout1038 _03178_ vssd1 vssd1 vccd1 vccd1 net1038 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout953_X net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1049 _03093_ vssd1 vssd1 vccd1 vccd1 net1049 sky130_fd_sc_hd__buf_2
XFILLER_59_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09543__C1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12802_ _07237_ _07255_ _07244_ vssd1 vssd1 vccd1 vccd1 _07256_ sky130_fd_sc_hd__o21ba_1
X_13782_ net10 net1051 net886 net4015 vssd1 vssd1 vccd1 vccd1 _02663_ sky130_fd_sc_hd__a22o_1
XANTENNA__08649__A1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10994_ net514 _06213_ net542 vssd1 vssd1 vccd1 vccd1 _06551_ sky130_fd_sc_hd__and3_1
X_12733_ _07191_ _07192_ vssd1 vssd1 vccd1 vccd1 _07193_ sky130_fd_sc_hd__nor2_1
XFILLER_16_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15521_ net1855 _01731_ net1225 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[321\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10456__B2 top.CPU.handler.toreg\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11653__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07857__C1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_67_Left_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15452_ net1786 _01662_ net1195 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[252\]
+ sky130_fd_sc_hd__dfrtp_1
X_12664_ top.CPU.alu.program_counter\[3\] _05021_ vssd1 vssd1 vccd1 vccd1 _07131_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_61_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14575__745 clknet_leaf_178_clk vssd1 vssd1 vccd1 vccd1 net2214 sky130_fd_sc_hd__inv_2
X_11615_ _06230_ net3417 net212 vssd1 vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__mux2_1
XANTENNA__11405__B1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15383_ net1717 _01593_ net1180 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[183\]
+ sky130_fd_sc_hd__dfrtp_1
X_12595_ top.SPI.command\[0\] top.SPI.command\[4\] vssd1 vssd1 vccd1 vccd1 _07096_
+ sky130_fd_sc_hd__or2_1
XFILLER_129_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09596__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11546_ net3475 net253 _06734_ _06520_ vssd1 vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__a22o_1
XANTENNA__08821__A1 _04459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14616__786 clknet_leaf_160_clk vssd1 vssd1 vccd1 vccd1 net2255 sky130_fd_sc_hd__inv_2
X_11477_ net3703 net254 _06729_ net484 vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__a22o_1
XANTENNA__14926__RESET_B net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16004_ net2338 _02214_ net1186 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[804\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11220__A net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13216_ net893 top.I2C.data_out\[23\] _02789_ vssd1 vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10428_ top.CPU.fetch.current_ra\[20\] net1040 net881 top.CPU.handler.toreg\[20\]
+ _06055_ vssd1 vssd1 vccd1 vccd1 _06056_ sky130_fd_sc_hd__a221o_4
XPHY_EDGE_ROW_164_Right_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_76_Left_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13147_ net126 _02738_ net1359 vssd1 vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10392__A0 _03755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10359_ net600 _05988_ _05989_ vssd1 vssd1 vccd1 vccd1 _05990_ sky130_fd_sc_hd__o21ai_4
XFILLER_3_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10931__A2 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13078_ top.CPU.data_out\[13\] net3159 net558 vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__mux2_1
XFILLER_111_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09534__C1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12029_ net362 _06724_ _06791_ _06790_ vssd1 vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__a31o_1
XANTENNA__08888__A1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11892__A0 _06373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07570_ net1047 _03163_ net1038 _03111_ vssd1 vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__a31o_1
XANTENNA__09837__B1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08675__S net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_85_Left_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11644__B1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15719_ net2053 _01929_ net1201 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[519\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07848__C1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09240_ top.CPU.registers.data\[741\] net1387 net809 top.CPU.registers.data\[709\]
+ net715 vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__a221o_1
XANTENNA__07863__A2 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13397__A0 top.CPU.control_unit.instruction\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11114__B net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09171_ net789 _04809_ vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__or2_1
XANTENNA__09065__A1 net1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08122_ top.CPU.registers.data\[949\] top.CPU.registers.data\[917\] top.CPU.registers.data\[821\]
+ top.CPU.registers.data\[789\] net992 net917 vssd1 vssd1 vccd1 vccd1 _03761_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_116_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10953__B net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08053_ net674 _03690_ _03691_ net604 vssd1 vssd1 vccd1 vccd1 _03692_ sky130_fd_sc_hd__a31o_1
XFILLER_147_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11130__A net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08025__C1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_131_Right_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08576__B1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09773__C1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1021_A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10922__A2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08955_ top.CPU.registers.data_out_r2_prev\[10\] _04593_ net686 vssd1 vssd1 vccd1
+ vccd1 _04594_ sky130_fd_sc_hd__mux2_1
XFILLER_102_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08328__B1 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout481_A net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07906_ top.CPU.registers.data\[60\] net1025 net944 vssd1 vssd1 vccd1 vccd1 _03545_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__09525__C1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10033__X _05672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08886_ top.CPU.registers.data\[971\] net1309 net840 top.CPU.registers.data\[1003\]
+ net764 vssd1 vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__a221o_1
XANTENNA__10135__B1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07837_ top.CPU.alu.program_counter\[29\] _03474_ net1037 vssd1 vssd1 vccd1 vccd1
+ _03476_ sky130_fd_sc_hd__mux2_4
XFILLER_84_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11883__B1 net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1390_A net1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout367_X net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout746_A net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09828__A0 top.CPU.alu.program_counter\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07768_ net1036 _03405_ _03376_ vssd1 vssd1 vccd1 vccd1 _03407_ sky130_fd_sc_hd__a21oi_4
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09507_ net629 _05141_ _05142_ net615 vssd1 vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__a31o_1
XFILLER_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11635__B1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13504__B _02966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14262__432 clknet_leaf_182_clk vssd1 vssd1 vccd1 vccd1 net1901 sky130_fd_sc_hd__inv_2
XFILLER_72_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout534_X net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout913_A net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07699_ top.CPU.registers.data\[543\] net1030 _03335_ net959 vssd1 vssd1 vccd1 vccd1
+ _03338_ sky130_fd_sc_hd__o211a_1
XFILLER_169_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1276_X net1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14559__729 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 net2198 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_23_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09438_ top.CPU.registers.data\[962\] net1294 net1015 top.CPU.registers.data\[994\]
+ net911 vssd1 vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__a221o_1
XFILLER_24_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09369_ top.CPU.registers.data\[675\] top.CPU.registers.data\[643\] top.CPU.registers.data\[547\]
+ top.CPU.registers.data\[515\] net990 net915 vssd1 vssd1 vccd1 vccd1 _05008_ sky130_fd_sc_hd__mux4_1
XANTENNA__09056__A1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout701_X net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14303__473 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 net1942 sky130_fd_sc_hd__inv_2
X_11400_ _06529_ net278 net268 net3386 vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__a22o_1
X_12380_ top.CPU.addressnew\[21\] top.CPU.addressnew\[20\] top.CPU.addressnew\[23\]
+ top.CPU.addressnew\[22\] vssd1 vssd1 vccd1 vccd1 _06918_ sky130_fd_sc_hd__or4_2
XANTENNA__08264__C1 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10863__B net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10610__A1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11331_ _03189_ net461 vssd1 vssd1 vccd1 vccd1 _06713_ sky130_fd_sc_hd__nor2_2
XANTENNA__09359__A2 net1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11262_ net480 net457 _06687_ net293 net2682 vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__a32o_1
XANTENNA__08016__C1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13001_ net3852 _07427_ _07428_ _06946_ vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__o211a_1
XANTENNA__08567__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13560__B1 _03002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09764__C1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10213_ net575 net519 net442 _05848_ vssd1 vssd1 vccd1 vccd1 _05849_ sky130_fd_sc_hd__and4_1
XANTENNA__12423__X _06948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11193_ net486 _06500_ _06648_ net298 net3000 vssd1 vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_37_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10144_ _05779_ _05780_ net387 vssd1 vssd1 vccd1 vccd1 _05781_ sky130_fd_sc_hd__mux2_1
XFILLER_0_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12115__A1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14851__1021 clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 net2490 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_54_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14952_ clknet_leaf_53_clk _01198_ net1133 vssd1 vssd1 vccd1 vccd1 top.I2C.bit_timer_counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_130_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10075_ _04567_ _04634_ net380 vssd1 vssd1 vccd1 vccd1 _05713_ sky130_fd_sc_hd__mux2_1
XFILLER_153_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10103__B _05664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16622_ top.I2C.sda_out vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__clkbuf_1
XFILLER_35_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09819__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16553_ clknet_leaf_64_clk net2607 net1163 vssd1 vssd1 vccd1 vccd1 top.mmio.m2 sky130_fd_sc_hd__dfrtp_1
X_13765_ net2 net1049 net884 net3700 vssd1 vssd1 vccd1 vccd1 _02646_ sky130_fd_sc_hd__o22a_1
XFILLER_44_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11626__B1 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10977_ net3594 net217 _06540_ net314 vssd1 vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__a22o_1
XANTENNA__11215__A net1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15504_ net1838 _01714_ net1194 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[304\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_149_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12716_ _07176_ _07177_ vssd1 vssd1 vccd1 vccd1 _07178_ sky130_fd_sc_hd__nand2_1
XFILLER_31_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13696_ net3708 _03049_ vssd1 vssd1 vccd1 vccd1 _03053_ sky130_fd_sc_hd__nor2_1
X_16484_ clknet_leaf_41_clk _02646_ net1116 vssd1 vssd1 vccd1 vccd1 top.mmio.mem_data_i\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12647_ net1411 net1341 net2973 vssd1 vssd1 vccd1 vccd1 _00018_ sky130_fd_sc_hd__and3_1
XFILLER_129_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15435_ net1769 _01645_ net1057 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[235\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09598__A2 net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12051__B1 _06781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08255__C1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15366_ net1700 _01576_ net1081 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[166\]
+ sky130_fd_sc_hd__dfrtp_1
X_12578_ _03101_ _07053_ _07055_ _07082_ vssd1 vssd1 vccd1 vccd1 _07083_ sky130_fd_sc_hd__o31a_1
XFILLER_157_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_96_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11529_ _06654_ net258 net251 net3632 vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__a22o_1
X_15297_ net1631 _01507_ net1225 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[97\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold307 top.CPU.registers.data\[675\] vssd1 vssd1 vccd1 vccd1 net2864 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold318 top.CPU.registers.data\[575\] vssd1 vssd1 vccd1 vccd1 net2875 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold329 top.CPU.registers.data\[975\] vssd1 vssd1 vccd1 vccd1 net2886 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13551__A0 top.CPU.alu.program_counter\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout809 net812 vssd1 vssd1 vccd1 vccd1 net809 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10904__A2 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09770__A2 net1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08740_ top.CPU.registers.data\[973\] net1371 net968 top.CPU.registers.data\[1005\]
+ net1364 vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__o221a_1
Xhold1007 top.CPU.registers.data\[248\] vssd1 vssd1 vccd1 vccd1 net3564 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1018 top.CPU.registers.data\[875\] vssd1 vssd1 vccd1 vccd1 net3575 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1029 top.CPU.registers.data\[438\] vssd1 vssd1 vccd1 vccd1 net3586 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout1380 net1385 vssd1 vssd1 vccd1 vccd1 net1380 sky130_fd_sc_hd__clkbuf_4
XFILLER_38_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1391 net1392 vssd1 vssd1 vccd1 vccd1 net1391 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11865__B1 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08671_ top.CPU.registers.data\[974\] net1378 net982 top.CPU.registers.data\[1006\]
+ net1365 vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__o221a_1
XFILLER_27_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11824__S net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07622_ _03258_ _03260_ _03247_ _03256_ vssd1 vssd1 vccd1 vccd1 _03261_ sky130_fd_sc_hd__a211oi_2
XTAP_TAPCELL_ROW_109_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14246__416 clknet_leaf_134_clk vssd1 vssd1 vccd1 vccd1 net1885 sky130_fd_sc_hd__inv_2
XFILLER_53_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10948__B _03170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11617__A0 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07553_ net563 _03183_ vssd1 vssd1 vccd1 vccd1 _03192_ sky130_fd_sc_hd__or2_1
XANTENNA__10300__Y _05933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07484_ top.I2C.within_byte_counter_writing\[2\] vssd1 vssd1 vccd1 vccd1 _03124_
+ sky130_fd_sc_hd__inv_2
XANTENNA__08494__C1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_153_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09223_ _04859_ _04860_ vssd1 vssd1 vccd1 vccd1 _04862_ sky130_fd_sc_hd__nand2_2
XFILLER_166_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09038__A1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09089__X _04728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1069_A net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09154_ top.CPU.control_unit.instruction\[27\] _04596_ _04597_ vssd1 vssd1 vccd1
+ vccd1 _04793_ sky130_fd_sc_hd__o21a_2
XANTENNA__12042__B1 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11396__A2 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08105_ top.CPU.registers.data\[341\] net1330 net861 top.CPU.registers.data\[373\]
+ net776 vssd1 vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_4_3_0_clk_X clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13790__B1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09085_ net1366 _04716_ _04715_ top.CPU.control_unit.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 _04724_ sky130_fd_sc_hd__o211a_1
XANTENNA__08261__A2 net1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1236_A net1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08036_ net743 _03673_ _03674_ net692 vssd1 vssd1 vccd1 vccd1 _03675_ sky130_fd_sc_hd__o211a_1
Xhold830 top.CPU.registers.data\[363\] vssd1 vssd1 vccd1 vccd1 net3387 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold841 top.CPU.registers.data\[241\] vssd1 vssd1 vccd1 vccd1 net3398 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11148__A2 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold852 top.SPI.parameters\[30\] vssd1 vssd1 vccd1 vccd1 net3409 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13486__S net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout696_A net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13542__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09746__C1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold863 top.CPU.registers.data\[401\] vssd1 vssd1 vccd1 vccd1 net3420 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold874 top.CPU.registers.data\[506\] vssd1 vssd1 vccd1 vccd1 net3431 sky130_fd_sc_hd__dlygate4sd3_1
Xhold885 top.CPU.registers.data\[243\] vssd1 vssd1 vccd1 vccd1 net3442 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1403_A net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold896 top.CPU.registers.data\[529\] vssd1 vssd1 vccd1 vccd1 net3453 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_67_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09987_ _04829_ net372 vssd1 vssd1 vccd1 vccd1 _05626_ sky130_fd_sc_hd__nor2_1
XFILLER_114_1008 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout863_A net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout484_X net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08938_ top.CPU.registers.data\[202\] net1374 net972 top.CPU.registers.data\[234\]
+ net928 vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_129_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10659__A1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout651_X net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08869_ top.CPU.registers.data\[171\] top.CPU.registers.data\[139\] net808 vssd1
+ vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__mux2_1
XANTENNA__11856__B1 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1393_X net1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout749_X net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11320__A2 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10900_ net485 net459 _06493_ net221 net3074 vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__a32o_1
X_11880_ net139 net3361 net188 vssd1 vssd1 vccd1 vccd1 _01683_ sky130_fd_sc_hd__mux2_1
XFILLER_26_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11608__A0 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10831_ net381 _06394_ vssd1 vssd1 vccd1 vccd1 _06440_ sky130_fd_sc_hd__nand2_1
XFILLER_16_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09277__A1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout916_X net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13550_ top.CPU.addressnew\[0\] _02996_ net580 vssd1 vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__mux2_1
XFILLER_16_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10762_ net572 net514 _06374_ vssd1 vssd1 vccd1 vccd1 _06375_ sky130_fd_sc_hd__and3_1
XANTENNA__11084__B2 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1006 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12501_ _04890_ _04918_ vssd1 vssd1 vccd1 vccd1 _07010_ sky130_fd_sc_hd__nor2_1
XANTENNA__07800__X _03439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13481_ net1396 net873 _02932_ net418 vssd1 vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__a31o_1
X_10693_ net511 _06308_ _06307_ vssd1 vssd1 vccd1 vccd1 _06309_ sky130_fd_sc_hd__a21oi_4
XANTENNA__10874__A net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08615__Y _04254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15220_ net1554 _01430_ net1080 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_12432_ net898 _06952_ vssd1 vssd1 vccd1 vccd1 _00057_ sky130_fd_sc_hd__nor2_1
XFILLER_139_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12033__B1 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08237__C1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10593__B net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11387__A2 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08788__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15151_ clknet_leaf_42_clk _01361_ net1117 vssd1 vssd1 vccd1 vccd1 top.I2C.data_out\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_166_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12363_ top.I2C.output_state\[2\] net1054 _06902_ _06905_ vssd1 vssd1 vccd1 vccd1
+ _00060_ sky130_fd_sc_hd__a22o_1
XANTENNA__10595__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11314_ net3083 net290 net358 _06230_ vssd1 vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__a22o_1
X_15082_ clknet_leaf_51_clk _00059_ net1134 vssd1 vssd1 vccd1 vccd1 top.I2C.output_state\[28\]
+ sky130_fd_sc_hd__dfrtp_4
X_13927__97 clknet_leaf_159_clk vssd1 vssd1 vccd1 vccd1 net1566 sky130_fd_sc_hd__inv_2
X_12294_ net2629 _04361_ net1076 vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__mux2_1
XANTENNA__11139__A2 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14390__560 clknet_leaf_182_clk vssd1 vssd1 vccd1 vccd1 net2029 sky130_fd_sc_hd__inv_2
XANTENNA__12336__A1 _04951_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09737__C1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11245_ net492 net468 _06677_ net296 net2641 vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_91_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09201__A1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14687__857 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 net2326 sky130_fd_sc_hd__inv_2
XFILLER_106_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10898__A1 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11176_ net3840 net300 _06649_ net495 vssd1 vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07763__A1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10127_ _05617_ _05722_ _05764_ vssd1 vssd1 vccd1 vccd1 _05765_ sky130_fd_sc_hd__a21bo_1
XFILLER_110_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10114__A net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15377__RESET_B net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14728__898 clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 net2367 sky130_fd_sc_hd__inv_2
X_15984_ net2318 _02194_ net1155 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[784\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09504__A2 net1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14935_ clknet_leaf_70_clk _01181_ net1169 vssd1 vssd1 vccd1 vccd1 top.CPU.alu.program_counter\[18\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_57_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10058_ net563 _03183_ _03185_ vssd1 vssd1 vccd1 vccd1 _05696_ sky130_fd_sc_hd__and3_2
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11847__B1 net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08712__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13817_ net2861 net335 net328 top.CPU.data_out\[19\] vssd1 vssd1 vccd1 vccd1 _02697_
+ sky130_fd_sc_hd__a22o_1
X_16536_ clknet_leaf_99_clk _02698_ net1256 vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__dfrtp_1
X_13748_ top.SPI.timem\[21\] top.SPI.timem\[20\] _03082_ vssd1 vssd1 vccd1 vccd1 _03085_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08476__C1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07710__X _03349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10822__A1 _05672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16467_ clknet_leaf_86_clk _02629_ net1272 vssd1 vssd1 vccd1 vccd1 top.SPI.timem\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10822__B2 _05665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13679_ net2667 net336 vssd1 vssd1 vccd1 vccd1 _02607_ sky130_fd_sc_hd__and2_1
XFILLER_85_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12024__B1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08228__C1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15418_ net1752 _01628_ net1252 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[218\]
+ sky130_fd_sc_hd__dfrtp_1
X_16398_ clknet_leaf_63_clk _00022_ net1162 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11378__A2 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09976__C1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14631__801 clknet_leaf_185_clk vssd1 vssd1 vccd1 vccd1 net2270 sky130_fd_sc_hd__inv_2
X_15349_ net1683 _01559_ net1216 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[149\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10586__B1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold104 top.CPU.registers.data\[298\] vssd1 vssd1 vccd1 vccd1 net2661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 net117 vssd1 vssd1 vccd1 vccd1 net2672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 top.SPI.parameters\[3\] vssd1 vssd1 vccd1 vccd1 net2683 sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 net115 vssd1 vssd1 vccd1 vccd1 net2694 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12327__A1 _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13524__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11819__S _06762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold148 top.CPU.registers.data\[562\] vssd1 vssd1 vccd1 vccd1 net2705 sky130_fd_sc_hd__dlygate4sd3_1
Xhold159 _00033_ vssd1 vssd1 vccd1 vccd1 net2716 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_160_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09910_ net381 _05192_ vssd1 vssd1 vccd1 vccd1 _05549_ sky130_fd_sc_hd__and2b_1
XFILLER_113_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10950__C net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout606 net609 vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__buf_4
Xfanout617 net619 vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__buf_4
X_09841_ net945 _05478_ _05479_ net960 vssd1 vssd1 vccd1 vccd1 _05480_ sky130_fd_sc_hd__o211a_1
XANTENNA__08400__C1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout628 net630 vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__buf_4
XANTENNA_clkload14_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout639 _03225_ vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__buf_4
XFILLER_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11550__A2 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09772_ top.CPU.registers.data\[251\] top.CPU.registers.data\[219\] net990 vssd1
+ vssd1 vccd1 vccd1 _05411_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_146_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13827__B2 top.CPU.data_out\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_13_Left_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08723_ _04361_ vssd1 vssd1 vccd1 vccd1 _04362_ sky130_fd_sc_hd__inv_2
XANTENNA__11838__B1 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08929__S1 net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout277_A net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08654_ top.CPU.alu.program_counter\[14\] net878 vssd1 vssd1 vccd1 vccd1 _04293_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_124_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11853__A3 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07605_ _03147_ net882 vssd1 vssd1 vccd1 vccd1 _03244_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_124_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10030__Y _05669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08585_ top.CPU.alu.program_counter\[15\] net878 vssd1 vssd1 vccd1 vccd1 _04224_
+ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout444_A net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11066__A1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07536_ net1402 net661 vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__and2_1
XFILLER_81_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08863__S net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08467__C1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11605__A3 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07467_ top.CPU.control_unit.instruction\[14\] vssd1 vssd1 vccd1 vccd1 _03107_ sky130_fd_sc_hd__inv_2
XANTENNA__10694__A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout232_X net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout611_A net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1353_A top.CPU.handler.state\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout709_A _03212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_22_Left_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14850__1020 clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 net2489 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_33_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09206_ top.CPU.registers.data\[582\] net1287 net1006 top.CPU.registers.data\[614\]
+ net930 vssd1 vssd1 vccd1 vccd1 _04845_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_33_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08164__A net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11302__B net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09137_ net683 _04774_ _04775_ net919 vssd1 vssd1 vccd1 vccd1 _04776_ sky130_fd_sc_hd__o211a_1
XFILLER_163_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08234__A2 net1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14374__544 clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 net2013 sky130_fd_sc_hd__inv_2
XFILLER_136_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09694__S net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09068_ _04705_ _04706_ net927 vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__mux2_1
XFILLER_162_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout980_A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12318__A1 _03915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout699_X net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09719__C1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08019_ top.CPU.registers.data\[436\] top.CPU.registers.data\[404\] net816 vssd1
+ vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__mux2_1
XFILLER_118_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold660 top.CPU.registers.data\[459\] vssd1 vssd1 vccd1 vccd1 net3217 sky130_fd_sc_hd__dlygate4sd3_1
Xhold671 top.CPU.registers.data\[790\] vssd1 vssd1 vccd1 vccd1 net3228 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1406_X net1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14415__585 clknet_leaf_177_clk vssd1 vssd1 vccd1 vccd1 net2054 sky130_fd_sc_hd__inv_2
X_11030_ net3938 net216 _06573_ net312 vssd1 vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_34_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold682 top.CPU.registers.data\[941\] vssd1 vssd1 vccd1 vccd1 net3239 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09195__B1 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold693 top.CPU.registers.data\[454\] vssd1 vssd1 vccd1 vccd1 net3250 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout866_X net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12981_ top.I2C.bit_timer_counter\[5\] _07411_ top.I2C.bit_timer_counter\[6\] vssd1
+ vssd1 vccd1 vccd1 _07413_ sky130_fd_sc_hd__a21o_1
XANTENNA__11829__B1 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09498__A1 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11464__S net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1360 top.I2C.data_out\[10\] vssd1 vssd1 vccd1 vccd1 net3917 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_40_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1371 top.I2C.data_out\[7\] vssd1 vssd1 vccd1 vccd1 net3928 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1382 top.mmio.mem_data_i\[24\] vssd1 vssd1 vccd1 vccd1 net3939 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11932_ net3678 net185 net342 _06465_ vssd1 vssd1 vccd1 vccd1 _01634_ sky130_fd_sc_hd__a22o_1
XANTENNA__10501__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1393 top.CPU.registers.data\[69\] vssd1 vssd1 vccd1 vccd1 net3950 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11844__A3 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11863_ _06699_ _06754_ net152 net3345 vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_150_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13602_ net3164 net579 _03027_ _03028_ vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__a22o_1
X_10814_ net549 _05127_ _05754_ _05889_ _06423_ vssd1 vssd1 vccd1 vccd1 _06424_ sky130_fd_sc_hd__o221a_1
XANTENNA__11057__A1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11794_ net429 net198 vssd1 vssd1 vccd1 vccd1 _06761_ sky130_fd_sc_hd__nand2_1
XANTENNA__08773__S net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07530__X _03169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16321_ clknet_leaf_66_clk _02530_ net1165 vssd1 vssd1 vccd1 vccd1 top.CPU.addressnew\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13533_ _05361_ net585 vssd1 vssd1 vccd1 vccd1 _02987_ sky130_fd_sc_hd__and2_1
X_10745_ _05273_ _05543_ vssd1 vssd1 vccd1 vccd1 _06358_ sky130_fd_sc_hd__nor2_1
X_13982__152 clknet_leaf_150_clk vssd1 vssd1 vccd1 vccd1 net1621 sky130_fd_sc_hd__inv_2
XFILLER_41_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xteam_08_1417 vssd1 vssd1 vccd1 vccd1 team_08_1417/HI gpio_oeb[3] sky130_fd_sc_hd__conb_1
Xteam_08_1428 vssd1 vssd1 vccd1 vccd1 team_08_1428/HI gpio_oeb[14] sky130_fd_sc_hd__conb_1
XFILLER_159_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16252_ clknet_leaf_61_clk _02462_ net1160 vssd1 vssd1 vccd1 vccd1 top.CPU.control_unit.instruction\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_13464_ top.CPU.handler.toreg\[21\] _02953_ net120 vssd1 vssd1 vccd1 vccd1 _02487_
+ sky130_fd_sc_hd__mux2_1
Xteam_08_1439 vssd1 vssd1 vccd1 vccd1 team_08_1439/HI gpio_out[24] sky130_fd_sc_hd__conb_1
X_10676_ net524 _06292_ vssd1 vssd1 vccd1 vccd1 _06293_ sky130_fd_sc_hd__nor2_1
XFILLER_159_83 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12415_ _06935_ _06937_ _06938_ _06940_ vssd1 vssd1 vccd1 vccd1 _06941_ sky130_fd_sc_hd__or4_4
X_15203_ net1537 _01413_ net1210 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13395_ top.mmio.mem_data_i\[24\] _07089_ net555 top.I2C.data_out\[24\] vssd1 vssd1
+ vccd1 vccd1 _02914_ sky130_fd_sc_hd__a22o_1
X_16183_ net2517 _02393_ net1182 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[983\]
+ sky130_fd_sc_hd__dfrtp_1
X_12346_ top.I2C.bit_timer_state\[1\] net1340 vssd1 vssd1 vccd1 vccd1 _06895_ sky130_fd_sc_hd__nand2_1
X_15134_ clknet_leaf_46_clk _01344_ net1137 vssd1 vssd1 vccd1 vccd1 top.I2C.data_out\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12309__A1 _03370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11780__A2 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15065_ clknet_leaf_52_clk _00044_ net1132 vssd1 vssd1 vccd1 vccd1 top.I2C.output_state\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_12277_ net3775 _03542_ net1235 vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__mux2_1
XFILLER_141_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11228_ _05933_ net545 net531 vssd1 vssd1 vccd1 vccd1 _06669_ sky130_fd_sc_hd__and3b_1
XANTENNA__08013__S net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11532__A2 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11159_ net521 _06448_ vssd1 vssd1 vccd1 vccd1 _06640_ sky130_fd_sc_hd__nor2_1
XANTENNA__13809__B2 top.CPU.data_out\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15967_ net2301 _02177_ net1219 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[767\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13285__A2 net1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10131__X _05769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12493__B1 _04952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08249__A _03887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15898_ net2232 _02108_ net1251 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[698\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11048__A1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08370_ top.CPU.registers.data\[466\] net1320 net851 top.CPU.registers.data\[498\]
+ net769 vssd1 vssd1 vccd1 vccd1 _04009_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_102_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11106__C net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09110__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16519_ clknet_leaf_92_clk _02681_ net1269 vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_82_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14061__231 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 net1700 sky130_fd_sc_hd__inv_2
XFILLER_149_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14358__528 clknet_leaf_181_clk vssd1 vssd1 vccd1 vccd1 net1997 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_30_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11122__B net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12933__S net1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14102__272 clknet_leaf_175_clk vssd1 vssd1 vccd1 vccd1 net1741 sky130_fd_sc_hd__inv_2
XFILLER_145_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09808__A net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12553__C_N top.CPU.done vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11771__A2 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_148_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15299__RESET_B net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09177__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout403 net404 vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09716__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout414 net415 vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__clkbuf_2
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout425 _06756_ vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout394_A net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11523__A2 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout436 _06467_ vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__buf_2
XANTENNA__08924__B1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout447 _05517_ vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__buf_2
X_09824_ net711 _05460_ _05461_ _05462_ vssd1 vssd1 vccd1 vccd1 _05463_ sky130_fd_sc_hd__a31o_1
Xfanout458 net463 vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_126_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout469 net470 vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12888__B _07322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09755_ _05392_ _05393_ net643 vssd1 vssd1 vccd1 vccd1 _05394_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout182_X net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout659_A net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08706_ _04335_ _04343_ _04344_ net702 vssd1 vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__a211o_1
X_09686_ top.CPU.registers.data\[345\] net1336 net869 top.CPU.registers.data\[377\]
+ net757 vssd1 vssd1 vccd1 vccd1 _05325_ sky130_fd_sc_hd__a221o_1
XFILLER_27_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08637_ top.CPU.registers.data\[46\] top.CPU.registers.data\[14\] net819 vssd1 vssd1
+ vccd1 vccd1 _04276_ sky130_fd_sc_hd__mux2_1
XFILLER_27_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15053__Q top.CPU.alu.program_counter\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout447_X net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout826_A net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14800__970 clknet_leaf_196_clk vssd1 vssd1 vccd1 vccd1 net2439 sky130_fd_sc_hd__inv_2
XANTENNA_fanout1189_X net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13966__136 clknet_leaf_166_clk vssd1 vssd1 vccd1 vccd1 net1605 sky130_fd_sc_hd__inv_2
X_08568_ net788 _04205_ _04206_ net641 vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__a31o_1
XANTENNA__12236__B1 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_30_Left_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07519_ net1409 net1408 top.CPU.control_unit.instruction\[6\] vssd1 vssd1 vccd1 vccd1
+ _03158_ sky130_fd_sc_hd__and3b_1
XFILLER_80_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13512__B _02966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08455__A2 _04090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout614_X net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08499_ net794 _04132_ _04133_ net745 vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__o211a_1
XFILLER_167_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12409__A _06918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10530_ _04397_ _04469_ _05284_ _05285_ vssd1 vssd1 vccd1 vccd1 _06153_ sky130_fd_sc_hd__o31a_1
XFILLER_128_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10461_ _05294_ _05297_ _06064_ vssd1 vssd1 vccd1 vccd1 _06087_ sky130_fd_sc_hd__a21bo_1
XANTENNA__08207__A2 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12200_ top.CPU.registers.data\[51\] net647 vssd1 vssd1 vccd1 vccd1 _06867_ sky130_fd_sc_hd__or2_1
X_13180_ top.I2C.I2C_state\[25\] top.I2C.I2C_state\[1\] top.I2C.within_byte_counter_writing\[0\]
+ top.I2C.within_byte_counter_writing\[1\] vssd1 vssd1 vccd1 vccd1 _02761_ sky130_fd_sc_hd__o211a_1
XFILLER_89_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10392_ _03755_ _03889_ net379 vssd1 vssd1 vccd1 vccd1 _06021_ sky130_fd_sc_hd__mux2_1
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout983_X net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07966__A1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12131_ net3966 net174 _06833_ _06736_ vssd1 vssd1 vccd1 vccd1 _01497_ sky130_fd_sc_hd__a22o_1
XANTENNA__11459__S net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07509__Y _03148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09168__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09707__A2 net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12062_ net568 net364 _06610_ net179 top.CPU.registers.data\[122\] vssd1 vssd1 vccd1
+ vccd1 _06800_ sky130_fd_sc_hd__a32o_1
Xhold490 net66 vssd1 vssd1 vccd1 vccd1 net3047 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07718__A1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11013_ net526 _06562_ vssd1 vssd1 vccd1 vccd1 _06563_ sky130_fd_sc_hd__nor2_1
XFILLER_150_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10722__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12798__B _04189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout970 net1003 vssd1 vssd1 vccd1 vccd1 net970 sky130_fd_sc_hd__buf_2
X_15821_ net2155 _02031_ net1071 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[621\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout981 net982 vssd1 vssd1 vccd1 vccd1 net981 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout992 net994 vssd1 vssd1 vccd1 vccd1 net992 sky130_fd_sc_hd__buf_4
XFILLER_46_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11278__B2 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15752_ net2086 _01962_ net1099 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[552\]
+ sky130_fd_sc_hd__dfrtp_1
X_12964_ net1411 _07401_ top.I2C.bit_timer_counter\[0\] vssd1 vssd1 vccd1 vccd1 _07402_
+ sky130_fd_sc_hd__mux2_1
X_14799__969 clknet_leaf_191_clk vssd1 vssd1 vccd1 vccd1 net2438 sky130_fd_sc_hd__inv_2
XFILLER_45_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08679__C1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08143__A1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1190 top.mmio.mem_data_i\[9\] vssd1 vssd1 vccd1 vccd1 net3747 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09340__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11915_ net3398 net185 net347 _06127_ vssd1 vssd1 vccd1 vccd1 _01651_ sky130_fd_sc_hd__a22o_1
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15683_ net2017 _01893_ net1206 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[483\]
+ sky130_fd_sc_hd__dfrtp_1
X_12895_ top.CPU.alu.program_counter\[25\] _05362_ vssd1 vssd1 vccd1 vccd1 _07340_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_47_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09599__S net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12227__B1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11846_ net464 _06677_ net239 net152 net2701 vssd1 vssd1 vccd1 vccd1 _01715_ sky130_fd_sc_hd__a32o_1
XFILLER_54_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14045__215 clknet_leaf_130_clk vssd1 vssd1 vccd1 vccd1 net1684 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_11_0_clk_X clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07701__A top.CPU.control_unit.instruction\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11777_ net462 _06620_ net236 net161 net2976 vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__a32o_1
X_16304_ clknet_leaf_107_clk _02513_ net1248 vssd1 vssd1 vccd1 vccd1 top.CPU.data_out\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13516_ top.CPU.data_out\[16\] net590 _02977_ net340 vssd1 vssd1 vccd1 vccd1 _02514_
+ sky130_fd_sc_hd__o22a_1
X_10728_ _05705_ _05715_ vssd1 vssd1 vccd1 vccd1 _06342_ sky130_fd_sc_hd__nor2_1
XANTENNA__08008__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08851__C1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11450__B2 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16235_ clknet_leaf_32_clk _02445_ net1125 vssd1 vssd1 vccd1 vccd1 top.CPU.control_unit.instruction\[11\]
+ sky130_fd_sc_hd__dfrtp_4
X_13447_ _02887_ _02937_ _02939_ vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__a21o_1
X_10659_ net548 _05279_ _06275_ vssd1 vssd1 vccd1 vccd1 _06276_ sky130_fd_sc_hd__o21ai_2
Xclkload13 clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clkload13/Y sky130_fd_sc_hd__clkinv_8
XFILLER_173_247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload24 clknet_leaf_200_clk vssd1 vssd1 vccd1 vccd1 clkload24/Y sky130_fd_sc_hd__inv_12
XANTENNA__11510__X _06733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload35 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 clkload35/Y sky130_fd_sc_hd__inv_6
Xclkload46 clknet_leaf_191_clk vssd1 vssd1 vccd1 vccd1 clkload46/Y sky130_fd_sc_hd__inv_16
XFILLER_173_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13378_ top.I2C.data_out\[19\] net556 _02901_ vssd1 vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__a21oi_1
XFILLER_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08603__C1 net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16166_ net2500 _02376_ net1072 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[966\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_142_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload57 clknet_leaf_177_clk vssd1 vssd1 vccd1 vccd1 clkload57/Y sky130_fd_sc_hd__clkinv_16
XFILLER_86_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload68 clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 clkload68/Y sky130_fd_sc_hd__clkinv_8
XFILLER_114_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload79 clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 clkload79/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__11753__A2 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15117_ net1499 _01330_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r2_prev\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_12329_ net2569 _04500_ net1236 vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__mux2_1
XFILLER_170_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16097_ net2431 _02307_ net1232 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[897\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_48_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15048_ clknet_leaf_93_clk _01293_ net1268 vssd1 vssd1 vccd1 vccd1 top.SPI.command\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_123_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12702__A1 top.CPU.alu.program_counter\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11505__A2 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07870_ _03508_ _03477_ net453 vssd1 vssd1 vccd1 vccd1 _03509_ sky130_fd_sc_hd__mux2_1
X_14743__913 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 net2382 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_143_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08382__A1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13911__81 clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 net1550 sky130_fd_sc_hd__inv_2
XFILLER_110_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12501__B _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07590__C1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09540_ top.CPU.registers.data\[33\] top.CPU.registers.data\[1\] net835 vssd1 vssd1
+ vccd1 vccd1 _05179_ sky130_fd_sc_hd__mux2_1
XANTENNA__12466__B1 _05330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09331__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09471_ top.CPU.registers.data\[962\] net1324 net855 top.CPU.registers.data\[994\]
+ net723 vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__a221o_1
XFILLER_36_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08685__A2 _04323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08422_ top.CPU.registers.data\[305\] top.CPU.registers.data\[273\] net825 vssd1
+ vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__mux2_1
XANTENNA__12218__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08353_ net694 _03991_ vssd1 vssd1 vccd1 vccd1 _03992_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_158_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout142_A _06253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08437__A2 net1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08284_ _03922_ vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__inv_2
Xclkload7 clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clkload7/Y sky130_fd_sc_hd__inv_6
XANTENNA__11992__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout407_A _05023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1051_A net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07757__S net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15409__RESET_B net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09493__S0 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11744__A2 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1316_A net1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout200 net201 vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__clkbuf_4
Xfanout1209 net1218 vssd1 vssd1 vccd1 vccd1 net1209 sky130_fd_sc_hd__buf_2
Xfanout211 _06753_ vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__buf_2
XANTENNA_fanout776_A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_892 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout222 net223 vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__clkbuf_8
XFILLER_8_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout233 net243 vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__clkbuf_4
Xfanout244 _06748_ vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10704__B1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout255 _06728_ vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__clkbuf_4
XFILLER_8_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14486__656 clknet_leaf_175_clk vssd1 vssd1 vccd1 vccd1 net2125 sky130_fd_sc_hd__inv_2
XANTENNA__09570__B1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout266 _06717_ vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__buf_4
XFILLER_75_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09807_ top.CPU.registers.data\[58\] top.CPU.registers.data\[26\] net838 vssd1 vssd1
+ vccd1 vccd1 _05446_ sky130_fd_sc_hd__mux2_1
Xfanout277 net278 vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__buf_4
XFILLER_75_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout288 _06712_ vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout564_X net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout299 _06645_ vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout943_A net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07999_ top.CPU.registers.data\[312\] net1010 net933 vssd1 vssd1 vccd1 vccd1 _03638_
+ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_105_Left_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09738_ top.CPU.registers.data\[59\] top.CPU.registers.data\[27\] net831 vssd1 vssd1
+ vccd1 vccd1 _05377_ sky130_fd_sc_hd__mux2_1
XFILLER_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10212__A net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12457__B1 _03541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09322__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14527__697 clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 net2166 sky130_fd_sc_hd__inv_2
XANTENNA_fanout731_X net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09669_ net757 _05306_ _05307_ _05305_ net642 vssd1 vssd1 vccd1 vccd1 _05308_ sky130_fd_sc_hd__a311o_1
XANTENNA_fanout829_X net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13523__A _03716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11700_ _06531_ net204 net422 net3306 vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__a22o_1
X_12680_ net125 _07141_ _03118_ vssd1 vssd1 vccd1 vccd1 _07146_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12209__B1 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11680__A1 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07884__B1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10866__B _05693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11631_ _05772_ net207 net427 net3176 vssd1 vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__a22o_1
XFILLER_24_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_145_Right_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11562_ _06539_ _06731_ vssd1 vssd1 vccd1 vccd1 _06742_ sky130_fd_sc_hd__nor2_1
XANTENNA__08833__C1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11432__B2 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10513_ net397 _06135_ _06136_ vssd1 vssd1 vccd1 vccd1 _06137_ sky130_fd_sc_hd__o21ai_1
X_13301_ top.mmio.mem_data_i\[0\] net592 net1344 vssd1 vssd1 vccd1 vccd1 _02844_ sky130_fd_sc_hd__a21o_1
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11983__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10640__C1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11493_ net482 net471 _06623_ net254 net2916 vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__a32o_1
XANTENNA__10882__A _05693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13232_ net2873 _02776_ _02799_ vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__mux2_1
XANTENNA__09389__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16020_ net2354 _02230_ net1120 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[820\]
+ sky130_fd_sc_hd__dfrtp_1
X_10444_ _05976_ _06070_ net389 vssd1 vssd1 vccd1 vccd1 _06071_ sky130_fd_sc_hd__mux2_1
XFILLER_171_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11735__A2 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13163_ net3936 top.I2C.output_state\[10\] top.I2C.output_state\[16\] _02750_ vssd1
+ vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__or4b_1
XANTENNA__10093__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08061__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10375_ _05759_ _06001_ _06000_ vssd1 vssd1 vccd1 vccd1 _06005_ sky130_fd_sc_hd__a21oi_1
XFILLER_124_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14430__600 clknet_leaf_152_clk vssd1 vssd1 vccd1 vccd1 net2069 sky130_fd_sc_hd__inv_2
XFILLER_124_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12114_ net354 net233 vssd1 vssd1 vccd1 vccd1 _06825_ sky130_fd_sc_hd__nand2_4
X_13094_ top.CPU.data_out\[29\] net2757 net558 vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__mux2_1
XFILLER_3_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12045_ _06594_ _06779_ net150 net3310 vssd1 vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_88_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08364__A1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12160__A2 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09561__B1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10171__A1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15804_ net2138 _02014_ net1195 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[604\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11218__A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15735_ net2069 _01945_ net1180 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[535\]
+ sky130_fd_sc_hd__dfrtp_1
X_12947_ _07384_ _07385_ vssd1 vssd1 vccd1 vccd1 _07387_ sky130_fd_sc_hd__xor2_1
XANTENNA__08667__A2 net1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11671__A1 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15666_ net2000 _01876_ net1103 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[466\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07875__B1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12878_ _07324_ _07321_ net126 vssd1 vssd1 vccd1 vccd1 _07325_ sky130_fd_sc_hd__mux2_1
XFILLER_60_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11829_ _06520_ _06648_ net241 net158 net2862 vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__a32o_1
X_15597_ net1931 _01807_ net1064 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[397\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_112_Right_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10631__C1 _06249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11974__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload102 clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 clkload102/Y sky130_fd_sc_hd__bufinv_16
Xclkload113 clknet_leaf_159_clk vssd1 vssd1 vccd1 vccd1 clkload113/Y sky130_fd_sc_hd__inv_6
X_16218_ net2552 _02428_ net1243 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[1018\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload124 clknet_leaf_165_clk vssd1 vssd1 vccd1 vccd1 clkload124/Y sky130_fd_sc_hd__inv_6
Xclkload135 clknet_leaf_143_clk vssd1 vssd1 vccd1 vccd1 clkload135/Y sky130_fd_sc_hd__clkinv_8
XFILLER_143_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08262__A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload146 clknet_leaf_122_clk vssd1 vssd1 vccd1 vccd1 clkload146/Y sky130_fd_sc_hd__inv_8
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11187__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload157 clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 clkload157/Y sky130_fd_sc_hd__inv_2
Xclkload168 clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 clkload168/Y sky130_fd_sc_hd__inv_6
XANTENNA__11726__A2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_111 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16149_ net2483 _02359_ net1217 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[949\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload179 clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 clkload179/Y sky130_fd_sc_hd__inv_6
XANTENNA__08052__B1 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14173__343 clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 net1812 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_77_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08971_ net640 _04606_ _04609_ vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__or3_1
XANTENNA__09227__S0 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13479__A2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13888__58 clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 net1527 sky130_fd_sc_hd__inv_2
XANTENNA__11827__S net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07922_ top.CPU.registers.data\[988\] net1302 net1023 top.CPU.registers.data\[1020\]
+ net919 vssd1 vssd1 vccd1 vccd1 _03561_ sky130_fd_sc_hd__a221o_1
Xhold19 top.CPU.registers.data_out_r2_prev\[27\] vssd1 vssd1 vccd1 vccd1 net2576 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_60_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12151__A2 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14214__384 clknet_leaf_125_clk vssd1 vssd1 vccd1 vccd1 net1853 sky130_fd_sc_hd__inv_2
XFILLER_96_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07853_ top.CPU.registers.data_out_r2_prev\[29\] net685 net618 _03485_ _03491_ vssd1
+ vssd1 vccd1 vccd1 _03492_ sky130_fd_sc_hd__o2111a_1
XFILLER_111_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11128__A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07784_ top.CPU.registers.data\[926\] net1303 net1025 top.CPU.registers.data\[958\]
+ net621 vssd1 vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__a221o_1
XFILLER_37_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09523_ top.CPU.registers.data\[897\] net1335 net868 top.CPU.registers.data\[929\]
+ net733 vssd1 vssd1 vccd1 vccd1 _05162_ sky130_fd_sc_hd__a221o_1
XANTENNA__11111__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10967__A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout357_A net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09454_ top.CPU.registers.data\[34\] top.CPU.registers.data\[2\] net823 vssd1 vssd1
+ vccd1 vccd1 _05093_ sky130_fd_sc_hd__mux2_1
XFILLER_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07866__B1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09032__S net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08405_ top.CPU.registers.data\[338\] net1291 net1012 top.CPU.registers.data\[370\]
+ net934 vssd1 vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__a221o_1
X_09385_ _05019_ _05022_ net454 vssd1 vssd1 vccd1 vccd1 _05024_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout145_X net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout524_A net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1266_A net1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08336_ _03973_ _03974_ net938 vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__mux2_1
XANTENNA__08724__X _04363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08815__C1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09083__A2 net1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11965__A2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08267_ top.CPU.registers.data\[758\] net1382 net998 top.CPU.registers.data\[726\]
+ net923 vssd1 vssd1 vccd1 vccd1 _03906_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_140_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_140_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout312_X net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1054_X net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09268__A net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08198_ net679 _03832_ _03833_ _03836_ net612 vssd1 vssd1 vccd1 vccd1 _03837_ sky130_fd_sc_hd__a311o_1
XANTENNA__11717__A2 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09240__C1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1319_X net1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09791__A0 _05428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11193__A3 _06648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10160_ net414 _05667_ _05787_ net510 _03511_ vssd1 vssd1 vccd1 vccd1 _05797_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_7_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout681_X net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout779_X net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1006 net1013 vssd1 vssd1 vccd1 vccd1 net1006 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16449__RESET_B net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10091_ _03958_ net373 vssd1 vssd1 vccd1 vccd1 _05729_ sky130_fd_sc_hd__nor2_1
Xfanout1017 net1022 vssd1 vssd1 vccd1 vccd1 net1017 sky130_fd_sc_hd__buf_2
XFILLER_126_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1028 net1029 vssd1 vssd1 vccd1 vccd1 net1028 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1039 _03177_ vssd1 vssd1 vccd1 vccd1 net1039 sky130_fd_sc_hd__buf_2
XANTENNA__12142__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09543__B1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout946_X net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11350__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12801_ _07232_ _07245_ vssd1 vssd1 vccd1 vccd1 _07255_ sky130_fd_sc_hd__nand2_1
XFILLER_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13781_ net9 net1049 net884 net3260 vssd1 vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__o22a_1
X_10993_ net2821 net216 _06550_ net314 vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_172_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10877__A net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11472__S net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15520_ net1854 _01730_ net1094 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[320\]
+ sky130_fd_sc_hd__dfrtp_1
X_12732_ top.CPU.alu.program_counter\[9\] _07173_ top.CPU.alu.program_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _07192_ sky130_fd_sc_hd__a21oi_1
XFILLER_37_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_52_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15451_ net1785 _01661_ net1213 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[251\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ top.CPU.alu.program_counter\[3\] _05021_ vssd1 vssd1 vccd1 vccd1 _07130_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_61_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11614_ _06212_ net3301 net212 vssd1 vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_187_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15382_ net1716 _01592_ net1228 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[182\]
+ sky130_fd_sc_hd__dfrtp_1
X_12594_ top.SPI.command\[1\] top.SPI.command\[5\] _07093_ _07094_ vssd1 vssd1 vccd1
+ vccd1 _07095_ sky130_fd_sc_hd__and4bb_1
XANTENNA__09074__A2 net1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11956__A2 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11545_ _06661_ net260 net252 net3232 vssd1 vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_67_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_131_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_131_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_98_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11476_ net563 net526 _05810_ vssd1 vssd1 vccd1 vccd1 _06729_ sky130_fd_sc_hd__and3_1
XANTENNA__08082__A _03683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_110_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14157__327 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 net1796 sky130_fd_sc_hd__inv_2
XFILLER_171_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16003_ net2337 _02213_ net1208 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[803\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11708__A2 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13215_ top.I2C.within_byte_counter_reading\[2\] _02753_ vssd1 vssd1 vccd1 vccd1
+ _02789_ sky130_fd_sc_hd__or2_2
X_10427_ net600 _06054_ vssd1 vssd1 vccd1 vccd1 _06055_ sky130_fd_sc_hd__nor2_1
XANTENNA__11220__B net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09231__C1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10916__B1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09782__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13146_ top.CPU.alu.program_counter\[0\] top.CPU.alu.program_counter\[1\] top.CPU.alu.program_counter\[31\]
+ _07390_ vssd1 vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__and4_1
X_10358_ top.CPU.fetch.current_ra\[23\] net1041 net633 top.CPU.handler.toreg\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05989_ sky130_fd_sc_hd__a22oi_4
XANTENNA__10392__A1 _03889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13077_ top.CPU.data_out\[12\] net3349 net559 vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__mux2_1
XANTENNA__09625__B net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10289_ _05786_ _05912_ net390 vssd1 vssd1 vccd1 vccd1 _05922_ sky130_fd_sc_hd__mux2_1
XANTENNA__10404__X _06033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_125_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08337__A1 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12133__A2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12028_ top.CPU.registers.data\[147\] net651 vssd1 vssd1 vccd1 vccd1 _06791_ sky130_fd_sc_hd__or2_1
XFILLER_111_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_198_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_198_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_38_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11341__B1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13094__A0 top.CPU.data_out\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09298__C1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15718_ net2052 _01928_ net1081 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[518\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10852__C1 _06141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16247__Q top.CPU.control_unit.instruction\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15649_ net1983 _01859_ net1224 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[449\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_22_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09170_ top.CPU.registers.data\[294\] top.CPU.registers.data\[262\] net814 vssd1
+ vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_155_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08121_ net941 _03757_ _03759_ net620 vssd1 vssd1 vccd1 vccd1 _03760_ sky130_fd_sc_hd__o211a_1
XANTENNA__11947__A2 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13610__B _05958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08273__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09470__C1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_122_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_122_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10080__A0 _04294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10953__C net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08052_ top.CPU.registers.data\[244\] net1379 net979 top.CPU.registers.data\[212\]
+ net905 vssd1 vssd1 vccd1 vccd1 _03691_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_12_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11130__B net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10027__A net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10907__B1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09773__B1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07784__C1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11580__B1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08954_ net611 _04572_ _04579_ _04592_ vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__a31o_2
XFILLER_88_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1014_A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09525__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12124__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07905_ net1036 _03541_ _03543_ vssd1 vssd1 vccd1 vccd1 _03544_ sky130_fd_sc_hd__a21oi_4
X_08885_ net786 _04523_ vssd1 vssd1 vccd1 vccd1 _04524_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_189_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_189_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08879__A2 net1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout474_A _03193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11332__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07836_ _03474_ vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__inv_2
XANTENNA__08866__S net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07623__X _03262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09828__A1 _05465_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07767_ _03405_ vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__inv_2
XANTENNA__09289__C1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10697__A net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout262_X net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout641_A net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1383_A net1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout739_A net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09506_ net622 _05143_ _05144_ vssd1 vssd1 vccd1 vccd1 _05145_ sky130_fd_sc_hd__and3_1
XANTENNA__07839__B1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07698_ net1409 _03154_ net1278 net1285 _03104_ vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__a2111o_1
X_14598__768 clknet_leaf_122_clk vssd1 vssd1 vccd1 vccd1 net2237 sky130_fd_sc_hd__inv_2
XFILLER_40_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09437_ net954 _05075_ _05074_ net606 vssd1 vssd1 vccd1 vccd1 _05076_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_23_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout527_X net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout906_A net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09368_ net679 _05005_ _05006_ vssd1 vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__and3_1
XANTENNA__11399__B1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11938__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08319_ net880 _03955_ _03957_ vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__o21ai_2
XFILLER_166_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09299_ top.CPU.registers.data\[580\] net1299 net1020 top.CPU.registers.data\[612\]
+ net940 vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_113_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_113_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09461__C1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11330_ net490 net474 _05695_ net287 net2717 vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__a32o_1
XANTENNA__10610__A2 _06228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout896_X net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11261_ net513 _06555_ vssd1 vssd1 vccd1 vccd1 _06687_ sky130_fd_sc_hd__nor2_1
XANTENNA__12851__S net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09213__C1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13000_ net1354 net1410 vssd1 vssd1 vccd1 vccd1 _07428_ sky130_fd_sc_hd__nand2_2
XANTENNA__12363__A2 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07945__S net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10212_ net661 _05847_ vssd1 vssd1 vccd1 vccd1 _05848_ sky130_fd_sc_hd__and2_1
XANTENNA__09726__A _05332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11192_ net143 net3597 net297 vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__mux2_1
XANTENNA__10374__A1 _05687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11571__B1 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10143_ _05633_ _05638_ net306 vssd1 vssd1 vccd1 vccd1 _05780_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08319__A1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09516__B1 net1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07790__A2 net1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input35_A gpio_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14951_ clknet_leaf_52_clk _01197_ net1133 vssd1 vssd1 vccd1 vccd1 top.I2C.bit_timer_counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10074_ _05711_ vssd1 vssd1 vccd1 vccd1 _05712_ sky130_fd_sc_hd__inv_2
XANTENNA__10126__A1 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11323__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10677__A2 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14542__712 clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 net2181 sky130_fd_sc_hd__inv_2
X_16621_ top.I2C.sda_oeb vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__clkbuf_1
XANTENNA__13076__A0 top.CPU.data_out\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16552_ clknet_leaf_64_clk net4000 net1162 vssd1 vssd1 vccd1 vccd1 top.mmio.s1 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11626__A1 _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13764_ net1346 net1052 top.wm.prev_BUSY_O vssd1 vssd1 vccd1 vccd1 _03095_ sky130_fd_sc_hd__or3b_2
XANTENNA__09295__A2 net1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10976_ net526 _06539_ vssd1 vssd1 vccd1 vccd1 _06540_ sky130_fd_sc_hd__nor2_1
X_15503_ net1837 _01713_ net1095 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[303\]
+ sky130_fd_sc_hd__dfrtp_1
X_12715_ top.CPU.alu.program_counter\[8\] _04728_ vssd1 vssd1 vccd1 vccd1 _07177_
+ sky130_fd_sc_hd__or2_1
XANTENNA__11215__B net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16483_ clknet_leaf_58_clk _02645_ net1143 vssd1 vssd1 vccd1 vccd1 top.I2C.which_data_address\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13695_ top.SPI.timem\[1\] _03049_ vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__and2_1
X_15434_ net1768 _01644_ net1085 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[234\]
+ sky130_fd_sc_hd__dfrtp_1
X_12646_ top.I2C.output_state\[20\] top.I2C.initiate_read_bit _06948_ vssd1 vssd1
+ vccd1 vccd1 _00019_ sky130_fd_sc_hd__and3_1
XFILLER_62_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11929__A2 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15365_ net1699 _01575_ net1062 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[165\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_104_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_104_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12577_ _07054_ _03101_ _03246_ vssd1 vssd1 vccd1 vccd1 _07082_ sky130_fd_sc_hd__or3b_1
XFILLER_12_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11528_ _06653_ net260 net252 net3347 vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__a22o_1
X_15296_ net1630 _01506_ net1096 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[96\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_116_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold308 top.CPU.registers.data\[21\] vssd1 vssd1 vccd1 vccd1 net2865 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08007__B1 _03408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold319 top.CPU.registers.data\[428\] vssd1 vssd1 vccd1 vccd1 net2876 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09204__C1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11459_ _06212_ net3163 net264 vssd1 vssd1 vccd1 vccd1 _02063_ sky130_fd_sc_hd__mux2_1
XANTENNA__13551__A1 _06445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09755__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13129_ top.SPI.command\[3\] top.SPI.command\[5\] _07093_ _02731_ vssd1 vssd1 vccd1
+ vccd1 _02732_ sky130_fd_sc_hd__and4_1
XFILLER_98_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13858__28 clknet_leaf_140_clk vssd1 vssd1 vccd1 vccd1 net1497 sky130_fd_sc_hd__inv_2
XANTENNA__12106__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09507__B1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07781__A2 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1008 top.CPU.registers.data\[918\] vssd1 vssd1 vccd1 vccd1 net3565 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1019 top.CPU.registers.data\[945\] vssd1 vssd1 vccd1 vccd1 net3576 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11314__B1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1370 net1377 vssd1 vssd1 vccd1 vccd1 net1370 sky130_fd_sc_hd__clkbuf_2
XFILLER_94_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08670_ net619 _04301_ _04307_ _04308_ vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__o22a_1
Xfanout1381 net1383 vssd1 vssd1 vccd1 vccd1 net1381 sky130_fd_sc_hd__clkbuf_4
Xfanout1392 net1393 vssd1 vssd1 vccd1 vccd1 net1392 sky130_fd_sc_hd__clkbuf_4
X_07621_ net1397 _03259_ vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__nor2_1
XANTENNA__13067__A0 top.CPU.data_out\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14285__455 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 net1924 sky130_fd_sc_hd__inv_2
XFILLER_26_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07552_ _03173_ net323 vssd1 vssd1 vccd1 vccd1 _03191_ sky130_fd_sc_hd__nand2_1
X_07483_ top.I2C.output_state\[20\] vssd1 vssd1 vccd1 vccd1 _03123_ sky130_fd_sc_hd__inv_2
XANTENNA__08494__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14326__496 clknet_leaf_179_clk vssd1 vssd1 vccd1 vccd1 net1965 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09222_ _04860_ vssd1 vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__inv_2
XFILLER_50_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_170_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09153_ net628 _04790_ _04791_ _04778_ vssd1 vssd1 vccd1 vccd1 _04792_ sky130_fd_sc_hd__a31o_4
XFILLER_159_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09443__C1 net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout222_A net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09994__A0 _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11141__A net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08104_ top.CPU.registers.data\[309\] top.CPU.registers.data\[277\] net830 vssd1
+ vssd1 vccd1 vccd1 _03743_ sky130_fd_sc_hd__mux2_1
XANTENNA__10053__B1 _05691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09084_ net1284 _04721_ _04722_ vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__or3_1
XFILLER_107_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10028__Y _05667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08035_ top.CPU.registers.data\[660\] net1319 net850 top.CPU.registers.data\[692\]
+ net719 vssd1 vssd1 vccd1 vccd1 _03674_ sky130_fd_sc_hd__a221o_1
XFILLER_135_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold820 top.CPU.registers.data\[328\] vssd1 vssd1 vccd1 vccd1 net3377 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_174_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1131_A net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold831 top.CPU.registers.data\[1002\] vssd1 vssd1 vccd1 vccd1 net3388 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08549__A1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13542__A1 top.CPU.data_out\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1229_A net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold842 top.CPU.registers.data\[536\] vssd1 vssd1 vccd1 vccd1 net3399 sky130_fd_sc_hd__dlygate4sd3_1
Xhold853 top.CPU.registers.data\[716\] vssd1 vssd1 vccd1 vccd1 net3410 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold864 top.CPU.registers.data\[372\] vssd1 vssd1 vccd1 vccd1 net3421 sky130_fd_sc_hd__dlygate4sd3_1
Xhold875 top.CPU.registers.data\[642\] vssd1 vssd1 vccd1 vccd1 net3432 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09210__A2 net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11553__B1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap594 net595 vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__clkbuf_1
XANTENNA_fanout689_A _03331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold886 top.CPU.registers.data\[757\] vssd1 vssd1 vccd1 vccd1 net3443 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_168_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold897 top.CPU.registers.data\[617\] vssd1 vssd1 vccd1 vccd1 net3454 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_107_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09986_ _04765_ net377 vssd1 vssd1 vccd1 vccd1 _05625_ sky130_fd_sc_hd__nor2_1
XFILLER_67_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1017_X net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10108__A1 _03613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08937_ top.CPU.registers.data\[74\] net1374 net972 top.CPU.registers.data\[106\]
+ net902 vssd1 vssd1 vccd1 vccd1 _04576_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_129_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout856_A net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout477_X net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11305__B1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08868_ net783 _04505_ _04506_ net737 vssd1 vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__o211a_1
XANTENNA__08596__S net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08721__A1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07819_ net1308 _03455_ _03456_ _03457_ vssd1 vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__o22a_1
X_13872__42 clknet_leaf_198_clk vssd1 vssd1 vccd1 vccd1 net1511 sky130_fd_sc_hd__inv_2
XANTENNA_fanout644_X net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08799_ top.CPU.registers.data\[44\] top.CPU.registers.data\[12\] net978 vssd1 vssd1
+ vccd1 vccd1 _04438_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1386_X net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10830_ _06438_ _06433_ _06436_ vssd1 vssd1 vccd1 vccd1 _06439_ sky130_fd_sc_hd__or3b_1
XFILLER_72_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08485__A0 _04122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11084__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10761_ net438 _06373_ vssd1 vssd1 vccd1 vccd1 _06374_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout811_X net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout909_X net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13531__A _03645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12500_ _07002_ _07003_ _07007_ _07008_ vssd1 vssd1 vccd1 vccd1 _07009_ sky130_fd_sc_hd__a22o_1
XFILLER_160_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13480_ net2744 _02961_ net123 vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__mux2_1
X_10692_ _04732_ _05564_ vssd1 vssd1 vccd1 vccd1 _06308_ sky130_fd_sc_hd__xor2_1
XANTENNA__08184__X _03823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12431_ net1341 top.I2C.output_state\[11\] net2741 vssd1 vssd1 vccd1 vccd1 _06952_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_157_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08237__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09434__C1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11051__A _06033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10593__C _06213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15150_ clknet_leaf_48_clk _01360_ net1128 vssd1 vssd1 vccd1 vccd1 top.I2C.data_out\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12362_ _03119_ _06904_ vssd1 vssd1 vccd1 vccd1 _06905_ sky130_fd_sc_hd__nor2_1
XFILLER_4_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11792__B1 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07996__C1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11313_ net2981 net289 net357 _06212_ vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__a22o_1
X_15081_ clknet_leaf_51_clk _00058_ net1132 vssd1 vssd1 vccd1 vccd1 top.I2C.output_state\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10890__A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12293_ net3766 _04292_ net1108 vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07528__X _03167_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09737__B1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11244_ net528 net442 net140 net545 vssd1 vssd1 vccd1 vccd1 _06677_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_91_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11544__B1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07748__C1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_51 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11175_ _05693_ _06479_ _06648_ vssd1 vssd1 vccd1 vccd1 _06649_ sky130_fd_sc_hd__and3_1
XANTENNA__10898__A2 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10126_ net404 _05643_ _05732_ _05756_ _05763_ vssd1 vssd1 vccd1 vccd1 _05764_ sky130_fd_sc_hd__o311a_1
XANTENNA__08960__A1 _04598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15983_ net2317 _02193_ net1095 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[783\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10114__B _05616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14269__439 clknet_leaf_133_clk vssd1 vssd1 vccd1 vccd1 net1908 sky130_fd_sc_hd__inv_2
X_14934_ clknet_leaf_70_clk _01180_ net1169 vssd1 vssd1 vccd1 vccd1 top.CPU.alu.program_counter\[17\]
+ sky130_fd_sc_hd__dfrtp_2
X_10057_ net3578 net227 net320 _05695_ vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__a22o_1
XANTENNA__11847__A1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08173__C1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07704__A top.CPU.control_unit.instruction\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14013__183 clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 net1652 sky130_fd_sc_hd__inv_2
XANTENNA_clkload0_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11226__A net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13816_ net2971 net335 net328 top.CPU.data_out\[18\] vssd1 vssd1 vccd1 vccd1 _02696_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10130__A net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16535_ clknet_leaf_99_clk _02697_ net1270 vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10807__C1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13747_ top.SPI.timem\[20\] _03082_ net3862 vssd1 vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__a21oi_1
X_10959_ net3402 net217 _06530_ net321 vssd1 vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_14_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16466_ clknet_leaf_86_clk _02628_ net1264 vssd1 vssd1 vccd1 vccd1 top.SPI.timem\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13678_ net2639 net336 vssd1 vssd1 vccd1 vccd1 _02606_ sky130_fd_sc_hd__and2_1
XANTENNA__08535__A net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15417_ net1751 _01627_ net1238 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[217\]
+ sky130_fd_sc_hd__dfrtp_1
X_12629_ net1340 top.I2C.output_state\[18\] top.I2C.output_state\[11\] vssd1 vssd1
+ vccd1 vccd1 _07120_ sky130_fd_sc_hd__a21o_1
XANTENNA__08228__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16397_ clknet_leaf_65_clk _00021_ net1162 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.next_counter_on
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10129__X _05767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14670__840 clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 net2309 sky130_fd_sc_hd__inv_2
X_15348_ net1682 _01558_ net1082 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[148\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10586__A1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11783__B1 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07987__C1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold105 top.CPU.registers.data\[572\] vssd1 vssd1 vccd1 vccd1 net2662 sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 net53 vssd1 vssd1 vccd1 vccd1 net2673 sky130_fd_sc_hd__dlygate4sd3_1
X_15279_ net1613 _01489_ net1105 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[79\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_171_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold127 _01209_ vssd1 vssd1 vccd1 vccd1 net2684 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 top.SPI.paroutput\[10\] vssd1 vssd1 vccd1 vccd1 net2695 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 net52 vssd1 vssd1 vccd1 vccd1 net2706 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14711__881 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 net2350 sky130_fd_sc_hd__inv_2
XFILLER_160_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11535__B1 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout607 net609 vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__clkbuf_4
X_09840_ top.CPU.registers.data\[666\] net1305 net1027 top.CPU.registers.data\[698\]
+ net921 vssd1 vssd1 vccd1 vccd1 _05479_ sky130_fd_sc_hd__a221o_1
XANTENNA__08400__B1 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout618 net619 vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__buf_4
Xfanout629 net630 vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__buf_2
XFILLER_101_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07754__A2 net1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09771_ top.CPU.registers.data\[187\] net1381 net990 top.CPU.registers.data\[155\]
+ net680 vssd1 vssd1 vccd1 vccd1 _05410_ sky130_fd_sc_hd__a221o_1
XANTENNA__10024__B net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08722_ top.CPU.registers.data_out_r1_prev\[13\] net871 net635 _04360_ _04346_ vssd1
+ vssd1 vccd1 vccd1 _04361_ sky130_fd_sc_hd__o221a_4
XTAP_TAPCELL_ROW_163_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08653_ _04291_ vssd1 vssd1 vccd1 vccd1 _04292_ sky130_fd_sc_hd__inv_2
XANTENNA__10510__A1 _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout172_A _06825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07911__C1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07604_ net417 vssd1 vssd1 vccd1 vccd1 _03243_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_124_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11136__A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09259__A2 net1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08584_ _04222_ vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_141_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13460__A0 top.CPU.handler.toreg\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12263__A1 _06311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08467__B1 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07535_ net1403 net572 vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__nand2_1
XANTENNA__11066__A2 _06230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10975__A net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout437_A _06467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1179_A net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10813__A2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07466_ top.CPU.alu.program_counter\[0\] vssd1 vssd1 vccd1 vccd1 _03106_ sky130_fd_sc_hd__inv_2
XANTENNA__10694__B _06309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09205_ top.CPU.registers.data\[966\] net1287 net1006 top.CPU.registers.data\[998\]
+ net904 vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_33_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout225_X net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout604_A net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1346_A net1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09136_ top.CPU.registers.data\[71\] net1304 net1024 top.CPU.registers.data\[103\]
+ net958 vssd1 vssd1 vccd1 vccd1 _04775_ sky130_fd_sc_hd__a221o_1
XFILLER_163_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11302__C _05694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11774__B1 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09067_ top.CPU.registers.data\[168\] top.CPU.registers.data\[136\] net969 vssd1
+ vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__mux2_1
XFILLER_118_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08451__Y _04090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13515__A1 _03369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08018_ top.CPU.registers.data\[244\] net1389 net816 top.CPU.registers.data\[212\]
+ net768 vssd1 vssd1 vccd1 vccd1 _03657_ sky130_fd_sc_hd__a221o_1
XFILLER_150_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold650 top.CPU.registers.data\[774\] vssd1 vssd1 vccd1 vccd1 net3207 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11526__B1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout973_A net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold661 top.CPU.registers.data\[915\] vssd1 vssd1 vccd1 vccd1 net3218 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold672 top.CPU.registers.data\[189\] vssd1 vssd1 vccd1 vccd1 net3229 sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 top.CPU.registers.data\[209\] vssd1 vssd1 vccd1 vccd1 net3240 sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 top.CPU.registers.data\[137\] vssd1 vssd1 vccd1 vccd1 net3251 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_34_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1301_X net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07745__A2 net1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09969_ _05527_ _05606_ vssd1 vssd1 vccd1 vccd1 _05608_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout859_X net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12980_ net2734 _07411_ _07412_ vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__a21oi_1
XFILLER_134_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1350 top.CPU.registers.data\[149\] vssd1 vssd1 vccd1 vccd1 net3907 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1361 top.mmio.mem_data_i\[10\] vssd1 vssd1 vccd1 vccd1 net3918 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1372 top.mmio.mem_data_i\[2\] vssd1 vssd1 vccd1 vccd1 net3929 sky130_fd_sc_hd__dlygate4sd3_1
X_11931_ net3561 net186 net351 _06449_ vssd1 vssd1 vccd1 vccd1 _01635_ sky130_fd_sc_hd__a22o_1
Xhold1383 top.CPU.registers.data\[81\] vssd1 vssd1 vccd1 vccd1 net3940 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1394 top.CPU.handler.state\[5\] vssd1 vssd1 vccd1 vccd1 net3951 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10501__B2 top.CPU.handler.toreg\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11046__A _05960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11862_ _06698_ net208 net155 net2692 vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__a22o_1
XFILLER_26_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13601_ top.CPU.alu.program_counter\[20\] net1348 net583 vssd1 vssd1 vccd1 vccd1
+ _03028_ sky130_fd_sc_hd__o21a_1
X_10813_ _05126_ net508 net504 _05124_ net443 vssd1 vssd1 vccd1 vccd1 _06423_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_0_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12254__A1 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11057__A2 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11793_ _06641_ net198 net160 net2975 vssd1 vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_49_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16320_ clknet_leaf_108_clk _02529_ net1249 vssd1 vssd1 vccd1 vccd1 top.CPU.data_out\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_13532_ net3984 net590 net340 _02986_ vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__o22a_1
X_10744_ net3881 net225 net313 _06357_ vssd1 vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__a22o_1
XFILLER_158_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09670__A2 net1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14654__824 clknet_leaf_152_clk vssd1 vssd1 vccd1 vccd1 net2293 sky130_fd_sc_hd__inv_2
X_16251_ clknet_leaf_60_clk _02461_ net1160 vssd1 vssd1 vccd1 vccd1 top.CPU.control_unit.instruction\[27\]
+ sky130_fd_sc_hd__dfrtp_2
Xteam_08_1418 vssd1 vssd1 vccd1 vccd1 team_08_1418/HI gpio_oeb[4] sky130_fd_sc_hd__conb_1
XFILLER_158_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13463_ net1396 net873 _02908_ net418 vssd1 vssd1 vccd1 vccd1 _02953_ sky130_fd_sc_hd__a31o_1
Xteam_08_1429 vssd1 vssd1 vccd1 vccd1 team_08_1429/HI gpio_out[0] sky130_fd_sc_hd__conb_1
XFILLER_13_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10675_ net551 _06291_ vssd1 vssd1 vccd1 vccd1 _06292_ sky130_fd_sc_hd__or2_1
XFILLER_159_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15202_ net1536 _01412_ net1175 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_12414_ _06920_ _06928_ _06939_ vssd1 vssd1 vccd1 vccd1 _06940_ sky130_fd_sc_hd__or3_1
XANTENNA__09958__B1 _05367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16182_ net2516 _02392_ net1227 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[982\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10568__A1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13394_ top.CPU.control_unit.instruction\[23\] _02913_ net667 vssd1 vssd1 vccd1 vccd1
+ _02457_ sky130_fd_sc_hd__mux2_1
XANTENNA__11765__B1 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15133_ clknet_leaf_48_clk _01343_ net1130 vssd1 vssd1 vccd1 vccd1 top.I2C.data_out\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_12345_ net1411 net1341 vssd1 vssd1 vccd1 vccd1 _06894_ sky130_fd_sc_hd__and2_1
XFILLER_4_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09186__A net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07984__A2 net1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15064_ clknet_leaf_50_clk _00043_ net1129 vssd1 vssd1 vccd1 vccd1 top.I2C.output_state\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_142_838 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12276_ net2635 _03474_ net1120 vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__mux2_1
XANTENNA__11517__B1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11227_ net495 net469 _06668_ net296 net2814 vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__a32o_1
XFILLER_122_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12190__B1 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08933__A1 net1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11158_ net3742 net303 _06639_ net488 vssd1 vssd1 vccd1 vccd1 _02276_ sky130_fd_sc_hd__a22o_1
XANTENNA__10740__A1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10109_ _05744_ _05746_ net384 vssd1 vssd1 vccd1 vccd1 _05747_ sky130_fd_sc_hd__mux2_1
X_11089_ _03186_ net501 vssd1 vssd1 vccd1 vccd1 _06600_ sky130_fd_sc_hd__nor2_1
X_15966_ net2300 _02176_ net1203 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[766\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15527__RESET_B net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12493__B2 _04986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15897_ net2231 _02107_ net1245 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[697\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_159_Right_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12994__B net1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08449__B1 net1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16518_ clknet_leaf_98_clk _02680_ net1257 vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07657__D1 net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16255__Q top.CPU.alu.immediate\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16449_ clknet_leaf_81_clk _02612_ net1242 vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__dfrtp_1
XFILLER_20_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14397__567 clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 net2036 sky130_fd_sc_hd__inv_2
XANTENNA__10008__A0 _03822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11122__C net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10559__A1 _05664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10559__B2 _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11756__B1 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07975__A2 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout404 net405 vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__clkbuf_4
XFILLER_99_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_165_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout415 net416 vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12181__B1 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout426 _06756_ vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__clkbuf_8
Xfanout437 _06467_ vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__buf_4
X_09823_ net698 _05458_ _05459_ net638 vssd1 vssd1 vccd1 vccd1 _05462_ sky130_fd_sc_hd__a31o_1
XFILLER_86_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout459 net463 vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__clkbuf_4
XFILLER_100_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15950__RESET_B net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout387_A net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09754_ net708 _05370_ _05373_ vssd1 vssd1 vccd1 vccd1 _05393_ sky130_fd_sc_hd__or3_1
XFILLER_100_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08705_ net784 _04337_ _04338_ vssd1 vssd1 vccd1 vccd1 _04344_ sky130_fd_sc_hd__and3_1
XANTENNA__10041__Y _05680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09685_ top.CPU.registers.data\[249\] net1394 net837 top.CPU.registers.data\[217\]
+ net732 vssd1 vssd1 vccd1 vccd1 _05324_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout554_A _02847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout175_X net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_93_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_93_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08152__A2 net1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1296_A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_169_Left_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_126_Right_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08636_ net706 _04273_ _04274_ _04268_ _04272_ vssd1 vssd1 vccd1 vccd1 _04275_ sky130_fd_sc_hd__o32a_1
X_13842__12 clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 net1481 sky130_fd_sc_hd__inv_2
XANTENNA__12236__A1 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14341__511 clknet_leaf_112_clk vssd1 vssd1 vccd1 vccd1 net1980 sky130_fd_sc_hd__inv_2
XANTENNA_fanout342_X net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08567_ top.CPU.registers.data\[751\] net1388 net812 top.CPU.registers.data\[719\]
+ net717 vssd1 vssd1 vccd1 vccd1 _04206_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout721_A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14638__808 clknet_leaf_165_clk vssd1 vssd1 vccd1 vccd1 net2277 sky130_fd_sc_hd__inv_2
XANTENNA_fanout819_A net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07518_ net1409 net1408 top.CPU.control_unit.instruction\[6\] top.CPU.control_unit.instruction\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03157_ sky130_fd_sc_hd__and4b_4
XFILLER_147_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08498_ net794 _04126_ _04127_ net721 vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__o211a_1
XFILLER_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11995__B1 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout607_X net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10460_ net3490 net226 net316 _06086_ vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__a22o_1
XANTENNA__09404__A2 net1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11747__B1 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09119_ top.CPU.registers.data\[807\] top.CPU.registers.data\[775\] net834 vssd1
+ vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__mux2_1
X_10391_ _06015_ _06019_ vssd1 vssd1 vccd1 vccd1 _06020_ sky130_fd_sc_hd__nor2_1
XANTENNA__13020__S net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12130_ top.CPU.registers.data\[87\] net651 net362 vssd1 vssd1 vccd1 vccd1 _06833_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__11762__A3 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout976_X net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12144__B net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10970__B2 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12061_ net566 net363 _06609_ _06799_ _06798_ vssd1 vssd1 vccd1 vccd1 _01533_ sky130_fd_sc_hd__a41o_1
XFILLER_1_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold480 top.CPU.registers.data\[164\] vssd1 vssd1 vccd1 vccd1 net3037 sky130_fd_sc_hd__dlygate4sd3_1
Xhold491 _02604_ vssd1 vssd1 vccd1 vccd1 net3048 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08915__A1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12172__B1 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11012_ net541 net501 _06355_ vssd1 vssd1 vccd1 vccd1 _06562_ sky130_fd_sc_hd__or3b_1
XFILLER_49_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout960 net961 vssd1 vssd1 vccd1 vccd1 net960 sky130_fd_sc_hd__clkbuf_4
X_15820_ net2154 _02030_ net1071 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[620\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout971 net973 vssd1 vssd1 vccd1 vccd1 net971 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout982 net985 vssd1 vssd1 vccd1 vccd1 net982 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08128__C1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout993 net994 vssd1 vssd1 vccd1 vccd1 net993 sky130_fd_sc_hd__buf_2
XFILLER_46_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15751_ net2085 _01961_ net1201 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[551\]
+ sky130_fd_sc_hd__dfrtp_1
X_12963_ net1411 top.I2C.bit_timer_state\[0\] vssd1 vssd1 vccd1 vccd1 _07401_ sky130_fd_sc_hd__nand2_1
XANTENNA__11278__A2 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08679__B1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13672__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_84_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_clk sky130_fd_sc_hd__clkbuf_8
Xhold1180 top.mmio.mem_data_i\[21\] vssd1 vssd1 vccd1 vccd1 net3737 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1191 top.CPU.registers.data\[748\] vssd1 vssd1 vccd1 vccd1 net3748 sky130_fd_sc_hd__dlygate4sd3_1
X_11914_ net3558 net187 net345 _06107_ vssd1 vssd1 vccd1 vccd1 _01652_ sky130_fd_sc_hd__a22o_1
X_15682_ net2016 _01892_ net1172 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[482\]
+ sky130_fd_sc_hd__dfrtp_1
X_12894_ top.CPU.alu.program_counter\[25\] _05362_ vssd1 vssd1 vccd1 vccd1 _07339_
+ sky130_fd_sc_hd__and2_1
XANTENNA__07541__X _03180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13424__A0 net1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11845_ _06676_ net200 net153 net3087 vssd1 vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__a22o_1
X_14084__254 clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 net1723 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07701__B net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ _06619_ net205 net162 net3177 vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__a22o_1
XANTENNA__10789__A1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16303_ clknet_leaf_107_clk _02512_ net1248 vssd1 vssd1 vccd1 vccd1 top.CPU.data_out\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11986__B1 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13515_ _03369_ net584 net589 vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__o21ai_1
X_10727_ _05712_ _05752_ _06139_ net412 vssd1 vssd1 vccd1 vccd1 _06341_ sky130_fd_sc_hd__o22a_1
XANTENNA__11450__A2 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14125__295 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 net1764 sky130_fd_sc_hd__inv_2
XFILLER_174_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16234_ clknet_leaf_43_clk _02444_ net1117 vssd1 vssd1 vccd1 vccd1 top.CPU.control_unit.instruction\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_146_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13446_ net3805 _02944_ net123 vssd1 vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__mux2_1
X_10658_ _04665_ net508 net503 _04664_ net443 vssd1 vssd1 vccd1 vccd1 _06275_ sky130_fd_sc_hd__o221a_1
XFILLER_127_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload14 clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clkload14/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__11738__B1 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload25 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 clkload25/Y sky130_fd_sc_hd__inv_8
XFILLER_103_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16165_ net2499 _02375_ net1083 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[965\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload36 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 clkload36/Y sky130_fd_sc_hd__inv_16
X_13377_ net1344 top.mmio.mem_data_i\[19\] net597 vssd1 vssd1 vccd1 vccd1 _02901_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__09628__B _05266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload47 clknet_leaf_192_clk vssd1 vssd1 vccd1 vccd1 clkload47/Y sky130_fd_sc_hd__inv_16
X_10589_ net444 _06209_ _06208_ _06195_ vssd1 vssd1 vccd1 vccd1 _06210_ sky130_fd_sc_hd__o211ai_4
Xclkload58 clknet_leaf_178_clk vssd1 vssd1 vccd1 vccd1 clkload58/Y sky130_fd_sc_hd__clkinv_8
Xclkload69 clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 clkload69/Y sky130_fd_sc_hd__inv_16
XFILLER_142_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15116_ net1498 _01329_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r2_prev\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07957__A2 net1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12328_ net3058 _04461_ net1157 vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__mux2_1
XFILLER_154_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16096_ net2430 _02306_ net1092 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[896\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_154_495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12054__B _06731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10961__B2 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15047_ clknet_leaf_92_clk _01292_ net1268 vssd1 vssd1 vccd1 vccd1 top.SPI.command\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_12259_ net3095 _06230_ net431 vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__mux2_1
XFILLER_69_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12163__B1 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07709__A2 net1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14782__952 clknet_leaf_153_clk vssd1 vssd1 vccd1 vccd1 net2421 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_143_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11910__B1 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08382__A2 _04019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09363__B net1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07590__B1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_160_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12466__A1 _03610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09867__C1 _03650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12466__B2 _05361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15949_ net2283 _02159_ net1069 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[749\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_75_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_clk sky130_fd_sc_hd__clkbuf_8
X_14823__993 clknet_leaf_185_clk vssd1 vssd1 vccd1 vccd1 net2462 sky130_fd_sc_hd__inv_2
XANTENNA__10302__B net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13989__159 clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 net1628 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_121_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09470_ top.CPU.registers.data\[834\] net1324 net855 top.CPU.registers.data\[866\]
+ net748 vssd1 vssd1 vccd1 vccd1 _05109_ sky130_fd_sc_hd__a221o_1
XFILLER_24_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08694__S net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08421_ _03925_ _04055_ _04058_ _04059_ vssd1 vssd1 vccd1 vccd1 _04060_ sky130_fd_sc_hd__o211a_1
XFILLER_51_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09619__C1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08352_ top.CPU.registers.data\[946\] top.CPU.registers.data\[914\] top.CPU.registers.data\[818\]
+ top.CPU.registers.data\[786\] net818 net720 vssd1 vssd1 vccd1 vccd1 _03991_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_158_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11977__B1 net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08283_ _03920_ _03921_ vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__nor2_1
XFILLER_20_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout135_A _05879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload8 clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clkload8/Y sky130_fd_sc_hd__inv_6
XFILLER_165_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08723__A _04361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11729__B1 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09398__A1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10464__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout302_A _06604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1044_A _03165_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10401__B1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09493__S1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07948__A2 net1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11744__A3 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10952__B2 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08869__S net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1211_A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12154__B1 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout201 net202 vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1309_A net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout212 _06752_ vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08358__C1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout223 _06469_ vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__buf_4
XANTENNA_fanout671_A _00000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout234 net243 vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__buf_4
Xfanout245 _06748_ vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout292_X net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout256 _06728_ vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout769_A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13933__103 clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 net1572 sky130_fd_sc_hd__inv_2
X_09806_ top.CPU.registers.data\[442\] net1395 net837 top.CPU.registers.data\[410\]
+ net698 vssd1 vssd1 vccd1 vccd1 _05445_ sky130_fd_sc_hd__a221o_1
Xfanout267 net270 vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10052__X _05691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout278 net279 vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__clkbuf_8
XFILLER_87_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout289 net292 vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__buf_6
X_07998_ top.CPU.registers.data\[408\] net983 _03636_ vssd1 vssd1 vccd1 vccd1 _03637_
+ sky130_fd_sc_hd__a21o_1
XFILLER_101_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12411__C top.CPU.addressnew\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09737_ top.CPU.registers.data\[251\] net1391 net827 top.CPU.registers.data\[219\]
+ net775 vssd1 vssd1 vccd1 vccd1 _05376_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout936_A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10212__B _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12457__B2 _03575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_66_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1299_X net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14068__238 clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 net1707 sky130_fd_sc_hd__inv_2
X_09668_ top.CPU.registers.data\[665\] net1336 net869 top.CPU.registers.data\[697\]
+ net710 vssd1 vssd1 vccd1 vccd1 _05307_ sky130_fd_sc_hd__a221o_1
XANTENNA__08530__C1 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08619_ _04225_ _04257_ vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__nor2_1
XANTENNA__13406__B1 net1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09599_ top.CPU.registers.data\[32\] top.CPU.registers.data\[0\] net810 vssd1 vssd1
+ vccd1 vccd1 _05238_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout724_X net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11680__A2 _06500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10866__C _06471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11630_ _05695_ net208 net427 net3592 vssd1 vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__a22o_1
X_14109__279 clknet_leaf_130_clk vssd1 vssd1 vccd1 vccd1 net1748 sky130_fd_sc_hd__inv_2
XFILLER_145_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11968__B1 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07636__B2 _03152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08833__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11561_ _06673_ net261 net248 net3182 vssd1 vssd1 vccd1 vccd1 _01975_ sky130_fd_sc_hd__a22o_1
XANTENNA__11432__A2 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13300_ _02832_ _02833_ _02836_ _02842_ vssd1 vssd1 vccd1 vccd1 _02843_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_42_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10512_ net392 _06040_ vssd1 vssd1 vccd1 vccd1 _06136_ sky130_fd_sc_hd__or2_1
XANTENNA__10640__B1 _05685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11492_ _06622_ net258 net255 net3608 vssd1 vssd1 vccd1 vccd1 _02032_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_21_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13231_ _02785_ _02793_ vssd1 vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__nor2_1
XFILLER_155_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10443_ _06021_ _06068_ net310 vssd1 vssd1 vccd1 vccd1 _06070_ sky130_fd_sc_hd__mux2_1
XFILLER_109_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08597__C1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13162_ top.I2C.output_state\[6\] top.I2C.output_state\[19\] top.I2C.output_state\[23\]
+ top.I2C.scl_out vssd1 vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__or4b_1
X_10374_ _05687_ _06000_ _06001_ _06002_ _06003_ vssd1 vssd1 vccd1 vccd1 _06004_ sky130_fd_sc_hd__o311a_1
X_12113_ net3964 net176 _06824_ _06641_ vssd1 vssd1 vccd1 vccd1 _01506_ sky130_fd_sc_hd__a22o_1
XFILLER_124_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14766__936 clknet_leaf_165_clk vssd1 vssd1 vccd1 vccd1 net2405 sky130_fd_sc_hd__inv_2
X_13093_ top.CPU.data_out\[28\] net2785 net560 vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__mux2_1
XANTENNA__08779__S net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12044_ _06593_ _06779_ _06781_ net3099 vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__a22o_1
XANTENNA__09010__B1 net1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11499__A2 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_88_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14510__680 clknet_leaf_165_clk vssd1 vssd1 vccd1 vccd1 net2149 sky130_fd_sc_hd__inv_2
XANTENNA__12160__A3 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14807__977 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 net2446 sky130_fd_sc_hd__inv_2
XANTENNA__10171__A2 _05806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07572__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout790 net791 vssd1 vssd1 vccd1 vccd1 net790 sky130_fd_sc_hd__clkbuf_2
X_15803_ net2137 _02013_ net1209 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[603\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11218__B net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09849__C1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_57_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08116__A2 _03754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15734_ net2068 _01944_ net1231 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[534\]
+ sky130_fd_sc_hd__dfrtp_1
X_12946_ _07366_ _07371_ _07375_ _07376_ _07384_ vssd1 vssd1 vccd1 vccd1 _07386_ sky130_fd_sc_hd__o311a_1
XFILLER_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15665_ net1999 _01875_ net1189 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[465\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12877_ _07322_ _07323_ vssd1 vssd1 vccd1 vccd1 _07324_ sky130_fd_sc_hd__nor2_1
XFILLER_34_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11234__A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11828_ _06661_ net500 net157 net3315 vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__a22o_1
X_15596_ net1930 _01806_ net1071 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[396\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08019__S net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11959__B1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12764__S net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11423__A2 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11759_ _06596_ net210 net195 net3017 vssd1 vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__a22o_1
XFILLER_174_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload103 clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 clkload103/Y sky130_fd_sc_hd__inv_6
Xclkload114 clknet_leaf_160_clk vssd1 vssd1 vccd1 vccd1 clkload114/Y sky130_fd_sc_hd__inv_4
X_16217_ net2551 _02427_ net1243 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[1017\]
+ sky130_fd_sc_hd__dfrtp_1
X_13429_ net3200 _02858_ net122 vssd1 vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__mux2_1
Xclkload125 clknet_leaf_166_clk vssd1 vssd1 vccd1 vccd1 clkload125/Y sky130_fd_sc_hd__inv_4
Xclkload136 clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 clkload136/Y sky130_fd_sc_hd__inv_12
XFILLER_60_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11187__A1 net1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload147 clknet_leaf_123_clk vssd1 vssd1 vccd1 vccd1 clkload147/Y sky130_fd_sc_hd__clkinv_8
Xclkload158 clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 clkload158/Y sky130_fd_sc_hd__inv_16
XFILLER_155_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload169 clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 clkload169/Y sky130_fd_sc_hd__inv_8
X_16148_ net2482 _02358_ net1120 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[948\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_114_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08970_ net783 _04607_ _04608_ net737 vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__o211a_1
X_16079_ net2413 _02289_ net1094 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[879\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_143_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09227__S1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12136__B1 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09374__A net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07921_ top.CPU.registers.data\[860\] net1302 net1023 top.CPU.registers.data\[892\]
+ net943 vssd1 vssd1 vccd1 vccd1 _03560_ sky130_fd_sc_hd__a221o_1
XFILLER_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07606__B net1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07852_ net674 _03486_ _03487_ _03490_ net610 vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__a311o_1
XFILLER_84_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput1 ACK_I vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07783_ top.CPU.registers.data\[670\] net1304 net1026 top.CPU.registers.data\[702\]
+ net628 vssd1 vssd1 vccd1 vccd1 _03422_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_48_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09304__A1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09522_ net758 _05160_ vssd1 vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__or2_1
XANTENNA__08277__X _03916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11111__A1 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09855__A2 net1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09453_ top.CPU.registers.data\[322\] net1324 net855 top.CPU.registers.data\[354\]
+ net773 vssd1 vssd1 vccd1 vccd1 _05092_ sky130_fd_sc_hd__a221o_1
XANTENNA__07866__A1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout252_A _06733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08404_ top.CPU.registers.data\[242\] net1378 net982 top.CPU.registers.data\[210\]
+ net908 vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__a221o_1
X_09384_ _05018_ _05021_ net454 vssd1 vssd1 vccd1 vccd1 _05023_ sky130_fd_sc_hd__mux2_2
XFILLER_51_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08335_ top.CPU.registers.data\[691\] top.CPU.registers.data\[659\] net989 vssd1
+ vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__mux2_1
XANTENNA__11414__A2 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08815__B1 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1161_A net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout517_A net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout138_X net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10622__A0 _04430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1259_A net1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08266_ top.CPU.registers.data\[598\] net1307 net1030 top.CPU.registers.data\[630\]
+ net947 vssd1 vssd1 vccd1 vccd1 _03905_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_134_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14453__623 clknet_leaf_171_clk vssd1 vssd1 vccd1 vccd1 net2092 sky130_fd_sc_hd__inv_2
X_08197_ net936 _03834_ _03835_ net954 vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__o211a_1
XANTENNA__08579__C1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_1001 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09240__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout886_A net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09791__A1 _05429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09284__A _04891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10090_ _03755_ net375 _05727_ vssd1 vssd1 vccd1 vccd1 _05728_ sky130_fd_sc_hd__o21ai_1
Xfanout1007 net1009 vssd1 vssd1 vccd1 vccd1 net1007 sky130_fd_sc_hd__buf_2
Xfanout1018 net1022 vssd1 vssd1 vccd1 vccd1 net1018 sky130_fd_sc_hd__clkbuf_4
Xfanout1029 net1031 vssd1 vssd1 vccd1 vccd1 net1029 sky130_fd_sc_hd__buf_2
XANTENNA_fanout674_X net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11319__A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout841_X net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout939_X net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_39_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_8
X_12800_ _07253_ vssd1 vssd1 vccd1 vccd1 _07254_ sky130_fd_sc_hd__inv_2
X_13780_ net8 net1049 net884 net3959 vssd1 vssd1 vccd1 vccd1 _02661_ sky130_fd_sc_hd__o22a_1
XFILLER_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10992_ net527 _06549_ vssd1 vssd1 vccd1 vccd1 _06550_ sky130_fd_sc_hd__nor2_1
XANTENNA__10877__B _05906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08503__C1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07532__A top.CPU.control_unit.instruction\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12731_ top.CPU.alu.program_counter\[10\] top.CPU.alu.program_counter\[9\] _07173_
+ vssd1 vssd1 vccd1 vccd1 _07191_ sky130_fd_sc_hd__and3_1
XFILLER_27_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11653__A2 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15450_ net1784 _01660_ net1252 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[250\]
+ sky130_fd_sc_hd__dfrtp_1
X_12662_ top.CPU.alu.program_counter\[2\] _07129_ net1359 vssd1 vssd1 vccd1 vccd1
+ _01165_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _06499_ net428 net206 net213 net2870 vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__a32o_1
X_15381_ net1715 _01591_ net1215 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[181\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11405__A2 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12593_ top.SPI.command\[3\] top.SPI.command\[2\] vssd1 vssd1 vccd1 vccd1 _07094_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__10893__A net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11544_ net489 net149 net356 net252 net2922 vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__a32o_1
XFILLER_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11475_ _06606_ net261 net257 net3272 vssd1 vssd1 vccd1 vccd1 _02048_ sky130_fd_sc_hd__a22o_1
X_14196__366 clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 net1835 sky130_fd_sc_hd__inv_2
X_16002_ net2336 _02212_ net1173 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[802\]
+ sky130_fd_sc_hd__dfrtp_1
X_13214_ net3810 _02779_ _02788_ _02773_ vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__a22o_1
X_10426_ net445 _06053_ _06052_ _06038_ vssd1 vssd1 vccd1 vccd1 _06054_ sky130_fd_sc_hd__o211a_2
XFILLER_152_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09231__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10916__A1 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09782__A1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13145_ net3867 top.CPU.data_out\[7\] net557 vssd1 vssd1 vccd1 vccd1 _01296_ sky130_fd_sc_hd__mux2_1
X_10357_ net446 _05969_ _05974_ net511 _05987_ vssd1 vssd1 vccd1 vccd1 _05988_ sky130_fd_sc_hd__a221oi_4
XFILLER_151_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13076_ top.CPU.data_out\[11\] net2756 net561 vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__mux2_1
X_10288_ _05617_ _05920_ vssd1 vssd1 vccd1 vccd1 _05921_ sky130_fd_sc_hd__nand2_1
XANTENNA__09534__A1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12027_ top.CPU.registers.data\[147\] _06781_ vssd1 vssd1 vccd1 vccd1 _06790_ sky130_fd_sc_hd__and2_1
XFILLER_93_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14935__RESET_B net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09298__B1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09837__A2 net1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09133__S net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12929_ _07348_ _07351_ _07357_ _07369_ _07356_ vssd1 vssd1 vccd1 vccd1 _07371_ sky130_fd_sc_hd__o311a_1
X_15717_ net2051 _01927_ net1062 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[517\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11644__A2 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_124_Left_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08972__S net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15648_ net1982 _01858_ net1090 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[448\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15579_ net1913 _01789_ net1214 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[379\]
+ sky130_fd_sc_hd__dfrtp_1
X_14140__310 clknet_leaf_138_clk vssd1 vssd1 vccd1 vccd1 net1779 sky130_fd_sc_hd__inv_2
XFILLER_147_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08120_ net917 _03758_ vssd1 vssd1 vccd1 vccd1 _03759_ sky130_fd_sc_hd__or2_1
X_14437__607 clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 net2076 sky130_fd_sc_hd__inv_2
XFILLER_174_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09470__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10080__A1 _04363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08051_ top.CPU.registers.data\[84\] net1288 net1008 top.CPU.registers.data\[116\]
+ net931 vssd1 vssd1 vccd1 vccd1 _03690_ sky130_fd_sc_hd__a221o_1
XANTENNA__10953__D net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08025__A1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11130__C _06213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10907__A1 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10027__B _05664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08576__A2 net1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11580__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07784__B1 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08953_ net617 _04591_ _04586_ _03342_ vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__o211a_1
XFILLER_131_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08328__A2 net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07904_ top.CPU.alu.program_counter\[28\] net1036 vssd1 vssd1 vccd1 vccd1 _03543_
+ sky130_fd_sc_hd__nor2_1
X_08884_ top.CPU.registers.data\[939\] top.CPU.registers.data\[907\] net805 vssd1
+ vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__mux2_1
XANTENNA__10135__A2 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1007_A net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07835_ top.CPU.registers.data_out_r1_prev\[29\] net873 net641 _03458_ _03473_ vssd1
+ vssd1 vccd1 vccd1 _03474_ sky130_fd_sc_hd__o221a_4
XANTENNA__12669__S net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10978__A net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11883__A2 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout467_A _03194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07766_ top.CPU.registers.data_out_r1_prev\[30\] net876 net638 _03404_ _03390_ vssd1
+ vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__o221ai_4
XANTENNA__09289__B1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09043__S net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10697__B _06311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09505_ top.CPU.registers.data\[737\] net1384 net1000 top.CPU.registers.data\[705\]
+ net921 vssd1 vssd1 vccd1 vccd1 _05144_ sky130_fd_sc_hd__a221o_1
XANTENNA__10189__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11635__A2 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout255_X net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07697_ net1047 _03262_ net1285 vssd1 vssd1 vccd1 vccd1 _03336_ sky130_fd_sc_hd__a21oi_2
XANTENNA_fanout1376_A net1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10843__B1 _06450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09436_ top.CPU.registers.data\[418\] top.CPU.registers.data\[386\] top.CPU.registers.data\[290\]
+ top.CPU.registers.data\[258\] net986 net911 vssd1 vssd1 vccd1 vccd1 _05075_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_23_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09367_ top.CPU.registers.data\[739\] net1381 net990 top.CPU.registers.data\[707\]
+ net915 vssd1 vssd1 vccd1 vccd1 _05006_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout801_A net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout422_X net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1164_X net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08318_ top.CPU.alu.program_counter\[19\] net878 vssd1 vssd1 vccd1 vccd1 _03957_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__08264__A1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09298_ top.CPU.registers.data\[740\] net1381 net992 top.CPU.registers.data\[708\]
+ net918 vssd1 vssd1 vccd1 vccd1 _04937_ sky130_fd_sc_hd__a221o_1
XFILLER_166_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08249_ _03887_ vssd1 vssd1 vccd1 vccd1 _03888_ sky130_fd_sc_hd__inv_2
XFILLER_153_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1331_X net1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11260_ net3175 net293 _06686_ net478 vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__a22o_1
XFILLER_137_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09213__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout791_X net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10211_ net602 _05845_ _05846_ vssd1 vssd1 vccd1 vccd1 _05847_ sky130_fd_sc_hd__a21o_4
XANTENNA__08567__A2 net1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13560__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13529__A _03854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11191_ net3534 net298 _06654_ net325 vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__a22o_1
XFILLER_122_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09218__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10142_ _05627_ _05635_ net305 vssd1 vssd1 vccd1 vccd1 _05779_ sky130_fd_sc_hd__mux2_1
XFILLER_97_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08319__A2 _03955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11049__A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14950_ clknet_leaf_52_clk _01196_ net1133 vssd1 vssd1 vccd1 vccd1 top.I2C.bit_timer_counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10073_ _05704_ _05710_ net386 vssd1 vssd1 vccd1 vccd1 _05711_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12115__A3 _06749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10126__A2 _05643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11323__B2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07961__S net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input28_A DAT_I[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14581__751 clknet_leaf_172_clk vssd1 vssd1 vccd1 vccd1 net2220 sky130_fd_sc_hd__inv_2
X_16620_ net1347 vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07533__Y _03172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09819__A2 net1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16551_ clknet_leaf_64_clk top.CPU.busy net1162 vssd1 vssd1 vccd1 vccd1 top.mmio.m1
+ sky130_fd_sc_hd__dfrtp_1
X_13763_ _03130_ top.wm.prev_BUSY_O net1050 vssd1 vssd1 vccd1 vccd1 _03094_ sky130_fd_sc_hd__and3_1
XFILLER_62_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11626__A2 _06701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10975_ net541 net501 _06057_ vssd1 vssd1 vccd1 vccd1 _06539_ sky130_fd_sc_hd__or3b_1
X_12714_ top.CPU.alu.program_counter\[8\] _04728_ vssd1 vssd1 vccd1 vccd1 _07176_
+ sky130_fd_sc_hd__nand2_1
X_14622__792 clknet_leaf_151_clk vssd1 vssd1 vccd1 vccd1 net2261 sky130_fd_sc_hd__inv_2
X_15502_ net1836 _01712_ net1107 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[302\]
+ sky130_fd_sc_hd__dfrtp_1
X_16482_ clknet_leaf_58_clk _02644_ net1143 vssd1 vssd1 vccd1 vccd1 top.I2C.which_data_address\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_71_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13694_ _03049_ _03051_ vssd1 vssd1 vccd1 vccd1 _02619_ sky130_fd_sc_hd__nor2_1
XANTENNA__11215__C net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15433_ net1767 _01643_ net1056 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[233\]
+ sky130_fd_sc_hd__dfrtp_1
X_12645_ _03135_ _06941_ vssd1 vssd1 vccd1 vccd1 _00020_ sky130_fd_sc_hd__nor2_1
XFILLER_157_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15364_ net1698 _01574_ net1221 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[164\]
+ sky130_fd_sc_hd__dfrtp_1
X_12576_ _07065_ _07076_ _07077_ _07080_ vssd1 vssd1 vccd1 vccd1 _07081_ sky130_fd_sc_hd__or4b_1
XANTENNA__12051__A2 _06779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11527_ _06652_ net258 net251 net3601 vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__a22o_1
XFILLER_156_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15295_ net1629 _01505_ net1223 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[95\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_156_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08007__A1 top.CPU.control_unit.instruction\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold309 top.CPU.registers.data\[17\] vssd1 vssd1 vccd1 vccd1 net2866 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09204__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11458_ net3807 net263 _06727_ net486 vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__a22o_1
XANTENNA__08380__X _04019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10409_ _05295_ _05964_ _03722_ _04056_ vssd1 vssd1 vccd1 vccd1 _06037_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_111_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11389_ net474 _06511_ net274 net3224 vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_74_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07766__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13128_ top.SPI.command\[2\] top.SPI.command\[4\] vssd1 vssd1 vccd1 vccd1 _02731_
+ sky130_fd_sc_hd__nor2_1
XFILLER_97_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09507__A1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13059_ top.SPI.parameters\[31\] top.SPI.paroutput\[23\] net1355 vssd1 vssd1 vccd1
+ vccd1 _07455_ sky130_fd_sc_hd__mux2_1
XFILLER_79_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1009 top.CPU.registers.data\[61\] vssd1 vssd1 vccd1 vccd1 net3566 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11314__B2 _06230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1360 net1362 vssd1 vssd1 vccd1 vccd1 net1360 sky130_fd_sc_hd__clkbuf_4
Xfanout1371 net1373 vssd1 vssd1 vccd1 vccd1 net1371 sky130_fd_sc_hd__clkbuf_4
Xfanout1382 net1383 vssd1 vssd1 vccd1 vccd1 net1382 sky130_fd_sc_hd__buf_2
XANTENNA__11865__A2 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1393 net1395 vssd1 vssd1 vccd1 vccd1 net1393 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08191__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07620_ top.CPU.control_unit.instruction\[14\] net1400 vssd1 vssd1 vccd1 vccd1 _03259_
+ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_109_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08268__A net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_132_Left_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07551_ net562 _03189_ vssd1 vssd1 vccd1 vccd1 _03190_ sky130_fd_sc_hd__nor2_4
XFILLER_35_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12248__A_N net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07482_ top.I2C.output_state\[26\] vssd1 vssd1 vccd1 vccd1 _03122_ sky130_fd_sc_hd__inv_2
XFILLER_62_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09221_ _04829_ _04857_ vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_17_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07900__A net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09152_ net683 _04782_ _04783_ net608 _04781_ vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__a311o_1
XANTENNA__12042__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12237__B net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08103_ net798 _03740_ _03741_ net752 vssd1 vssd1 vccd1 vccd1 _03742_ sky130_fd_sc_hd__o211a_1
XANTENNA__09994__A1 _04567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12952__S net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13790__A2 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09083_ top.CPU.registers.data\[584\] net1373 net970 top.CPU.registers.data\[616\]
+ net901 vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__o221a_1
XFILLER_163_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10038__A net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout215_A _06752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_141_Left_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08034_ top.CPU.registers.data\[564\] top.CPU.registers.data\[532\] net817 vssd1
+ vssd1 vccd1 vccd1 _03673_ sky130_fd_sc_hd__mux2_1
XANTENNA__09827__A _05465_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold810 top.CPU.registers.data\[378\] vssd1 vssd1 vccd1 vccd1 net3367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold821 top.CPU.registers.data\[263\] vssd1 vssd1 vccd1 vccd1 net3378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold832 top.CPU.registers.data\[527\] vssd1 vssd1 vccd1 vccd1 net3389 sky130_fd_sc_hd__dlygate4sd3_1
Xhold843 top.SPI.timem\[5\] vssd1 vssd1 vccd1 vccd1 net3400 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09746__A1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_171_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold854 top.CPU.registers.data\[687\] vssd1 vssd1 vccd1 vccd1 net3411 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold865 top.CPU.registers.data\[667\] vssd1 vssd1 vccd1 vccd1 net3422 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11553__A1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold876 top.CPU.registers.data\[207\] vssd1 vssd1 vccd1 vccd1 net3433 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap595 _02733_ vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__clkbuf_1
Xhold887 top.CPU.registers.data\[775\] vssd1 vssd1 vccd1 vccd1 net3444 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_168_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_51_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold898 top.CPU.registers.data\[138\] vssd1 vssd1 vccd1 vccd1 net3455 sky130_fd_sc_hd__dlygate4sd3_1
X_09985_ _05621_ _05623_ net381 vssd1 vssd1 vccd1 vccd1 _05624_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout584_A net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08936_ _04573_ _04574_ net928 vssd1 vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__mux2_1
XANTENNA__10108__A2 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14565__735 clknet_leaf_110_clk vssd1 vssd1 vccd1 vccd1 net2204 sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_186_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08706__C1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11305__B2 _06056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08867_ top.CPU.registers.data\[747\] net1386 net805 top.CPU.registers.data\[715\]
+ net761 vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout751_A net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11856__A2 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_150_Left_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_66_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout849_A net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07818_ net743 _03446_ _03447_ top.CPU.control_unit.instruction\[16\] vssd1 vssd1
+ vccd1 vccd1 _03457_ sky130_fd_sc_hd__a31o_1
XFILLER_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08798_ net1366 _04433_ _04436_ vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__o21a_1
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14606__776 clknet_leaf_164_clk vssd1 vssd1 vccd1 vccd1 net2245 sky130_fd_sc_hd__inv_2
X_07749_ _03386_ _03387_ net700 vssd1 vssd1 vccd1 vccd1 _03388_ sky130_fd_sc_hd__a21o_1
XFILLER_25_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1281_X net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout637_X net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1379_X net1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09131__C1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08485__A1 _04123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10760_ top.CPU.fetch.current_ra\[5\] net1040 net633 top.CPU.handler.toreg\[5\] _06372_
+ vssd1 vssd1 vccd1 vccd1 _06373_ sky130_fd_sc_hd__a221o_4
XFILLER_53_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09682__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08906__A net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09419_ net409 _05055_ vssd1 vssd1 vccd1 vccd1 _05058_ sky130_fd_sc_hd__nand2_1
XFILLER_73_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10691_ net446 _06306_ _06304_ _06301_ vssd1 vssd1 vccd1 vccd1 _06307_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout804_X net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13023__S net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10874__C net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_124_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12430_ _06894_ _06951_ vssd1 vssd1 vccd1 vccd1 _00058_ sky130_fd_sc_hd__nor2_1
XANTENNA__09434__B1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12033__A2 _06779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11051__B net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08788__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12361_ top.I2C.I2C_state\[19\] top.I2C.I2C_state\[13\] vssd1 vssd1 vccd1 vccd1 _06904_
+ sky130_fd_sc_hd__or2_1
XANTENNA__11241__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11312_ net3876 net290 _06709_ net492 vssd1 vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__a22o_1
X_15080_ clknet_leaf_55_clk _00018_ net1134 vssd1 vssd1 vccd1 vccd1 top.I2C.output_state\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12292_ net2582 _04223_ net1105 vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_139_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10890__B _05693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11243_ net2974 net294 _06676_ net314 vssd1 vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_91_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12741__A0 top.CPU.alu.program_counter\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11544__A1 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07748__B1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08945__C1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_19_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11174_ _03181_ net473 vssd1 vssd1 vccd1 vccd1 _06648_ sky130_fd_sc_hd__nor2_4
XFILLER_164_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10125_ net411 _05760_ _05762_ vssd1 vssd1 vccd1 vccd1 _05763_ sky130_fd_sc_hd__a21o_1
XFILLER_67_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15982_ net2316 _02192_ net1193 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[782\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14933_ clknet_leaf_71_clk _01179_ net1169 vssd1 vssd1 vccd1 vccd1 top.CPU.alu.program_counter\[16\]
+ sky130_fd_sc_hd__dfrtp_2
X_10056_ net1406 net576 net520 net138 vssd1 vssd1 vccd1 vccd1 _05695_ sky130_fd_sc_hd__and4_1
XANTENNA__11847__A2 _06678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08173__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09370__C1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08712__A2 net1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07704__B net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07920__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13815_ net3556 net337 net329 top.CPU.data_out\[17\] vssd1 vssd1 vccd1 vccd1 _02695_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10130__B _05767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13746_ net4004 _03082_ _03083_ vssd1 vssd1 vccd1 vccd1 _02639_ sky130_fd_sc_hd__o21a_1
X_16534_ clknet_leaf_99_clk net2972 net1256 vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08476__A1 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10958_ net519 net442 _05848_ net545 vssd1 vssd1 vccd1 vccd1 _06530_ sky130_fd_sc_hd__and4_1
XFILLER_32_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11480__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13677_ net2992 net331 net330 net4026 vssd1 vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__a22o_1
X_16465_ clknet_leaf_86_clk _02627_ net1265 vssd1 vssd1 vccd1 vccd1 top.SPI.timem\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10889_ net662 _06010_ _06471_ vssd1 vssd1 vccd1 vccd1 _06487_ sky130_fd_sc_hd__and3_1
XANTENNA__11242__A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12628_ net2780 top.I2C.I2C_state\[21\] _06901_ _07119_ vssd1 vssd1 vccd1 vccd1 top.I2C.sda_oeb_n
+ sky130_fd_sc_hd__or4_1
X_15416_ net1750 _01626_ net1148 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[216\]
+ sky130_fd_sc_hd__dfrtp_1
X_16396_ clknet_leaf_64_clk _00001_ net1162 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__12024__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15347_ net1681 _01557_ net1184 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[147\]
+ sky130_fd_sc_hd__dfrtp_1
X_12559_ _05806_ _05876_ _07063_ vssd1 vssd1 vccd1 vccd1 _07064_ sky130_fd_sc_hd__or3_1
XFILLER_129_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07987__B1 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13918__88 clknet_leaf_150_clk vssd1 vssd1 vccd1 vccd1 net1557 sky130_fd_sc_hd__inv_2
Xhold106 top.CPU.registers.data\[819\] vssd1 vssd1 vccd1 vccd1 net2663 sky130_fd_sc_hd__dlygate4sd3_1
X_15278_ net1612 _01488_ net1109 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[78\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold117 top.CPU.registers.data_out_r1_prev\[27\] vssd1 vssd1 vccd1 vccd1 net2674
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold128 top.CPU.registers.data\[313\] vssd1 vssd1 vccd1 vccd1 net2685 sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 top.CPU.registers.data\[927\] vssd1 vssd1 vccd1 vccd1 net2696 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12732__B1 top.CPU.alu.program_counter\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14252__422 clknet_leaf_190_clk vssd1 vssd1 vccd1 vccd1 net1891 sky130_fd_sc_hd__inv_2
Xfanout608 net609 vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__buf_4
XFILLER_99_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14549__719 clknet_leaf_170_clk vssd1 vssd1 vccd1 vccd1 net2188 sky130_fd_sc_hd__inv_2
Xfanout619 net623 vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_107_Right_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09770_ top.CPU.registers.data\[91\] net1297 net1018 top.CPU.registers.data\[123\]
+ net956 vssd1 vssd1 vccd1 vccd1 _05409_ sky130_fd_sc_hd__a221o_1
XANTENNA__08697__S net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10799__Y _06410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08721_ net702 _04356_ _04357_ _04358_ _04359_ vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__o32a_1
XFILLER_113_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11838__A2 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1190 net1192 vssd1 vssd1 vccd1 vccd1 net1190 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07614__B _03252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08652_ top.CPU.registers.data_out_r1_prev\[14\] net871 net644 _04275_ _04290_ vssd1
+ vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__o221ai_4
XFILLER_66_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07911__B1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07603_ top.CPU.alu.program_counter\[31\] _03241_ net1036 vssd1 vssd1 vccd1 vccd1
+ _03242_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_124_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08583_ _04201_ _04208_ _04214_ _04221_ vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__a22oi_4
XFILLER_82_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09113__C1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout165_A _06757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07534_ net1403 net572 vssd1 vssd1 vccd1 vccd1 _03173_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_141_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11066__A3 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10975__B net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07465_ top.CPU.control_unit.instruction\[6\] vssd1 vssd1 vccd1 vccd1 _03105_ sky130_fd_sc_hd__inv_2
XANTENNA__11471__B1 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout332_A _03047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1074_A net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09204_ top.CPU.registers.data\[838\] net1287 net1006 top.CPU.registers.data\[870\]
+ net930 vssd1 vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__a221o_1
XANTENNA__09416__A0 top.CPU.alu.program_counter\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12015__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09135_ top.CPU.registers.data\[39\] top.CPU.registers.data\[7\] net995 vssd1 vssd1
+ vccd1 vccd1 _04774_ sky130_fd_sc_hd__mux2_1
XANTENNA__11223__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10991__A _06190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1241_A net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout218_X net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09066_ top.CPU.registers.data\[40\] top.CPU.registers.data\[8\] net969 vssd1 vssd1
+ vccd1 vccd1 _04705_ sky130_fd_sc_hd__mux2_1
XFILLER_163_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09719__A1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout799_A net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08017_ top.CPU.registers.data\[180\] top.CPU.registers.data\[148\] net816 vssd1
+ vssd1 vccd1 vccd1 _03656_ sky130_fd_sc_hd__mux2_1
XFILLER_151_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold640 top.CPU.registers.data\[587\] vssd1 vssd1 vccd1 vccd1 net3197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold651 top.I2C.output_state\[4\] vssd1 vssd1 vccd1 vccd1 net3208 sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 top.CPU.registers.data\[682\] vssd1 vssd1 vccd1 vccd1 net3219 sky130_fd_sc_hd__dlygate4sd3_1
Xhold673 top.CPU.registers.data\[585\] vssd1 vssd1 vccd1 vccd1 net3230 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09195__A2 net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold684 top.CPU.registers.data\[530\] vssd1 vssd1 vccd1 vccd1 net3241 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10734__C1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold695 top.CPU.registers.data\[262\] vssd1 vssd1 vccd1 vccd1 net3252 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout966_A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08942__A2 net1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09968_ _05606_ vssd1 vssd1 vccd1 vccd1 _05607_ sky130_fd_sc_hd__inv_2
XANTENNA__12711__A top.CPU.alu.program_counter\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08919_ net636 _04554_ _04557_ vssd1 vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__or3_1
XFILLER_76_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09899_ _04430_ _04464_ vssd1 vssd1 vccd1 vccd1 _05538_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout754_X net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11829__A2 _06648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1340 top.CPU.handler.toreg\[0\] vssd1 vssd1 vccd1 vccd1 net3897 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13018__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1351 top.CPU.fetch.current_ra\[2\] vssd1 vssd1 vccd1 vccd1 net3908 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11930_ net3357 net185 net347 _06430_ vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__a22o_1
XFILLER_100_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1362 top.I2C.output_state\[15\] vssd1 vssd1 vccd1 vccd1 net3919 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1373 top.CPU.registers.data\[76\] vssd1 vssd1 vccd1 vccd1 net3930 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1384 top.CPU.registers.data\[72\] vssd1 vssd1 vccd1 vccd1 net3941 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1395 top.mmio.mem_data_i\[31\] vssd1 vssd1 vccd1 vccd1 net3952 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout921_X net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11861_ _06697_ net205 net153 net2678 vssd1 vssd1 vccd1 vccd1 _01700_ sky130_fd_sc_hd__a22o_1
XANTENNA__11046__B _06575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12857__S net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13600_ net1349 _06054_ vssd1 vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__nand2_1
XANTENNA__09104__C1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10812_ _05127_ _05269_ vssd1 vssd1 vccd1 vccd1 _06422_ sky130_fd_sc_hd__xnor2_1
XFILLER_60_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11057__A3 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11792_ _06640_ net208 net163 net3283 vssd1 vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__a22o_1
XFILLER_129_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10885__B net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13531_ _03645_ net585 vssd1 vssd1 vccd1 vccd1 _02986_ sky130_fd_sc_hd__and2_1
XANTENNA__11462__A0 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10743_ net526 _06356_ vssd1 vssd1 vccd1 vccd1 _06357_ sky130_fd_sc_hd__nor2_1
XANTENNA__11062__A _06190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16250_ clknet_leaf_61_clk _02460_ net1160 vssd1 vssd1 vccd1 vccd1 top.CPU.control_unit.instruction\[26\]
+ sky130_fd_sc_hd__dfrtp_2
X_14693__863 clknet_leaf_110_clk vssd1 vssd1 vccd1 vccd1 net2332 sky130_fd_sc_hd__inv_2
Xteam_08_1419 vssd1 vssd1 vccd1 vccd1 team_08_1419/HI gpio_oeb[5] sky130_fd_sc_hd__conb_1
X_13462_ net3997 _02952_ net120 vssd1 vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__mux2_1
XFILLER_174_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10674_ net438 _06290_ vssd1 vssd1 vccd1 vccd1 _06291_ sky130_fd_sc_hd__nand2_1
XFILLER_139_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15201_ net1535 _01411_ net1224 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12413_ top.CPU.addressnew\[15\] top.CPU.addressnew\[14\] _03133_ vssd1 vssd1 vccd1
+ vccd1 _06939_ sky130_fd_sc_hd__nand3_1
XANTENNA__09958__A1 _05332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16181_ net2515 _02391_ net1210 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[981\]
+ sky130_fd_sc_hd__dfrtp_1
X_13393_ net888 _02912_ vssd1 vssd1 vccd1 vccd1 _02913_ sky130_fd_sc_hd__and2_1
XFILLER_139_696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12962__B1 top.CPU.alu.program_counter\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15132_ clknet_leaf_48_clk _01342_ net1130 vssd1 vssd1 vccd1 vccd1 top.I2C.data_out\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_12344_ net3983 _06893_ net1054 vssd1 vssd1 vccd1 vccd1 _00043_ sky130_fd_sc_hd__o21a_1
XFILLER_126_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08091__C1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14236__406 clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 net1875 sky130_fd_sc_hd__inv_2
XFILLER_4_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15063_ clknet_leaf_49_clk _00066_ net1129 vssd1 vssd1 vccd1 vccd1 top.I2C.output_state\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_12275_ net3758 _03406_ net1240 vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__mux2_1
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10406__A net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11517__A1 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08918__C1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11226_ net521 _06532_ vssd1 vssd1 vccd1 vccd1 _06668_ sky130_fd_sc_hd__nor2_1
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12190__A1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08394__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11157_ net464 _06638_ vssd1 vssd1 vccd1 vccd1 _06639_ sky130_fd_sc_hd__and2_1
XFILLER_122_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10740__A2 _06352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10108_ _03613_ net379 _05745_ vssd1 vssd1 vccd1 vccd1 _05746_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11508__Y _06731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11088_ _03184_ _06598_ vssd1 vssd1 vccd1 vccd1 _06599_ sky130_fd_sc_hd__nor2_1
X_15965_ net2299 _02175_ net1113 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[765\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09343__C1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10039_ top.CPU.alu.immediate\[31\] net506 vssd1 vssd1 vccd1 vccd1 _05678_ sky130_fd_sc_hd__nand2_1
XFILLER_49_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15896_ net2230 _02106_ net1150 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[696\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_86_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11048__A3 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09110__A2 net1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11453__A0 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16517_ clknet_leaf_86_clk _02679_ net1265 vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__dfrtp_1
X_13729_ _03072_ _03073_ vssd1 vssd1 vccd1 vccd1 _02632_ sky130_fd_sc_hd__nor2_1
XANTENNA__10287__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16448_ clknet_leaf_81_clk _02611_ net1242 vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08980__S net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10008__A1 _03889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16379_ clknet_leaf_69_clk _02588_ net1165 vssd1 vssd1 vccd1 vccd1 top.CPU.fetch.current_ra\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11122__D net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12953__A0 top.CPU.alu.program_counter\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11756__A1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07609__B net1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08909__C1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09177__A2 net1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout405 _05024_ vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__buf_2
Xfanout416 _04957_ vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__clkbuf_4
Xfanout427 _06756_ vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__buf_4
X_09822_ top.CPU.registers.data\[474\] net1335 net867 top.CPU.registers.data\[506\]
+ net732 vssd1 vssd1 vccd1 vccd1 _05461_ sky130_fd_sc_hd__a221o_1
XANTENNA__13627__A net1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08924__A2 net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10603__X _06223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout438 net439 vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_126_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09753_ net696 _05388_ _05391_ vssd1 vssd1 vccd1 vccd1 _05392_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_126_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout282_A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09334__C1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08704_ net738 _04336_ net763 vssd1 vssd1 vccd1 vccd1 _04343_ sky130_fd_sc_hd__o21a_1
XANTENNA__11147__A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09684_ top.CPU.registers.data\[89\] net1336 net869 top.CPU.registers.data\[121\]
+ net757 vssd1 vssd1 vccd1 vccd1 _05323_ sky130_fd_sc_hd__a221o_1
XFILLER_66_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11692__A0 _06428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08635_ net792 _04264_ _04265_ vssd1 vssd1 vccd1 vccd1 _04274_ sky130_fd_sc_hd__and3_1
XANTENNA__07896__C1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10986__A net1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout168_X net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14380__550 clknet_leaf_189_clk vssd1 vssd1 vccd1 vccd1 net2019 sky130_fd_sc_hd__inv_2
XANTENNA_fanout1289_A net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08566_ top.CPU.registers.data\[591\] net1314 net845 top.CPU.registers.data\[623\]
+ net740 vssd1 vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__a221o_1
XFILLER_70_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14677__847 clknet_leaf_171_clk vssd1 vssd1 vccd1 vccd1 net2316 sky130_fd_sc_hd__inv_2
X_07517_ _03153_ _03155_ vssd1 vssd1 vccd1 vccd1 _03156_ sky130_fd_sc_hd__nand2_1
XFILLER_168_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08497_ net706 _04134_ _04135_ vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__or3_1
XFILLER_22_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout714_A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08860__A1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14421__591 clknet_leaf_171_clk vssd1 vssd1 vccd1 vccd1 net2060 sky130_fd_sc_hd__inv_2
X_14718__888 clknet_leaf_154_clk vssd1 vssd1 vccd1 vccd1 net2357 sky130_fd_sc_hd__inv_2
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout502_X net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09118_ net754 _04755_ _04756_ net700 vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__o211a_1
XANTENNA__08073__C1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10390_ _05733_ _05781_ _05790_ _05753_ _06018_ vssd1 vssd1 vccd1 vccd1 _06019_ sky130_fd_sc_hd__a221o_1
XFILLER_109_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09049_ top.CPU.registers.data\[296\] top.CPU.registers.data\[264\] net811 vssd1
+ vssd1 vccd1 vccd1 _04688_ sky130_fd_sc_hd__mux2_1
XFILLER_136_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10970__A2 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09168__A2 net1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12060_ top.CPU.registers.data\[123\] net653 vssd1 vssd1 vccd1 vccd1 _06799_ sky130_fd_sc_hd__or2_1
Xhold470 top.CPU.registers.data\[0\] vssd1 vssd1 vccd1 vccd1 net3027 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold481 top.SPI.paroutput\[16\] vssd1 vssd1 vccd1 vccd1 net3038 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout871_X net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout969_X net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08376__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold492 top.CPU.registers.data\[809\] vssd1 vssd1 vccd1 vccd1 net3049 sky130_fd_sc_hd__dlygate4sd3_1
X_11011_ net3621 net219 _06561_ net321 vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__a22o_1
XANTENNA__13537__A _05428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09573__C1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10722__A2 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout950 net951 vssd1 vssd1 vccd1 vccd1 net950 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07535__A net1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout961 net962 vssd1 vssd1 vccd1 vccd1 net961 sky130_fd_sc_hd__clkbuf_4
Xfanout972 net973 vssd1 vssd1 vccd1 vccd1 net972 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout983 net985 vssd1 vssd1 vccd1 vccd1 net983 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout994 net1003 vssd1 vssd1 vccd1 vccd1 net994 sky130_fd_sc_hd__clkbuf_4
XFILLER_161_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12962_ _07398_ _07400_ top.CPU.alu.program_counter\[31\] _03118_ vssd1 vssd1 vccd1
+ vccd1 _01194_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15750_ net2084 _01960_ net1081 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[550\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1170 top.CPU.registers.data\[201\] vssd1 vssd1 vccd1 vccd1 net3727 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13672__B2 top.CPU.addressnew\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input10_A DAT_I[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1181 top.SPI.paroutput\[12\] vssd1 vssd1 vccd1 vccd1 net3738 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09340__A2 net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11913_ net3442 net185 net347 _06086_ vssd1 vssd1 vccd1 vccd1 _01653_ sky130_fd_sc_hd__a22o_1
Xhold1192 top.CPU.registers.data\[921\] vssd1 vssd1 vccd1 vccd1 net3749 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11683__B1 net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12893_ _07336_ _07337_ vssd1 vssd1 vccd1 vccd1 _07338_ sky130_fd_sc_hd__nor2_1
X_15681_ net2015 _01891_ net1230 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[481\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11844_ net465 _06675_ net238 net154 net2681 vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__a32o_1
XANTENNA__12227__A2 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10238__A1 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11435__A0 _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11775_ net461 _06618_ net236 net161 net2857 vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__a32o_1
XFILLER_159_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16302_ clknet_leaf_107_clk _02511_ net1246 vssd1 vssd1 vccd1 vccd1 top.CPU.data_out\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10726_ _06000_ _06139_ _06339_ vssd1 vssd1 vccd1 vccd1 _06340_ sky130_fd_sc_hd__or3_1
X_13514_ _04188_ net584 vssd1 vssd1 vccd1 vccd1 _02977_ sky130_fd_sc_hd__and2_1
XFILLER_147_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08851__A1 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13445_ _02884_ _02937_ _02939_ vssd1 vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__a21o_1
X_16233_ clknet_leaf_33_clk _02443_ net1125 vssd1 vssd1 vccd1 vccd1 top.CPU.control_unit.instruction\[9\]
+ sky130_fd_sc_hd__dfrtp_4
X_10657_ _04730_ _05277_ _05279_ net370 vssd1 vssd1 vccd1 vccd1 _06274_ sky130_fd_sc_hd__a31o_1
XFILLER_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload15 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 clkload15/Y sky130_fd_sc_hd__inv_8
XFILLER_126_110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload26 clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 clkload26/Y sky130_fd_sc_hd__inv_12
X_13376_ top.CPU.control_unit.instruction\[18\] _02900_ net668 vssd1 vssd1 vccd1 vccd1
+ _02452_ sky130_fd_sc_hd__mux2_1
X_16164_ net2498 _02374_ net1210 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[964\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload37 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 clkload37/Y sky130_fd_sc_hd__inv_8
X_10588_ _04396_ _05568_ vssd1 vssd1 vccd1 vccd1 _06209_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09800__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload48 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 clkload48/Y sky130_fd_sc_hd__inv_8
Xclkload59 clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 clkload59/Y sky130_fd_sc_hd__inv_16
X_15115_ net1497 _01328_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r2_prev\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_86_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12327_ net2564 _04391_ net1157 vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__mux2_1
XFILLER_170_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16095_ net2429 _02305_ net1224 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[895\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_173_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10961__A2 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15046_ clknet_leaf_92_clk _01291_ net1268 vssd1 vssd1 vccd1 vccd1 top.SPI.command\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_12258_ net3141 _06212_ net431 vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__mux2_1
XANTENNA__12163__A1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09564__C1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11209_ net571 net487 _06660_ net299 net3425 vssd1 vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__a32o_1
X_12189_ net475 _06669_ _06861_ net170 net3549 vssd1 vssd1 vccd1 vccd1 _01467_ sky130_fd_sc_hd__a32o_1
XFILLER_150_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08975__S net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15948_ net2282 _02158_ net1070 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[748\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12466__A2 _03645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10302__C net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07732__X _03371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14364__534 clknet_leaf_137_clk vssd1 vssd1 vccd1 vccd1 net2003 sky130_fd_sc_hd__inv_2
XANTENNA__09331__A2 net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11674__B1 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07878__C1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15879_ net2213 _02089_ net1203 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[679\]
+ sky130_fd_sc_hd__dfrtp_1
X_08420_ _03858_ _03920_ _03857_ vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__a21boi_1
XFILLER_92_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12218__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09619__B1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08351_ top.CPU.alu.program_counter\[18\] net1033 vssd1 vssd1 vccd1 vccd1 _03990_
+ sky130_fd_sc_hd__or2_1
XANTENNA__11426__B1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14405__575 clknet_leaf_112_clk vssd1 vssd1 vccd1 vccd1 net2044 sky130_fd_sc_hd__inv_2
XFILLER_149_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_158_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08282_ _03889_ _03917_ vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__nor2_1
Xclkload9 clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clkload9/X sky130_fd_sc_hd__clkbuf_8
XFILLER_164_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11729__A1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout128_A net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11430__A net1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08055__C1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10952__A2 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08358__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout202 _06753_ vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__clkbuf_4
Xfanout213 _06752_ vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__buf_4
XFILLER_59_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout224 _05762_ vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__clkbuf_4
Xfanout235 net237 vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1204_A net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10704__A2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout246 net249 vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__buf_4
X_13972__142 clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 net1611 sky130_fd_sc_hd__inv_2
XFILLER_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13902__72 clknet_leaf_169_clk vssd1 vssd1 vccd1 vccd1 net1541 sky130_fd_sc_hd__inv_2
XANTENNA_input2_A DAT_I[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09805_ top.CPU.registers.data\[186\] net1394 net837 top.CPU.registers.data\[154\]
+ net710 vssd1 vssd1 vccd1 vccd1 _05444_ sky130_fd_sc_hd__a221o_1
Xfanout257 _06728_ vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__buf_2
Xfanout268 net270 vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__buf_4
Xfanout279 _06713_ vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__clkbuf_4
X_07997_ top.CPU.registers.data\[440\] net1010 net907 vssd1 vssd1 vccd1 vccd1 _03636_
+ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout664_A net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout285_X net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09307__C1 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09736_ net797 _05374_ vssd1 vssd1 vccd1 vccd1 _05375_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_2_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12457__A2 _03508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15418__RESET_B net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10468__A1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09322__A2 net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11665__B1 net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09667_ top.CPU.registers.data\[921\] net1336 net869 top.CPU.registers.data\[953\]
+ net698 vssd1 vssd1 vccd1 vccd1 _05306_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout452_X net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout831_A net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout929_A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08618_ _04255_ _04256_ net453 vssd1 vssd1 vccd1 vccd1 _04257_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_19_Left_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09598_ top.CPU.registers.data\[320\] net1313 net846 top.CPU.registers.data\[352\]
+ net766 vssd1 vssd1 vccd1 vccd1 _05237_ sky130_fd_sc_hd__a221o_1
XANTENNA__12209__A2 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07884__A2 net1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11680__A3 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11417__B1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08549_ net626 _04174_ _04176_ _04187_ vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__a31o_2
XANTENNA_fanout1361_X net1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09086__A1 _03116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout717_X net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11560_ net496 net475 _06672_ net249 net2665 vssd1 vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__a32o_1
XANTENNA__08294__C1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10511_ _06088_ _06134_ net306 vssd1 vssd1 vccd1 vccd1 _06135_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_42_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11491_ net562 net481 _06621_ net254 net3873 vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__a32o_1
XANTENNA__12436__A net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10882__C _06471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13230_ _02776_ net3265 _02798_ vssd1 vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__mux2_1
XFILLER_109_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire658 _03179_ vssd1 vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__clkbuf_4
X_10442_ _03684_ _03959_ net376 vssd1 vssd1 vccd1 vccd1 _06069_ sky130_fd_sc_hd__mux2_1
XANTENNA__09389__A2 net1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08125__S net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13161_ net3616 _02747_ _02749_ vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__a21o_1
X_10373_ _05721_ _05733_ _05754_ _05732_ vssd1 vssd1 vccd1 vccd1 _06003_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08061__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12112_ top.CPU.registers.data\[96\] net647 _06770_ vssd1 vssd1 vccd1 vccd1 _06824_
+ sky130_fd_sc_hd__o21a_1
XFILLER_152_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13092_ top.CPU.data_out\[27\] net2848 net561 vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__mux2_1
XFILLER_123_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13342__A0 top.CPU.control_unit.instruction\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12145__A1 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12043_ net3625 net151 _06793_ vssd1 vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__a21o_1
XFILLER_172_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09561__A2 net1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14051__221 clknet_leaf_114_clk vssd1 vssd1 vccd1 vccd1 net1690 sky130_fd_sc_hd__inv_2
XANTENNA__07572__A1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout780 net781 vssd1 vssd1 vccd1 vccd1 net780 sky130_fd_sc_hd__buf_4
X_14348__518 clknet_leaf_189_clk vssd1 vssd1 vccd1 vccd1 net1987 sky130_fd_sc_hd__inv_2
XFILLER_37_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15802_ net2136 _02012_ net1252 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[602\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout791 net794 vssd1 vssd1 vccd1 vccd1 net791 sky130_fd_sc_hd__buf_2
XFILLER_93_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11218__C _05771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11656__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15733_ net2067 _01943_ net1228 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[533\]
+ sky130_fd_sc_hd__dfrtp_1
X_12945_ _07366_ _07371_ _07375_ _07376_ vssd1 vssd1 vccd1 vccd1 _07385_ sky130_fd_sc_hd__o31a_1
XFILLER_45_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15664_ net1998 _01874_ net1156 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[464\]
+ sky130_fd_sc_hd__dfrtp_1
X_12876_ top.CPU.alu.program_counter\[23\] _07313_ vssd1 vssd1 vccd1 vccd1 _07323_
+ sky130_fd_sc_hd__nor2_1
XFILLER_34_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07875__A2 net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11671__A3 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11408__B1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11234__B _06010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11827_ net148 net3649 net157 vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__mux2_1
X_15595_ net1929 _01805_ net1067 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[395\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_159_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11758_ _06595_ net498 net192 net2956 vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__a22o_1
XANTENNA__12081__B1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10709_ net398 _06323_ net399 vssd1 vssd1 vccd1 vccd1 _06324_ sky130_fd_sc_hd__o21a_1
XFILLER_146_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11689_ _06513_ net198 net164 net3195 vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__a22o_1
Xclkload104 clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 clkload104/Y sky130_fd_sc_hd__clkinv_2
XFILLER_174_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16216_ net2550 _02426_ net1121 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[1016\]
+ sky130_fd_sc_hd__dfrtp_1
X_13428_ net4017 _02855_ net122 vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__mux2_1
Xclkload115 clknet_leaf_161_clk vssd1 vssd1 vccd1 vccd1 clkload115/Y sky130_fd_sc_hd__inv_8
Xclkload126 clknet_leaf_168_clk vssd1 vssd1 vccd1 vccd1 clkload126/Y sky130_fd_sc_hd__inv_6
Xclkload137 clknet_leaf_145_clk vssd1 vssd1 vccd1 vccd1 clkload137/Y sky130_fd_sc_hd__inv_16
XFILLER_115_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11187__A2 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload148 clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 clkload148/Y sky130_fd_sc_hd__inv_2
XANTENNA__09785__C1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload159 clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 clkload159/Y sky130_fd_sc_hd__inv_12
X_13359_ top.mmio.mem_data_i\[14\] _07089_ net554 top.I2C.data_out\[14\] vssd1 vssd1
+ vccd1 vccd1 _02888_ sky130_fd_sc_hd__a22o_1
X_16147_ net2481 _02357_ net1187 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[947\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_53_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08052__A2 net1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07874__S net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16078_ net2412 _02288_ net1106 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[878\]
+ sky130_fd_sc_hd__dfrtp_1
X_13956__126 clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 net1595 sky130_fd_sc_hd__inv_2
X_07920_ top.CPU.registers.data_out_r2_prev\[28\] net688 net621 _03552_ _03558_ vssd1
+ vssd1 vccd1 vccd1 _03559_ sky130_fd_sc_hd__o2111a_1
XANTENNA__10147__A0 _03407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15029_ clknet_leaf_90_clk _01274_ net1275 vssd1 vssd1 vccd1 vccd1 top.SPI.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_142_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11895__A0 _06428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07851_ net932 _03488_ _03489_ net952 vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__o211a_1
Xinput2 DAT_I[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
X_07782_ net920 _03418_ _03420_ vssd1 vssd1 vccd1 vccd1 _03421_ sky130_fd_sc_hd__and3_1
XFILLER_49_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09521_ top.CPU.registers.data\[801\] top.CPU.registers.data\[769\] net838 vssd1
+ vssd1 vccd1 vccd1 _05160_ sky130_fd_sc_hd__mux2_1
XANTENNA__11647__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07903__A _03541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11111__A2 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10967__C net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09452_ top.CPU.registers.data\[290\] top.CPU.registers.data\[258\] net823 vssd1
+ vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__mux2_1
XANTENNA__12020__S net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08403_ top.CPU.registers.data\[82\] net1291 net1012 top.CPU.registers.data\[114\]
+ net934 vssd1 vssd1 vccd1 vccd1 _04042_ sky130_fd_sc_hd__a221o_1
X_09383_ _05021_ vssd1 vssd1 vccd1 vccd1 _05022_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout245_A _06748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08334_ top.CPU.registers.data\[563\] top.CPU.registers.data\[531\] net989 vssd1
+ vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__mux2_1
XANTENNA__12072__B1 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10622__A1 _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08265_ net681 _03895_ _03896_ _03903_ net607 vssd1 vssd1 vccd1 vccd1 _03904_ sky130_fd_sc_hd__a311o_1
XANTENNA__10328__X _05960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16370__RESET_B net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08453__B net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08028__C1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08196_ top.CPU.registers.data\[663\] net1294 net1014 top.CPU.registers.data\[695\]
+ net912 vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__a221o_1
X_14492__662 clknet_leaf_135_clk vssd1 vssd1 vccd1 vccd1 net2131 sky130_fd_sc_hd__inv_2
XFILLER_146_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08579__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14789__959 clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 net2428 sky130_fd_sc_hd__inv_2
XANTENNA__12690__S net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout200_X net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10386__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08674__S0 net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1321_A net1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout781_A net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout879_A _03198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14035__205 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 net1674 sky130_fd_sc_hd__inv_2
X_13879__49 clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 net1518 sky130_fd_sc_hd__inv_2
XFILLER_120_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1008 net1009 vssd1 vssd1 vccd1 vccd1 net1008 sky130_fd_sc_hd__buf_2
XFILLER_126_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1019 net1022 vssd1 vssd1 vccd1 vccd1 net1019 sky130_fd_sc_hd__clkbuf_2
XFILLER_120_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11886__A0 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09543__A2 net1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11319__B net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11350__A2 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_27_Left_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11638__B1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09719_ net946 _05335_ _05336_ net960 vssd1 vssd1 vccd1 vccd1 _05358_ sky130_fd_sc_hd__o211a_1
XFILLER_16_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10991_ _06190_ net541 vssd1 vssd1 vccd1 vccd1 _06549_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout834_X net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13026__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08503__B1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09700__C1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10877__C _06471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12730_ top.CPU.alu.program_counter\[9\] _07190_ net1360 vssd1 vssd1 vccd1 vccd1
+ _01172_ sky130_fd_sc_hd__mux2_1
XFILLER_42_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07532__B net1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07857__A2 net1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12661_ _03100_ _07128_ net126 vssd1 vssd1 vccd1 vccd1 _07129_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11612_ net143 net3389 net213 vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08267__C1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12592_ top.SPI.command\[7\] top.SPI.command\[6\] vssd1 vssd1 vccd1 vccd1 _07093_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__08806__A1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15380_ net1714 _01590_ net1080 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[180\]
+ sky130_fd_sc_hd__dfrtp_1
X_14733__903 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 net2372 sky130_fd_sc_hd__inv_2
XFILLER_128_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11543_ net565 net491 _06660_ net252 net3288 vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__a32o_1
XANTENNA__11810__B1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_36_Left_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_98_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11474_ _06605_ net282 net257 net2938 vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_98_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13213_ net892 top.I2C.data_out\[22\] _02787_ vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__mux2_1
XFILLER_137_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16001_ net2335 _02211_ net1250 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[801\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_143_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10425_ _03723_ _05970_ vssd1 vssd1 vccd1 vccd1 _06053_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09767__C1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10916__A2 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13144_ net3904 top.CPU.data_out\[6\] net557 vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__mux2_1
X_10356_ _05983_ _05984_ _05986_ vssd1 vssd1 vccd1 vccd1 _05987_ sky130_fd_sc_hd__or3b_2
XFILLER_112_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07793__A1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13075_ top.CPU.data_out\[10\] net2792 net559 vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__mux2_1
XFILLER_112_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10287_ _05918_ _05919_ net401 vssd1 vssd1 vccd1 vccd1 _05920_ sky130_fd_sc_hd__mux2_1
XFILLER_105_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12026_ _06056_ net3456 net150 vssd1 vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__mux2_1
XANTENNA__11877__A0 _06056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11341__A2 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_45_Left_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09481__Y _05120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13893__63 clknet_leaf_109_clk vssd1 vssd1 vccd1 vccd1 net1532 sky130_fd_sc_hd__inv_2
XANTENNA__12453__A1_N _03405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15716_ net2050 _01926_ net1219 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[516\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_62_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12928_ _07348_ _07351_ _07357_ _07356_ vssd1 vssd1 vccd1 vccd1 _07370_ sky130_fd_sc_hd__o31a_1
XANTENNA__12775__S net1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15647_ net1981 _01857_ net1220 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[447\]
+ sky130_fd_sc_hd__dfrtp_1
X_12859_ top.CPU.alu.program_counter\[22\] _03916_ vssd1 vssd1 vccd1 vccd1 _07307_
+ sky130_fd_sc_hd__xor2_1
XFILLER_61_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15578_ net1912 _01788_ net1244 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[378\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_155_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14476__646 clknet_leaf_190_clk vssd1 vssd1 vccd1 vccd1 net2115 sky130_fd_sc_hd__inv_2
XANTENNA__11801__B1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08273__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08050_ top.CPU.registers.data\[148\] net979 _03688_ vssd1 vssd1 vccd1 vccd1 _03689_
+ sky130_fd_sc_hd__a21o_1
XFILLER_147_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14220__390 clknet_leaf_194_clk vssd1 vssd1 vccd1 vccd1 net1859 sky130_fd_sc_hd__inv_2
XANTENNA__13554__B1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14517__687 clknet_leaf_173_clk vssd1 vssd1 vccd1 vccd1 net2156 sky130_fd_sc_hd__inv_2
XFILLER_143_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10907__A2 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09773__A2 net1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08981__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11580__A2 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08952_ _04587_ _04588_ _04589_ _04590_ net673 net902 vssd1 vssd1 vccd1 vccd1 _04591_
+ sky130_fd_sc_hd__mux4_1
XFILLER_102_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09525__A2 net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11868__A0 _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07903_ _03541_ vssd1 vssd1 vccd1 vccd1 _03542_ sky130_fd_sc_hd__inv_2
X_08883_ net786 _04520_ _04521_ net713 vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__o211a_1
XFILLER_57_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11332__A2 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07834_ _03469_ _03472_ net636 vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__a21o_1
XANTENNA__10978__B net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07765_ net700 _03402_ _03403_ _03400_ _03401_ vssd1 vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__o32a_1
XANTENNA_fanout362_A net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09504_ top.CPU.registers.data\[577\] net1305 net1028 top.CPU.registers.data\[609\]
+ net945 vssd1 vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__a221o_1
XFILLER_25_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07696_ top.CPU.registers.data\[575\] net999 vssd1 vssd1 vccd1 vccd1 _03335_ sky130_fd_sc_hd__or2_1
XFILLER_24_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09435_ net677 _05072_ _05073_ vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__and3_1
XFILLER_13_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout150_X net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10994__A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1271_A net1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout248_X net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout627_A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1369_A net1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09366_ top.CPU.registers.data\[579\] net1297 net1018 top.CPU.registers.data\[611\]
+ net939 vssd1 vssd1 vccd1 vccd1 _05005_ sky130_fd_sc_hd__a221o_1
XANTENNA__12045__B1 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11399__A2 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08317_ _03955_ vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__inv_2
XANTENNA__13793__B1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09461__A1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09297_ net680 _04934_ _04935_ net607 _04933_ vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__a311o_1
XANTENNA__10058__X _05696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout415_X net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08248_ net642 _03885_ _03886_ vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__o21ai_4
XANTENNA__08751__X _04390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13545__A0 top.CPU.data_out\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout996_A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09749__C1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08179_ net795 _03810_ _03817_ net643 vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__a211o_1
XANTENNA__12714__A top.CPU.alu.program_counter\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1324_X net1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10210_ top.CPU.fetch.current_ra\[28\] net1044 net882 top.CPU.handler.toreg\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05846_ sky130_fd_sc_hd__a22o_1
XFILLER_137_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11190_ net146 net429 vssd1 vssd1 vccd1 vccd1 _06654_ sky130_fd_sc_hd__and2_1
XFILLER_161_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11571__A2 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10141_ net394 _05776_ _05777_ vssd1 vssd1 vccd1 vccd1 _05778_ sky130_fd_sc_hd__o21ai_1
XFILLER_122_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10234__A net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10072_ net305 _05708_ _05709_ _05707_ vssd1 vssd1 vccd1 vccd1 _05710_ sky130_fd_sc_hd__o31ai_1
XANTENNA__11859__B1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11049__B _05694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout951_X net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11323__A2 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07543__A net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13831_ net3677 net336 _03096_ vssd1 vssd1 vccd1 vccd1 _02711_ sky130_fd_sc_hd__a21o_1
XFILLER_29_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16550_ clknet_leaf_64_clk net2559 net1164 vssd1 vssd1 vccd1 vccd1 top.mmio.s2 sky130_fd_sc_hd__dfrtp_1
XFILLER_16_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13762_ top.wm.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1 _03093_ sky130_fd_sc_hd__nand2_2
X_10974_ net3258 net218 _06538_ net317 vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__a22o_1
XANTENNA__08488__C1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11626__A3 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15501_ net1835 _01711_ net1076 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[301\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12713_ _07173_ _07174_ vssd1 vssd1 vccd1 vccd1 _07175_ sky130_fd_sc_hd__nor2_1
XFILLER_71_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16481_ clknet_leaf_58_clk _02643_ net1143 vssd1 vssd1 vccd1 vccd1 top.I2C.which_data_address\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_14163__333 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 net1802 sky130_fd_sc_hd__inv_2
X_13693_ _07113_ _03050_ vssd1 vssd1 vccd1 vccd1 _03051_ sky130_fd_sc_hd__nand2_1
XFILLER_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12036__B1 _06781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15432_ net1766 _01642_ net1066 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[232\]
+ sky130_fd_sc_hd__dfrtp_1
X_12644_ top.I2C.byte_manager_done net4016 vssd1 vssd1 vccd1 vccd1 _00002_ sky130_fd_sc_hd__and2_1
XFILLER_129_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12575_ _05988_ _07079_ vssd1 vssd1 vccd1 vccd1 _07080_ sky130_fd_sc_hd__and2_1
X_15363_ net1697 _01573_ net1212 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[163\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_129_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14204__374 clknet_leaf_139_clk vssd1 vssd1 vccd1 vccd1 net1843 sky130_fd_sc_hd__inv_2
XFILLER_7_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11526_ _06651_ net260 net252 net3316 vssd1 vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__a22o_1
XANTENNA__08660__C1 net1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15294_ net1628 _01504_ net1237 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[94\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12339__A1 _05154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13536__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11939__S net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_150_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11457_ net564 _06588_ vssd1 vssd1 vccd1 vccd1 _06727_ sky130_fd_sc_hd__and2_1
X_10408_ net3605 net226 net317 _06036_ vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__a22o_1
XANTENNA__11011__B2 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11388_ net482 net471 _06507_ net271 net3210 vssd1 vssd1 vccd1 vccd1 _02122_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_74_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13127_ _07094_ _02727_ _02729_ top.SPI.command\[1\] vssd1 vssd1 vccd1 vccd1 _02730_
+ sky130_fd_sc_hd__and4b_1
X_10339_ _05575_ _05577_ _05588_ vssd1 vssd1 vccd1 vccd1 _05970_ sky130_fd_sc_hd__o21ai_1
X_13058_ net3596 _07454_ net894 vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__mux2_1
XFILLER_78_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11314__A2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1350 net1352 vssd1 vssd1 vccd1 vccd1 net1350 sky130_fd_sc_hd__clkbuf_4
X_12009_ _06578_ _06779_ _06781_ net3418 vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__a22o_1
XFILLER_94_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1361 net1362 vssd1 vssd1 vccd1 vccd1 net1361 sky130_fd_sc_hd__buf_4
XFILLER_16_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1372 net1373 vssd1 vssd1 vccd1 vccd1 net1372 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08810__S0 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08191__A1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1383 net1385 vssd1 vssd1 vccd1 vccd1 net1383 sky130_fd_sc_hd__buf_4
Xfanout1394 net1395 vssd1 vssd1 vccd1 vccd1 net1394 sky130_fd_sc_hd__buf_4
XANTENNA__11246__Y _06678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07550_ net648 _03186_ vssd1 vssd1 vccd1 vccd1 _03189_ sky130_fd_sc_hd__nand2_2
XANTENNA__11078__B2 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08479__C1 net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08983__S net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07481_ top.I2C.output_state\[7\] vssd1 vssd1 vccd1 vccd1 _03121_ sky130_fd_sc_hd__inv_2
XANTENNA__08494__A2 net1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09220_ _04829_ _04857_ vssd1 vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_17_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16274__Q top.CPU.handler.toreg\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09151_ net683 _04787_ _04788_ _04789_ vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_170_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09443__A1 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_8_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08102_ top.CPU.registers.data\[469\] net1330 net861 top.CPU.registers.data\[501\]
+ net777 vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__a221o_1
XANTENNA__10053__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09082_ top.CPU.registers.data\[712\] net1373 net969 top.CPU.registers.data\[744\]
+ net927 vssd1 vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__o221a_1
XANTENNA__11250__B2 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08033_ net705 _03670_ _03671_ _03669_ vssd1 vssd1 vccd1 vccd1 _03672_ sky130_fd_sc_hd__a31o_1
Xhold800 top.CPU.registers.data\[226\] vssd1 vssd1 vccd1 vccd1 net3357 sky130_fd_sc_hd__dlygate4sd3_1
Xhold811 top.I2C.data_out\[26\] vssd1 vssd1 vccd1 vccd1 net3368 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12534__A _03650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout208_A net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09319__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold822 top.CPU.registers.data\[331\] vssd1 vssd1 vccd1 vccd1 net3379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold833 top.CPU.registers.data\[23\] vssd1 vssd1 vccd1 vccd1 net3390 sky130_fd_sc_hd__dlygate4sd3_1
Xhold844 top.CPU.registers.data\[251\] vssd1 vssd1 vccd1 vccd1 net3401 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08403__C1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08223__S net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold855 top.CPU.registers.data\[792\] vssd1 vssd1 vccd1 vccd1 net3412 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold866 top.CPU.registers.data\[820\] vssd1 vssd1 vccd1 vccd1 net3423 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11553__A2 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold877 top.CPU.registers.data\[200\] vssd1 vssd1 vccd1 vccd1 net3434 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_168_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold888 top.CPU.registers.data\[269\] vssd1 vssd1 vccd1 vccd1 net3445 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10054__A net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09984_ _05546_ _05622_ vssd1 vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__nor2_1
Xhold899 top.CPU.registers.data\[148\] vssd1 vssd1 vccd1 vccd1 net3456 sky130_fd_sc_hd__dlygate4sd3_1
X_13849__19 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 net1488 sky130_fd_sc_hd__inv_2
X_08935_ top.CPU.registers.data\[170\] top.CPU.registers.data\[138\] net972 vssd1
+ vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__mux2_1
XANTENNA__10989__A net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout198_X net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout577_A _03169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11305__A2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08866_ top.CPU.registers.data\[683\] top.CPU.registers.data\[651\] net813 vssd1
+ vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__mux2_1
XFILLER_57_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07817_ net705 _03450_ _03451_ net719 vssd1 vssd1 vccd1 vccd1 _03456_ sky130_fd_sc_hd__o211a_1
X_08797_ net1283 _04434_ _04435_ vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__or3_1
XFILLER_45_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout365_X net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout744_A net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14147__317 clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 net1786 sky130_fd_sc_hd__inv_2
X_07748_ top.CPU.registers.data\[862\] net1333 net863 top.CPU.registers.data\[894\]
+ net754 vssd1 vssd1 vccd1 vccd1 _03387_ sky130_fd_sc_hd__a221o_1
XANTENNA__08893__S net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07679_ _03298_ _03304_ vssd1 vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout911_A net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout532_X net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09682__A1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09418_ net409 _05055_ vssd1 vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__or2_1
X_10690_ _05277_ _06305_ vssd1 vssd1 vccd1 vccd1 _06306_ sky130_fd_sc_hd__and2_1
XFILLER_12_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09349_ net416 _04987_ vssd1 vssd1 vccd1 vccd1 _04988_ sky130_fd_sc_hd__and2_1
XANTENNA__08237__A2 net1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12360_ _06902_ vssd1 vssd1 vccd1 vccd1 _06903_ sky130_fd_sc_hd__inv_2
XFILLER_138_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11241__A1 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08642__C1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14869__1039 clknet_leaf_172_clk vssd1 vssd1 vccd1 vccd1 net2508 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_95_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11311_ net477 net519 _05694_ _06499_ vssd1 vssd1 vccd1 vccd1 _06709_ sky130_fd_sc_hd__and4_1
XANTENNA__07996__A1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11792__A2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12291_ net3832 _04156_ net1235 vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__mux2_1
XFILLER_119_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10890__C _06010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11242_ net516 _06543_ vssd1 vssd1 vccd1 vccd1 _06676_ sky130_fd_sc_hd__nor2_1
XANTENNA__09737__A2 net1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_91_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11173_ net135 net3521 net299 vssd1 vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__mux2_1
XANTENNA__10752__B1 _06139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10124_ _05671_ _05761_ vssd1 vssd1 vccd1 vccd1 _05762_ sky130_fd_sc_hd__or2_2
XANTENNA__09753__A net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15981_ net2315 _02191_ net1076 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[781\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10899__A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10195__A1_N _03576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14932_ clknet_leaf_62_clk _01178_ net1164 vssd1 vssd1 vccd1 vccd1 top.CPU.alu.program_counter\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10055_ net552 _03180_ vssd1 vssd1 vccd1 vccd1 _05694_ sky130_fd_sc_hd__nand2_4
XANTENNA__11847__A3 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13425__D _07080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13863__33 clknet_leaf_159_clk vssd1 vssd1 vccd1 vccd1 net1502 sky130_fd_sc_hd__inv_2
X_13814_ net3142 net337 net329 top.CPU.data_out\[16\] vssd1 vssd1 vccd1 vccd1 _02694_
+ sky130_fd_sc_hd__a22o_1
XFILLER_29_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09122__B1 net1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16533_ clknet_leaf_85_clk _02695_ net1263 vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10807__A1 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13745_ top.SPI.timem\[20\] _03082_ _07113_ vssd1 vssd1 vccd1 vccd1 _03083_ sky130_fd_sc_hd__a21boi_1
X_10957_ net3600 net217 _06529_ net314 vssd1 vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__a22o_1
XFILLER_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12009__B1 _06781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16464_ clknet_leaf_86_clk _02626_ net1265 vssd1 vssd1 vccd1 vccd1 top.SPI.timem\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13676_ net3047 net331 net330 top.CPU.addressnew\[9\] vssd1 vssd1 vccd1 vccd1 _02604_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_14_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10888_ net488 net464 _06486_ net222 net3168 vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__a32o_1
XFILLER_32_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15415_ net1749 _01625_ net1183 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[215\]
+ sky130_fd_sc_hd__dfrtp_1
X_12627_ top.I2C.I2C_state\[8\] top.I2C.I2C_state\[11\] top.I2C.I2C_state\[9\] top.I2C.I2C_state\[10\]
+ vssd1 vssd1 vccd1 vccd1 _07119_ sky130_fd_sc_hd__or4_1
X_16395_ clknet_leaf_50_clk _00068_ net1131 vssd1 vssd1 vccd1 vccd1 top.I2C.initiate_read_bit
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08228__A2 net1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15346_ net1680 _01556_ net1099 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[146\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_156_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12558_ _05845_ _05904_ _05931_ _05958_ vssd1 vssd1 vccd1 vccd1 _07063_ sky130_fd_sc_hd__or4b_1
XANTENNA__11783__A2 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11509_ _06466_ _06731_ vssd1 vssd1 vccd1 vccd1 _06732_ sky130_fd_sc_hd__nor2_1
XANTENNA__10426__X _06054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15277_ net1611 _01487_ net1071 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[77\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10466__B1_N _05762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12489_ net449 _04727_ _04633_ _04658_ vssd1 vssd1 vccd1 vccd1 _06998_ sky130_fd_sc_hd__o2bb2a_1
Xhold107 top.CPU.registers.data\[62\] vssd1 vssd1 vccd1 vccd1 net2664 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold118 top.CPU.registers.data\[426\] vssd1 vssd1 vccd1 vccd1 net2675 sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 net118 vssd1 vssd1 vccd1 vccd1 net2686 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_153_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14291__461 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 net1930 sky130_fd_sc_hd__inv_2
XANTENNA__12732__A1 top.CPU.alu.program_counter\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11535__A2 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14588__758 clknet_leaf_139_clk vssd1 vssd1 vccd1 vccd1 net2227 sky130_fd_sc_hd__inv_2
XANTENNA__08400__A2 net1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout609 _03349_ vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__buf_4
XFILLER_39_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08720_ net738 _04350_ _04351_ net691 vssd1 vssd1 vccd1 vccd1 _04359_ sky130_fd_sc_hd__a31o_1
XANTENNA__11299__B2 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14629__799 clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 net2268 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_163_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1180 net1188 vssd1 vssd1 vccd1 vccd1 net1180 sky130_fd_sc_hd__clkbuf_4
X_08651_ _04282_ _04289_ net636 vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__a21o_1
Xfanout1191 net1192 vssd1 vssd1 vccd1 vccd1 net1191 sky130_fd_sc_hd__clkbuf_4
XFILLER_27_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07602_ _03097_ net875 net642 _03224_ _03240_ vssd1 vssd1 vccd1 vccd1 _03241_ sky130_fd_sc_hd__o221ai_4
XFILLER_26_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08582_ _04219_ _04220_ net703 vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_124_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09113__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07533_ net1405 net576 vssd1 vssd1 vccd1 vccd1 _03172_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_141_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08467__A2 net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout158_A net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07464_ net1408 vssd1 vssd1 vccd1 vccd1 _03104_ sky130_fd_sc_hd__inv_2
XANTENNA__11471__A1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09203_ top.CPU.registers.data_out_r2_prev\[6\] net685 net952 _04839_ _04841_ vssd1
+ vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__o2111a_1
XANTENNA__09416__A1 _05054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout325_A _03190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1067_A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09134_ net958 _04772_ _04771_ net943 vssd1 vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__o211a_1
XANTENNA__10026__A2 _03292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11223__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10991__B net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11774__A2 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09065_ net1366 _04700_ _04703_ vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__o21a_1
XFILLER_162_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09557__B net1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14532__702 clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 net2171 sky130_fd_sc_hd__inv_2
XFILLER_163_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09049__S net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08016_ top.CPU.registers.data\[84\] net1318 net849 top.CPU.registers.data\[116\]
+ net768 vssd1 vssd1 vccd1 vccd1 _03655_ sky130_fd_sc_hd__a221o_1
Xhold630 top.CPU.registers.data\[440\] vssd1 vssd1 vccd1 vccd1 net3187 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10055__Y _05694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold641 top.CPU.registers.data\[564\] vssd1 vssd1 vccd1 vccd1 net3198 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout694_A net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11526__A2 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold652 top.CPU.registers.data\[221\] vssd1 vssd1 vccd1 vccd1 net3209 sky130_fd_sc_hd__dlygate4sd3_1
Xhold663 top.CPU.registers.data\[515\] vssd1 vssd1 vccd1 vccd1 net3220 sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 top.CPU.registers.data\[713\] vssd1 vssd1 vccd1 vccd1 net3231 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1022_X net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1401_A net1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold685 top.CPU.registers.data\[33\] vssd1 vssd1 vccd1 vccd1 net3242 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10734__B1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold696 top.CPU.addressnew\[21\] vssd1 vssd1 vccd1 vccd1 net3253 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09967_ _03374_ _03445_ _05525_ _05605_ vssd1 vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout861_A net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout482_X net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout959_A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08918_ net787 _04555_ _04556_ net716 vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__o211a_1
XFILLER_103_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10512__A net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09898_ _04396_ _04468_ vssd1 vssd1 vccd1 vccd1 _05537_ sky130_fd_sc_hd__nor2_1
XANTENNA__11829__A3 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1330 top.CPU.registers.data\[759\] vssd1 vssd1 vccd1 vccd1 net3887 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09860__X _05499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1341 top.CPU.registers.data\[55\] vssd1 vssd1 vccd1 vccd1 net3898 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1352 top.CPU.registers.data\[997\] vssd1 vssd1 vccd1 vccd1 net3909 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1363 top.CPU.handler.toreg\[11\] vssd1 vssd1 vccd1 vccd1 net3920 sky130_fd_sc_hd__dlygate4sd3_1
X_08849_ top.CPU.registers.data\[203\] net1370 net967 top.CPU.registers.data\[235\]
+ net927 vssd1 vssd1 vccd1 vccd1 _04488_ sky130_fd_sc_hd__o221a_1
XFILLER_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1391_X net1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1374 top.I2C.data_out\[3\] vssd1 vssd1 vccd1 vccd1 net3931 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout747_X net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1385 top.CPU.registers.data\[106\] vssd1 vssd1 vccd1 vccd1 net3942 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1396 top.CPU.fetch.current_ra\[12\] vssd1 vssd1 vccd1 vccd1 net3953 sky130_fd_sc_hd__dlygate4sd3_1
X_11860_ _06696_ net204 net154 net2779 vssd1 vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__a22o_1
XFILLER_72_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10811_ net444 _05551_ _06420_ vssd1 vssd1 vccd1 vccd1 _06421_ sky130_fd_sc_hd__or3_1
XFILLER_14_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11791_ _06639_ net238 net162 net3538 vssd1 vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout914_X net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13034__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13530_ top.CPU.data_out\[23\] net589 net339 _02985_ vssd1 vssd1 vccd1 vccd1 _02521_
+ sky130_fd_sc_hd__o22a_1
X_10742_ net551 net501 _06355_ vssd1 vssd1 vccd1 vccd1 _06356_ sky130_fd_sc_hd__or3b_1
XFILLER_14_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11062__B _06575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10673_ net603 _06288_ _06289_ vssd1 vssd1 vccd1 vccd1 _06290_ sky130_fd_sc_hd__a21o_2
X_13461_ net1396 net872 _02905_ net418 vssd1 vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_173_Right_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15200_ net1534 _01410_ net1096 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12412_ top.CPU.addressnew\[0\] top.CPU.addressnew\[1\] top.CPU.addressnew\[19\]
+ top.CPU.addressnew\[18\] vssd1 vssd1 vccd1 vccd1 _06938_ sky130_fd_sc_hd__or4_1
XFILLER_138_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16180_ net2514 _02390_ net1112 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[980\]
+ sky130_fd_sc_hd__dfrtp_1
X_13392_ top.I2C.data_out\[23\] net556 _02911_ net597 vssd1 vssd1 vccd1 vccd1 _02912_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07969__A1 top.CPU.control_unit.instruction\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15131_ clknet_leaf_46_clk _01341_ net1137 vssd1 vssd1 vccd1 vccd1 top.I2C.data_out\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11765__A2 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12962__B2 _03118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12343_ top.I2C.output_state\[17\] _06892_ net1339 vssd1 vssd1 vccd1 vccd1 _06893_
+ sky130_fd_sc_hd__o21a_1
XFILLER_154_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14275__445 clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 net1914 sky130_fd_sc_hd__inv_2
XFILLER_142_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15062_ clknet_leaf_51_clk _00065_ net1132 vssd1 vssd1 vccd1 vccd1 top.I2C.output_state\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12274_ net2619 _03241_ net1203 vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__mux2_1
XFILLER_153_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10406__B net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11225_ net489 net466 _06667_ net295 net2949 vssd1 vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__a32o_1
XANTENNA__12902__A top.CPU.alu.program_counter\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14316__486 clknet_leaf_195_clk vssd1 vssd1 vccd1 vccd1 net1955 sky130_fd_sc_hd__inv_2
XANTENNA__08394__A1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12190__A2 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11156_ net574 net528 _06429_ vssd1 vssd1 vccd1 vccd1 _06638_ sky130_fd_sc_hd__and3_1
X_10107_ _03822_ net375 vssd1 vssd1 vccd1 vccd1 _05745_ sky130_fd_sc_hd__or2_1
X_11087_ net648 _03185_ vssd1 vssd1 vccd1 vccd1 _06598_ sky130_fd_sc_hd__nand2_1
XFILLER_67_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15964_ net2298 _02174_ net1195 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[764\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09343__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10038_ net506 vssd1 vssd1 vccd1 vccd1 _05677_ sky130_fd_sc_hd__inv_2
X_15895_ net2229 _02105_ net1180 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[695\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11150__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07731__A _03369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_170_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11989_ _06551_ net343 net180 net2822 vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__a22o_1
XANTENNA__11253__A net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16516_ clknet_leaf_92_clk _02678_ net1269 vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__dfrtp_1
X_13728_ top.SPI.timem\[13\] top.SPI.timem\[12\] _03068_ vssd1 vssd1 vccd1 vccd1 _03073_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08854__C1 net1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_50_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12068__B net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16447_ clknet_leaf_85_clk _02610_ net1263 vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__dfrtp_1
X_13659_ net2860 _07399_ net665 vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__mux2_1
XFILLER_83_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15536__RESET_B net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_140_Right_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_185_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16378_ clknet_leaf_62_clk _02587_ net1163 vssd1 vssd1 vccd1 vccd1 top.CPU.fetch.current_ra\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_129_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11756__A2 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15329_ net1663 _01539_ net1231 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[129\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10156__X _05793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_65_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08909__B1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09031__C1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout406 net407 vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__buf_2
XANTENNA_wire450_X net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12181__A2 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout417 _03242_ vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__clkbuf_4
X_09821_ top.CPU.registers.data\[346\] net1335 net867 top.CPU.registers.data\[378\]
+ net758 vssd1 vssd1 vccd1 vccd1 _05460_ sky130_fd_sc_hd__a221o_1
XFILLER_140_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout428 _06701_ vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__buf_4
XANTENNA_clkload12_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout439 _05697_ vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__buf_4
XFILLER_99_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07625__B top.CPU.control_unit.instruction\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09752_ net799 _05389_ _05390_ net751 vssd1 vssd1 vccd1 vccd1 _05391_ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_123_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_448 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13666__C1 _07089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08137__A1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09334__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08703_ net784 _04339_ _04340_ _04341_ net690 vssd1 vssd1 vccd1 vccd1 _04342_ sky130_fd_sc_hd__a311o_1
XFILLER_104_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09683_ net698 _05319_ _05320_ _05321_ vssd1 vssd1 vccd1 vccd1 _05322_ sky130_fd_sc_hd__a31o_1
XANTENNA__09885__A1 _03476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14868__1038 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 net2507 sky130_fd_sc_hd__inv_2
XANTENNA_fanout275_A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08634_ net744 _04261_ _04262_ net769 vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__o211a_1
XANTENNA__10986__B _03170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_138_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08565_ net740 _04202_ _04203_ net766 vssd1 vssd1 vccd1 vccd1 _04204_ sky130_fd_sc_hd__o211a_1
XANTENNA__09098__C1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout442_A _05697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11163__A net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10247__A2 _05367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07516_ top.CPU.control_unit.instruction\[3\] top.CPU.control_unit.instruction\[2\]
+ top.CPU.control_unit.instruction\[0\] top.CPU.control_unit.instruction\[1\] vssd1
+ vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__and4b_1
XANTENNA_clkbuf_leaf_18_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08496_ net793 _04130_ _04131_ net745 vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__o211a_1
XFILLER_168_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11995__A2 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout230_X net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_170_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_170_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08860__A2 _04497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout707_A net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14259__429 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 net1898 sky130_fd_sc_hd__inv_2
XANTENNA__08472__A net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11747__A2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09117_ top.CPU.registers.data\[647\] net1333 net864 top.CPU.registers.data\[679\]
+ net729 vssd1 vssd1 vccd1 vccd1 _04756_ sky130_fd_sc_hd__a221o_1
XANTENNA__09270__C1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09048_ top.CPU.registers.data\[72\] net1312 net843 top.CPU.registers.data\[104\]
+ net763 vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__a221o_1
X_14003__173 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 net1642 sky130_fd_sc_hd__inv_2
XFILLER_159_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout697_X net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold460 top.CPU.registers.data\[385\] vssd1 vssd1 vccd1 vccd1 net3017 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12722__A top.CPU.alu.program_counter\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold471 top.CPU.registers.data\[267\] vssd1 vssd1 vccd1 vccd1 net3028 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1404_X net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold482 top.CPU.fetch.current_ra\[4\] vssd1 vssd1 vccd1 vccd1 net3039 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08376__A1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11010_ net532 _06560_ vssd1 vssd1 vccd1 vccd1 _06561_ sky130_fd_sc_hd__nor2_1
XFILLER_89_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold493 top.SPI.parameters\[6\] vssd1 vssd1 vccd1 vccd1 net3050 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12172__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout864_X net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout940 net942 vssd1 vssd1 vccd1 vccd1 net940 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07584__C1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11380__B1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout951 net963 vssd1 vssd1 vccd1 vccd1 net951 sky130_fd_sc_hd__buf_4
XANTENNA__07535__B net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout962 net963 vssd1 vssd1 vccd1 vccd1 net962 sky130_fd_sc_hd__clkbuf_4
Xfanout973 net976 vssd1 vssd1 vccd1 vccd1 net973 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08128__A1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout984 net985 vssd1 vssd1 vccd1 vccd1 net984 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09325__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout995 net997 vssd1 vssd1 vccd1 vccd1 net995 sky130_fd_sc_hd__clkbuf_4
X_12961_ net128 _07399_ net1361 vssd1 vssd1 vccd1 vccd1 _07400_ sky130_fd_sc_hd__o21ai_1
XFILLER_161_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12868__S net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08679__A2 net1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14660__830 clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 net2299 sky130_fd_sc_hd__inv_2
Xhold1160 top.CPU.handler.toreg\[14\] vssd1 vssd1 vccd1 vccd1 net3717 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1171 top.CPU.registers.data\[127\] vssd1 vssd1 vccd1 vccd1 net3728 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1182 top.CPU.registers.data\[877\] vssd1 vssd1 vccd1 vccd1 net3739 sky130_fd_sc_hd__dlygate4sd3_1
X_11912_ net3972 net187 net344 _06058_ vssd1 vssd1 vccd1 vccd1 _01654_ sky130_fd_sc_hd__a22o_1
X_15680_ net2014 _01890_ net1090 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[480\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11683__A1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12892_ top.CPU.alu.program_counter\[25\] top.CPU.alu.program_counter\[24\] _07322_
+ vssd1 vssd1 vccd1 vccd1 _07337_ sky130_fd_sc_hd__and3_1
Xhold1193 top.CPU.registers.data\[492\] vssd1 vssd1 vccd1 vccd1 net3750 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07551__A net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11843_ _06674_ net235 net153 net3482 vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__a22o_1
XFILLER_72_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12227__A3 _06796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11073__A _06333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14701__871 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 net2340 sky130_fd_sc_hd__inv_2
XFILLER_13_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08836__C1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11774_ _06617_ net205 net162 net3174 vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_64_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ clknet_leaf_107_clk _02510_ net1248 vssd1 vssd1 vccd1 vccd1 top.CPU.data_out\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13513_ top.CPU.data_out\[15\] net588 _02969_ _02976_ vssd1 vssd1 vccd1 vccd1 _02513_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11986__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10725_ _05671_ _05759_ _06001_ vssd1 vssd1 vccd1 vccd1 _06339_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_161_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_161_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_81_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16232_ clknet_leaf_44_clk _02442_ net1126 vssd1 vssd1 vccd1 vccd1 top.CPU.control_unit.instruction\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13444_ net3920 _02943_ net121 vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__mux2_1
X_10656_ _04730_ _05277_ _05279_ vssd1 vssd1 vccd1 vccd1 _06273_ sky130_fd_sc_hd__a21oi_1
XFILLER_173_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11738__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16163_ net2497 _02373_ net1206 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[963\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload16 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 clkload16/Y sky130_fd_sc_hd__inv_2
XFILLER_166_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10587_ _05643_ _05783_ _06205_ _06207_ vssd1 vssd1 vccd1 vccd1 _06208_ sky130_fd_sc_hd__o211a_1
X_13375_ _02830_ _02899_ vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__nor2_1
XFILLER_127_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08603__A2 net1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload27 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 clkload27/Y sky130_fd_sc_hd__clkinv_8
XFILLER_126_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload38 clknet_leaf_179_clk vssd1 vssd1 vccd1 vccd1 clkload38/Y sky130_fd_sc_hd__inv_4
Xclkload49 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 clkload49/Y sky130_fd_sc_hd__inv_2
X_15114_ net1496 _01327_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r2_prev\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_170_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12326_ net2606 _04324_ net1157 vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__mux2_1
X_16094_ net2428 _02304_ net1202 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[894\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_86_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15045_ clknet_leaf_94_clk _01290_ net1267 vssd1 vssd1 vccd1 vccd1 top.SPI.command\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_141_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09484__Y _05123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12699__B1 net1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09013__C1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12257_ net3140 _06191_ net431 vssd1 vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__mux2_1
XFILLER_107_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09564__B1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11208_ net147 net430 vssd1 vssd1 vccd1 vccd1 _06660_ sky130_fd_sc_hd__and2_1
X_12188_ top.CPU.registers.data\[57\] net656 _03185_ vssd1 vssd1 vccd1 vccd1 _06861_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__11371__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11910__A2 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11248__A net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11139_ net480 net457 _06628_ net301 net2697 vssd1 vssd1 vccd1 vccd1 _02284_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_143_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07590__A2 net1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15947_ net2281 _02157_ net1057 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[747\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11123__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11674__A1 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15878_ net2212 _02088_ net1081 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[678\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_121_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08350_ _03958_ _03987_ vssd1 vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__nand2_1
XANTENNA__11977__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08281_ _03919_ vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_152_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_152_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_20_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11729__A2 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08055__B1 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12154__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout203 net204 vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09327__S net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout214 _06752_ vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__buf_6
XANTENNA_fanout392_A net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11362__B1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout225 net228 vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__buf_6
Xfanout236 net237 vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__clkbuf_4
XFILLER_8_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout247 net249 vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__buf_4
X_09804_ net758 _05441_ _05442_ net644 vssd1 vssd1 vccd1 vccd1 _05443_ sky130_fd_sc_hd__a31o_1
Xfanout258 net259 vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__buf_4
XANTENNA__10062__A _05123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14644__814 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 net2283 sky130_fd_sc_hd__inv_2
Xfanout269 net270 vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__clkbuf_8
X_07996_ net675 _03630_ _03631_ _03634_ net610 vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__a311o_1
XFILLER_28_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09735_ top.CPU.registers.data\[187\] top.CPU.registers.data\[155\] net827 vssd1
+ vssd1 vccd1 vccd1 _05374_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout180_X net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout278_X net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout657_A net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11665__A1 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09666_ _05302_ _05304_ net732 vssd1 vssd1 vccd1 vccd1 _05305_ sky130_fd_sc_hd__o21a_1
XFILLER_83_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08617_ net1390 _03160_ _03985_ vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__o21a_2
XFILLER_131_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout445_X net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09597_ top.CPU.registers.data\[288\] top.CPU.registers.data\[256\] net810 vssd1
+ vssd1 vccd1 vccd1 _05236_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout824_A net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09997__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08818__C1 top.CPU.control_unit.instruction\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08548_ net605 _04185_ _04186_ _04184_ vssd1 vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__o31a_1
XFILLER_23_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_702 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11968__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout612_X net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08294__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_143_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_143_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_51_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08479_ net938 _04095_ _04096_ net954 vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__o211a_1
XANTENNA__08833__A2 net1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10510_ _04093_ _04158_ net373 vssd1 vssd1 vccd1 vccd1 _06134_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_42_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10640__A2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11490_ _06620_ net258 net255 net3165 vssd1 vssd1 vccd1 vccd1 _02034_ sky130_fd_sc_hd__a22o_1
XFILLER_168_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10441_ _03683_ _03958_ net375 vssd1 vssd1 vccd1 vccd1 _06068_ sky130_fd_sc_hd__mux2_1
XANTENNA__08046__B1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09243__C1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13160_ net1411 top.I2C.bit_timer_state\[0\] _07414_ _07416_ vssd1 vssd1 vccd1 vccd1
+ _02749_ sky130_fd_sc_hd__and4b_1
X_10372_ net548 _03923_ _05712_ _05982_ _05996_ vssd1 vssd1 vccd1 vccd1 _06002_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout981_X net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12111_ net3991 net655 _06823_ vssd1 vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__o21a_1
XFILLER_152_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13091_ top.CPU.data_out\[26\] net2723 net560 vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__mux2_1
XFILLER_108_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12042_ top.CPU.registers.data\[135\] net657 net477 _06592_ net364 vssd1 vssd1 vccd1
+ vccd1 _06793_ sky130_fd_sc_hd__o2111a_1
XANTENNA__07546__A top.CPU.control_unit.instruction\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12145__A2 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold290 top.SPI.parameters\[23\] vssd1 vssd1 vccd1 vccd1 net2847 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10243__Y _05878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11353__B1 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14090__260 clknet_leaf_146_clk vssd1 vssd1 vccd1 vccd1 net1729 sky130_fd_sc_hd__inv_2
XFILLER_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_88_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14387__557 clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 net2026 sky130_fd_sc_hd__inv_2
X_15801_ net2135 _02011_ net1224 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[601\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout770 net771 vssd1 vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__clkbuf_4
Xfanout781 net782 vssd1 vssd1 vccd1 vccd1 net781 sky130_fd_sc_hd__buf_2
Xfanout792 net793 vssd1 vssd1 vccd1 vccd1 net792 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11105__B1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09849__A1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11218__D net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15732_ net2066 _01942_ net1081 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[532\]
+ sky130_fd_sc_hd__dfrtp_1
X_12944_ top.CPU.alu.program_counter\[30\] _03409_ vssd1 vssd1 vccd1 vccd1 _07384_
+ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_66_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14428__598 clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 net2067 sky130_fd_sc_hd__inv_2
X_15663_ net1997 _01873_ net1096 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[463\]
+ sky130_fd_sc_hd__dfrtp_1
X_12875_ top.CPU.alu.program_counter\[23\] _07313_ vssd1 vssd1 vccd1 vccd1 _07322_
+ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_83_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11826_ _06660_ net500 net157 net3383 vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__a22o_1
X_15594_ net1928 _01804_ net1088 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[394\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11234__C _06523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11959__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12081__A1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11757_ net148 net3427 net194 vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_134_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_134_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_147_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10708_ _06278_ _06322_ net306 vssd1 vssd1 vccd1 vccd1 _06323_ sky130_fd_sc_hd__mux2_1
XFILLER_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11688_ net459 _06512_ net235 net165 net3250 vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__a32o_1
X_16215_ net2549 _02425_ net1182 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[1015\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload105 clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 clkload105/Y sky130_fd_sc_hd__clkinv_8
X_13427_ top.CPU.handler.toreg\[1\] _02852_ net120 vssd1 vssd1 vccd1 vccd1 _02467_
+ sky130_fd_sc_hd__mux2_1
X_10639_ _04603_ _06235_ vssd1 vssd1 vccd1 vccd1 _06257_ sky130_fd_sc_hd__or2_1
XANTENNA__09234__C1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload116 clknet_leaf_162_clk vssd1 vssd1 vccd1 vccd1 clkload116/Y sky130_fd_sc_hd__inv_6
Xclkload127 clknet_leaf_169_clk vssd1 vssd1 vccd1 vccd1 clkload127/Y sky130_fd_sc_hd__inv_12
XFILLER_155_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload138 clknet_leaf_146_clk vssd1 vssd1 vccd1 vccd1 clkload138/Y sky130_fd_sc_hd__clkinv_8
XFILLER_127_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14867__1037 clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 net2506 sky130_fd_sc_hd__inv_2
X_16146_ net2480 _02356_ net1104 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[946\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload149 clknet_leaf_130_clk vssd1 vssd1 vccd1 vccd1 clkload149/Y sky130_fd_sc_hd__clkinv_8
X_13358_ net1396 _02887_ net668 vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__mux2_1
XFILLER_128_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07796__C1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12309_ net2612 _03370_ net1246 vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_114_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16077_ net2411 _02287_ net1069 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[877\]
+ sky130_fd_sc_hd__dfrtp_1
X_13289_ _02831_ vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__inv_2
XFILLER_142_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13995__165 clknet_leaf_149_clk vssd1 vssd1 vccd1 vccd1 net1634 sky130_fd_sc_hd__inv_2
X_14331__501 clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 net1970 sky130_fd_sc_hd__inv_2
XANTENNA__09537__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12136__A2 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15028_ clknet_leaf_98_clk _01273_ net1256 vssd1 vssd1 vccd1 vccd1 top.SPI.parameters\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10147__A1 _03476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11344__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07850_ top.CPU.registers.data\[669\] net1289 net1009 top.CPU.registers.data\[701\]
+ net906 vssd1 vssd1 vccd1 vccd1 _03489_ sky130_fd_sc_hd__a221o_1
X_07781_ top.CPU.registers.data\[830\] net1025 net621 _03419_ vssd1 vssd1 vccd1 vccd1
+ _03420_ sky130_fd_sc_hd__a211o_1
Xinput3 DAT_I[10] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
X_09520_ top.CPU.alu.program_counter\[1\] net879 vssd1 vssd1 vccd1 vccd1 _05159_ sky130_fd_sc_hd__nand2_1
XFILLER_65_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08512__A1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16277__Q top.CPU.handler.toreg\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09451_ _05085_ _05088_ net454 vssd1 vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__mux2_1
XANTENNA__07720__C1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08402_ net625 _04036_ _04037_ _04040_ vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__a31o_1
XFILLER_24_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09382_ net1402 net1048 _04953_ _05020_ vssd1 vssd1 vccd1 vccd1 _05021_ sky130_fd_sc_hd__a22o_2
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08333_ net677 _03970_ _03971_ vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_125_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_125_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout140_A _06126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout238_A net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08264_ net941 _03890_ _03891_ net957 vssd1 vssd1 vccd1 vccd1 _03903_ sky130_fd_sc_hd__o211a_1
XFILLER_20_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09225__C1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08195_ top.CPU.registers.data\[567\] top.CPU.registers.data\[535\] net986 vssd1
+ vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1147_A net1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13572__A1 _03009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09240__A2 net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11583__B1 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08674__S1 net1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_754 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1314_A net1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12127__A2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14074__244 clknet_leaf_163_clk vssd1 vssd1 vccd1 vccd1 net1713 sky130_fd_sc_hd__inv_2
XFILLER_114_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10504__B net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11335__B1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout774_A net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1009 net1013 vssd1 vssd1 vccd1 vccd1 net1009 sky130_fd_sc_hd__buf_2
XANTENNA__08200__B1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11319__C _05694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07653__X _03292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08751__A1 _03342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14115__285 clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 net1754 sky130_fd_sc_hd__inv_2
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout562_X net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout941_A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07979_ top.CPU.registers.data\[88\] net1290 net1010 top.CPU.registers.data\[120\]
+ net933 vssd1 vssd1 vccd1 vccd1 _03618_ sky130_fd_sc_hd__a221o_1
XFILLER_74_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13307__S net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09718_ net946 _05333_ _05334_ net960 vssd1 vssd1 vccd1 vccd1 _05357_ sky130_fd_sc_hd__o211a_1
X_10990_ net3648 net216 _06548_ net312 vssd1 vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__a22o_1
XANTENNA__09700__B1 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09649_ _04470_ _04603_ _05283_ _05287_ vssd1 vssd1 vccd1 vccd1 _05288_ sky130_fd_sc_hd__o31a_1
XANTENNA__07532__C net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout827_X net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12660_ _07123_ _07127_ vssd1 vssd1 vccd1 vccd1 _07128_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_26_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08484__X _04123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09059__A2 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ _06149_ net3329 net213 vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__mux2_1
XANTENNA__08267__B1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12591_ _07091_ _07092_ vssd1 vssd1 vccd1 vccd1 _00074_ sky130_fd_sc_hd__nand2_1
XFILLER_24_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09464__C1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_116_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_116_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13042__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10893__C net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14772__942 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 net2411 sky130_fd_sc_hd__inv_2
X_11542_ net3776 net250 _06738_ net480 vssd1 vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__a22o_1
XANTENNA__11810__A1 net1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13012__B1 _07431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11473_ net551 _03181_ net462 _06603_ vssd1 vssd1 vccd1 vccd1 _06728_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_98_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16000_ net2334 _02210_ net1092 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[800\]
+ sky130_fd_sc_hd__dfrtp_1
X_13212_ top.I2C.within_byte_counter_reading\[2\] top.I2C.within_byte_counter_reading\[1\]
+ top.I2C.within_byte_counter_reading\[0\] vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__or3b_2
XANTENNA__13563__A1 top.CPU.addressnew\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10424_ net416 _06051_ _06050_ _06046_ vssd1 vssd1 vccd1 vccd1 _06052_ sky130_fd_sc_hd__o211a_1
X_14813__983 clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 net2452 sky130_fd_sc_hd__inv_2
X_13979__149 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 net1618 sky130_fd_sc_hd__inv_2
XANTENNA__10377__A1 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13143_ top.SPI.command\[5\] top.CPU.data_out\[5\] net557 vssd1 vssd1 vccd1 vccd1
+ _01294_ sky130_fd_sc_hd__mux2_1
XANTENNA__12497__A2_N _05190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10355_ _03857_ net504 _05742_ _05979_ _05985_ vssd1 vssd1 vccd1 vccd1 _05986_ sky130_fd_sc_hd__o221a_1
XANTENNA__13315__A1 _02855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13074_ top.CPU.data_out\[9\] net2713 net560 vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__mux2_1
X_10286_ _05776_ _05779_ net387 vssd1 vssd1 vccd1 vccd1 _05919_ sky130_fd_sc_hd__mux2_1
X_12025_ net3907 net151 _06789_ _06723_ vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__a22o_1
XFILLER_120_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09491__A net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10430__A net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09298__A2 net1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15715_ net2049 _01925_ net1206 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[515\]
+ sky130_fd_sc_hd__dfrtp_1
X_12927_ _07368_ vssd1 vssd1 vccd1 vccd1 _07369_ sky130_fd_sc_hd__inv_2
XFILLER_18_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15646_ net1980 _01856_ net1238 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[446\]
+ sky130_fd_sc_hd__dfrtp_1
X_12858_ top.CPU.alu.program_counter\[21\] _07306_ net1359 vssd1 vssd1 vccd1 vccd1
+ _01184_ sky130_fd_sc_hd__mux2_1
XFILLER_61_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11809_ _06057_ net3822 net156 vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__mux2_1
XANTENNA__10576__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_107_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_107_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09455__C1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15577_ net1911 _01787_ net1223 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[377\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_155_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12357__A net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12789_ top.CPU.alu.program_counter\[15\] _04256_ vssd1 vssd1 vccd1 vccd1 _07244_
+ sky130_fd_sc_hd__nor2_1
XFILLER_159_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_1_Left_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11261__A net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10604__A2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11801__A1 net1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09470__A2 net1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09207__C1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13554__A1 _03100_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09758__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14058__228 clknet_leaf_148_clk vssd1 vssd1 vccd1 vccd1 net1697 sky130_fd_sc_hd__inv_2
XANTENNA__11565__B1 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16129_ net2463 _02339_ net1232 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[929\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_116_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12109__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07784__A2 net1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08951_ top.CPU.registers.data\[874\] top.CPU.registers.data\[842\] net971 vssd1
+ vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__mux2_1
XFILLER_103_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07617__C _03154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11317__B1 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07902_ top.CPU.registers.data_out_r1_prev\[28\] net876 _03525_ _03540_ vssd1 vssd1
+ vccd1 vccd1 _03541_ sky130_fd_sc_hd__o211ai_4
X_08882_ top.CPU.registers.data\[843\] net1309 net840 top.CPU.registers.data\[875\]
+ net761 vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_4_4_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08194__C1 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07833_ net693 _03470_ _03471_ vssd1 vssd1 vccd1 vccd1 _03472_ sky130_fd_sc_hd__or3_1
XANTENNA__13609__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11436__A net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10978__C net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout188_A net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12031__S net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07764_ net801 _03394_ _03395_ net755 vssd1 vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__o211a_1
XANTENNA__09289__A2 net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09503_ top.CPU.registers.data\[961\] net1305 net1028 top.CPU.registers.data\[993\]
+ net921 vssd1 vssd1 vccd1 vccd1 _05142_ sky130_fd_sc_hd__a221o_1
XANTENNA__13490__A0 top.CPU.data_out\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07695_ net1409 _03154_ net1278 net1290 _03104_ vssd1 vssd1 vccd1 vccd1 _03334_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout355_A net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1097_A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09434_ top.CPU.registers.data\[450\] net1294 net1015 top.CPU.registers.data\[482\]
+ net911 vssd1 vssd1 vccd1 vccd1 _05073_ sky130_fd_sc_hd__a221o_1
XFILLER_80_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10994__B _06213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14756__926 clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 net2395 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_23_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10486__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09365_ top.CPU.registers.data\[163\] net1381 net990 top.CPU.registers.data\[131\]
+ net679 vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__a221o_1
XFILLER_12_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout143_X net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout522_A net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11171__A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08316_ top.CPU.registers.data_out_r1_prev\[19\] net875 _03940_ _03954_ vssd1 vssd1
+ vccd1 vccd1 _03955_ sky130_fd_sc_hd__o211ai_4
X_14500__670 clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 net2139 sky130_fd_sc_hd__inv_2
X_09296_ top.CPU.registers.data\[68\] net1299 net1020 top.CPU.registers.data\[100\]
+ net940 vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__a221o_1
XFILLER_138_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout310_X net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08247_ top.CPU.registers.data_out_r1_prev\[22\] net875 net638 _03872_ vssd1 vssd1
+ vccd1 vccd1 _03886_ sky130_fd_sc_hd__o22a_1
XFILLER_165_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1052_X net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout408_X net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13545__A1 _03370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10359__A1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08178_ _03813_ _03816_ net1308 vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__o21a_1
XANTENNA__09213__A2 net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11556__B1 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12714__B _04728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout989_A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10515__A _05665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1317_X net1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10140_ net394 _05775_ vssd1 vssd1 vccd1 vccd1 _05777_ sky130_fd_sc_hd__nand2_1
XFILLER_161_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11308__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout777_X net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10071_ _05055_ net372 vssd1 vssd1 vccd1 vccd1 _05709_ sky130_fd_sc_hd__nor2_1
XFILLER_43_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout944_X net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13037__S net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15473__RESET_B net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07932__C1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13830_ _03130_ _03046_ _03045_ vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__o21bai_1
XANTENNA__07543__B net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13761_ top.wm.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1 _03092_ sky130_fd_sc_hd__and2_1
XFILLER_46_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08488__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13481__B1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14866__1036 clknet_leaf_201_clk vssd1 vssd1 vccd1 vccd1 net2505 sky130_fd_sc_hd__inv_2
X_10973_ net517 _06035_ net546 vssd1 vssd1 vccd1 vccd1 _06538_ sky130_fd_sc_hd__and3_1
XANTENNA__09685__C1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15500_ net1834 _01710_ net1079 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[300\]
+ sky130_fd_sc_hd__dfrtp_1
X_12712_ top.CPU.alu.program_counter\[8\] _07164_ vssd1 vssd1 vccd1 vccd1 _07174_
+ sky130_fd_sc_hd__nor2_1
X_16480_ clknet_leaf_89_clk _02642_ net1273 vssd1 vssd1 vccd1 vccd1 top.SPI.timem\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13692_ net1354 top.SPI.state\[4\] top.SPI.timem\[0\] vssd1 vssd1 vccd1 vccd1 _03050_
+ sky130_fd_sc_hd__a21o_1
X_15431_ net1765 _01641_ net1199 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[231\]
+ sky130_fd_sc_hd__dfrtp_1
X_14499__669 clknet_leaf_170_clk vssd1 vssd1 vccd1 vccd1 net2138 sky130_fd_sc_hd__inv_2
X_12643_ top.I2C.byte_manager_done net4023 vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__and2_1
XANTENNA__09437__C1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11081__A net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15362_ net1696 _01572_ net1171 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[162\]
+ sky130_fd_sc_hd__dfrtp_1
X_12574_ _06008_ _06031_ _06054_ _07078_ vssd1 vssd1 vccd1 vccd1 _07079_ sky130_fd_sc_hd__and4bb_1
XFILLER_50_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11525_ net484 _06057_ net355 net251 net2891 vssd1 vssd1 vccd1 vccd1 _02006_ sky130_fd_sc_hd__a32o_1
XANTENNA__08660__B1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15293_ net1627 _01503_ net1113 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[93\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12905__A top.CPU.alu.program_counter\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_150_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11456_ net3547 net264 net259 _06587_ vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__a22o_1
XANTENNA__08390__A net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09204__A2 net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11547__B1 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08412__A0 _04048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10407_ net574 net517 _06035_ vssd1 vssd1 vccd1 vccd1 _06036_ sky130_fd_sc_hd__and3_1
XANTENNA__11011__A2 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11387_ _06506_ net275 net271 net3231 vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_111_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07766__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13126_ top.SPI.command\[3\] top.SPI.command\[2\] top.SPI.command\[4\] vssd1 vssd1
+ vccd1 vccd1 _02729_ sky130_fd_sc_hd__a21boi_1
XFILLER_140_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10338_ _03859_ _05968_ vssd1 vssd1 vccd1 vccd1 _05969_ sky130_fd_sc_hd__xor2_1
XANTENNA__10770__A1 _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13057_ top.SPI.parameters\[30\] top.SPI.paroutput\[22\] net1355 vssd1 vssd1 vccd1
+ vccd1 _07454_ sky130_fd_sc_hd__mux2_1
X_10269_ _05503_ _05598_ vssd1 vssd1 vccd1 vccd1 _05903_ sky130_fd_sc_hd__or2_1
XANTENNA__08176__C1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1340 net1342 vssd1 vssd1 vccd1 vccd1 net1340 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09425__S net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07734__A net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12008_ _06577_ net350 net151 net3332 vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__a22o_1
Xfanout1351 net1352 vssd1 vssd1 vccd1 vccd1 net1351 sky130_fd_sc_hd__clkbuf_2
Xfanout1362 top.CPU.counter_on vssd1 vssd1 vccd1 vccd1 net1362 sky130_fd_sc_hd__buf_2
XFILLER_39_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1373 net1377 vssd1 vssd1 vccd1 vccd1 net1373 sky130_fd_sc_hd__buf_2
XANTENNA__08810__S1 net1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1384 net1385 vssd1 vssd1 vccd1 vccd1 net1384 sky130_fd_sc_hd__buf_4
XANTENNA__11256__A net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1395 top.CPU.control_unit.instruction\[15\] vssd1 vssd1 vccd1 vccd1 net1395
+ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_109_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14443__613 clknet_leaf_123_clk vssd1 vssd1 vccd1 vccd1 net2082 sky130_fd_sc_hd__inv_2
XANTENNA__11078__A2 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07480_ top.I2C.output_state\[14\] vssd1 vssd1 vccd1 vccd1 _03120_ sky130_fd_sc_hd__inv_2
XANTENNA__09160__S net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09428__C1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15629_ net1963 _01839_ net1064 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[429\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09150_ net958 _04785_ _04786_ net614 vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_170_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10589__A1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11786__B1 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08101_ top.CPU.registers.data\[437\] top.CPU.registers.data\[405\] net830 vssd1
+ vssd1 vccd1 vccd1 _03740_ sky130_fd_sc_hd__mux2_1
XFILLER_147_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11250__A2 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09081_ net929 _04719_ _04718_ net1367 vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__a211o_1
XANTENNA__08651__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09396__A net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08032_ top.CPU.registers.data\[852\] net1318 net849 top.CPU.registers.data\[884\]
+ net743 vssd1 vssd1 vccd1 vccd1 _03671_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_131_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold801 top.CPU.registers.data\[494\] vssd1 vssd1 vccd1 vccd1 net3358 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16290__Q top.CPU.data_out\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold812 top.CPU.registers.data\[540\] vssd1 vssd1 vccd1 vccd1 net3369 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold823 top.CPU.registers.data\[705\] vssd1 vssd1 vccd1 vccd1 net3380 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold834 top.CPU.registers.data\[797\] vssd1 vssd1 vccd1 vccd1 net3391 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08403__B1 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09600__C1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12026__S net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold845 top.CPU.registers.data\[956\] vssd1 vssd1 vccd1 vccd1 net3402 sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 top.CPU.registers.data\[205\] vssd1 vssd1 vccd1 vccd1 net3413 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10210__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold867 top.CPU.registers.data\[869\] vssd1 vssd1 vccd1 vccd1 net3424 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08954__A1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap586 _02965_ vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__clkbuf_2
Xhold878 top.CPU.registers.data\[897\] vssd1 vssd1 vccd1 vccd1 net3435 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_168_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09983_ _05192_ net377 vssd1 vssd1 vccd1 vccd1 _05622_ sky130_fd_sc_hd__nor2_1
XFILLER_27_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold889 top.CPU.registers.data\[159\] vssd1 vssd1 vccd1 vccd1 net3446 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_168_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10054__B _03180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08934_ top.CPU.registers.data\[42\] top.CPU.registers.data\[10\] net972 vssd1 vssd1
+ vccd1 vccd1 _04573_ sky130_fd_sc_hd__mux2_1
XFILLER_131_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1012_A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08167__C1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10989__B net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08865_ net783 _04502_ _04503_ net713 vssd1 vssd1 vccd1 vccd1 _04504_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout472_A net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11710__B1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07914__C1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07816_ net719 _03452_ _03453_ _03454_ vssd1 vssd1 vccd1 vccd1 _03455_ sky130_fd_sc_hd__a31o_1
X_08796_ top.CPU.registers.data\[332\] net1372 net968 top.CPU.registers.data\[364\]
+ net1280 vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__o221a_1
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14186__356 clknet_leaf_146_clk vssd1 vssd1 vccd1 vccd1 net1825 sky130_fd_sc_hd__inv_2
XANTENNA__12266__A1 _06373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07747_ top.CPU.registers.data\[990\] net1332 net863 top.CPU.registers.data\[1022\]
+ net729 vssd1 vssd1 vccd1 vccd1 _03386_ sky130_fd_sc_hd__a221o_1
XANTENNA__13463__B1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout260_X net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09667__C1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_154_Right_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout737_A net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1381_A net1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout358_X net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10277__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09131__A1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_64_Left_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10816__A2 _06419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07678_ _03305_ net550 vssd1 vssd1 vccd1 vccd1 _03317_ sky130_fd_sc_hd__nor2_1
XFILLER_73_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09417_ net409 _05055_ vssd1 vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__nor2_1
XFILLER_25_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14227__397 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 net1866 sky130_fd_sc_hd__inv_2
XANTENNA_fanout904_A net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout525_X net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09348_ top.CPU.alu.program_counter\[4\] _04986_ net1035 vssd1 vssd1 vccd1 vccd1
+ _04987_ sky130_fd_sc_hd__mux2_2
XANTENNA__09434__A2 net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11777__B1 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11900__Y _06770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09279_ _04909_ _04912_ _04917_ vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__a21o_4
XANTENNA__11241__A2 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13518__A1 top.CPU.data_out\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11310_ net3126 net289 net357 net143 vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_95_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12290_ net3796 _04091_ net1192 vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout894_X net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11529__B1 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10890__D _06471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11241_ net487 net465 _06675_ net295 net2663 vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_73_Left_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10245__A net1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07748__A2 net1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11544__A3 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11172_ net1402 net492 _06647_ net300 net3154 vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__a32o_1
XANTENNA__10752__A1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10123_ net417 net410 vssd1 vssd1 vccd1 vccd1 _05761_ sky130_fd_sc_hd__nor2_1
X_15980_ net2314 _02190_ net1076 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[780\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12460__A net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08158__C1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10899__B _06105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14931_ clknet_leaf_62_clk _01177_ net1160 vssd1 vssd1 vccd1 vccd1 top.CPU.alu.program_counter\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_input33_A DAT_I[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14130__300 clknet_leaf_201_clk vssd1 vssd1 vccd1 vccd1 net1769 sky130_fd_sc_hd__inv_2
X_10054_ net552 _03180_ vssd1 vssd1 vccd1 vccd1 _05693_ sky130_fd_sc_hd__and2_2
XANTENNA__11701__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09370__A1 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08173__A2 net1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13813_ net2836 net334 net327 top.CPU.data_out\[15\] vssd1 vssd1 vccd1 vccd1 _02693_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07920__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13454__A0 top.CPU.handler.toreg\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_82_Left_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_121_Right_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11363__X _06714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16532_ clknet_leaf_86_clk net3143 net1265 vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__dfrtp_1
X_13744_ _03081_ _03082_ vssd1 vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__nor2_1
XFILLER_17_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10956_ net515 _06528_ vssd1 vssd1 vccd1 vccd1 _06529_ sky130_fd_sc_hd__and2_1
XANTENNA__08385__A net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08330__C1 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16463_ clknet_leaf_86_clk _02625_ net1265 vssd1 vssd1 vccd1 vccd1 top.SPI.timem\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_104_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13675_ net3536 net331 net330 top.CPU.addressnew\[8\] vssd1 vssd1 vccd1 vccd1 _02603_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11480__A2 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10887_ net133 net437 vssd1 vssd1 vccd1 vccd1 _06486_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_14_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15414_ net1748 _01624_ net1230 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[214\]
+ sky130_fd_sc_hd__dfrtp_1
X_12626_ top.I2C.output_state\[7\] top.I2C.I2C_state\[3\] net1053 _03128_ net2560
+ vssd1 vssd1 vccd1 vccd1 _00026_ sky130_fd_sc_hd__a32o_1
X_16394_ clknet_leaf_50_clk _00019_ net1134 vssd1 vssd1 vccd1 vccd1 top.I2C.read_byte_done
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_129_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11768__B1 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15345_ net1679 _01555_ net1191 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[145\]
+ sky130_fd_sc_hd__dfrtp_1
X_12557_ _03101_ _07054_ net634 vssd1 vssd1 vccd1 vccd1 _07062_ sky130_fd_sc_hd__or3b_1
XANTENNA__08633__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12635__A top.I2C.output_state\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13509__A1 top.CPU.data_out\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13509__B2 _02974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11508_ net567 net532 vssd1 vssd1 vccd1 vccd1 _06731_ sky130_fd_sc_hd__nand2_4
XPHY_EDGE_ROW_91_Left_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07987__A2 net1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15276_ net1610 _01486_ net1076 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[76\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_145_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12488_ _04566_ _04594_ _04633_ _04658_ vssd1 vssd1 vccd1 vccd1 _06997_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_89_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold108 top.CPU.registers.data\[566\] vssd1 vssd1 vccd1 vccd1 net2665 sky130_fd_sc_hd__dlygate4sd3_1
Xhold119 top.CPU.registers.data\[303\] vssd1 vssd1 vccd1 vccd1 net2676 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11439_ top.CPU.registers.data\[665\] net265 vssd1 vssd1 vccd1 vccd1 _06720_ sky130_fd_sc_hd__and2_1
XANTENNA__10155__A net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08397__C1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11940__B1 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13109_ net2680 _02719_ net897 vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__mux2_1
XFILLER_98_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09155__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11299__A2 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_163_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1170 net1277 vssd1 vssd1 vccd1 vccd1 net1170 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_163_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1181 net1188 vssd1 vssd1 vccd1 vccd1 net1181 sky130_fd_sc_hd__clkbuf_2
X_08650_ net701 _04285_ _04288_ vssd1 vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__or3_1
Xfanout1192 net1205 vssd1 vssd1 vccd1 vccd1 net1192 sky130_fd_sc_hd__buf_2
XFILLER_93_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07601_ _03232_ _03239_ net638 vssd1 vssd1 vccd1 vccd1 _03240_ sky130_fd_sc_hd__o21bai_1
XANTENNA__07911__A2 net1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08581_ net788 _04215_ _04216_ net635 vssd1 vssd1 vccd1 vccd1 _04220_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_124_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10259__B1 _05892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13405__S net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07532_ top.CPU.control_unit.instruction\[7\] net1407 net659 vssd1 vssd1 vccd1 vccd1
+ _03171_ sky130_fd_sc_hd__and3_1
XANTENNA__07470__Y _03110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07463_ net1409 vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__inv_2
XANTENNA__11471__A2 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09202_ net618 _04837_ _04840_ net604 vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__a211o_1
XFILLER_22_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11759__B1 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09133_ top.CPU.registers.data\[231\] top.CPU.registers.data\[199\] net995 vssd1
+ vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__mux2_1
XANTENNA__11223__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout220_A _06469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09821__C1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout318_A net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10431__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07978__A2 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09064_ net1283 _04701_ _04702_ vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__or3_1
X_14571__741 clknet_leaf_164_clk vssd1 vssd1 vccd1 vccd1 net2210 sky130_fd_sc_hd__inv_2
XFILLER_163_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13909__79 clknet_leaf_168_clk vssd1 vssd1 vccd1 vccd1 net1548 sky130_fd_sc_hd__inv_2
X_08015_ top.CPU.registers.data\[52\] top.CPU.registers.data\[20\] net816 vssd1 vssd1
+ vccd1 vccd1 _03654_ sky130_fd_sc_hd__mux2_1
Xhold620 top.CPU.registers.data\[369\] vssd1 vssd1 vccd1 vccd1 net3177 sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 top.CPU.registers.data\[264\] vssd1 vssd1 vccd1 vccd1 net3188 sky130_fd_sc_hd__dlygate4sd3_1
Xhold642 top.CPU.registers.data\[325\] vssd1 vssd1 vccd1 vccd1 net3199 sky130_fd_sc_hd__dlygate4sd3_1
X_14865__1035 clknet_leaf_188_clk vssd1 vssd1 vccd1 vccd1 net2504 sky130_fd_sc_hd__inv_2
XANTENNA__08388__C1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold653 top.CPU.registers.data\[712\] vssd1 vssd1 vccd1 vccd1 net3210 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold664 top.SPI.parameters\[5\] vssd1 vssd1 vccd1 vccd1 net3221 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold675 top.CPU.registers.data\[578\] vssd1 vssd1 vccd1 vccd1 net3232 sky130_fd_sc_hd__dlygate4sd3_1
X_14612__782 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 net2251 sky130_fd_sc_hd__inv_2
Xhold686 top.SPI.parameters\[22\] vssd1 vssd1 vccd1 vccd1 net3243 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11931__B1 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold697 top.CPU.registers.data\[2\] vssd1 vssd1 vccd1 vccd1 net3254 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_34_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout687_A _03332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09966_ _03374_ _03407_ _03441_ _05604_ vssd1 vssd1 vccd1 vccd1 _05605_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout1015_X net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08917_ top.CPU.registers.data\[330\] net1314 net845 top.CPU.registers.data\[362\]
+ net772 vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__a221o_1
X_09897_ _04603_ _05283_ _05532_ _05534_ _05535_ vssd1 vssd1 vccd1 vccd1 _05536_ sky130_fd_sc_hd__a311o_1
XANTENNA__12487__B2 _04531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1320 net114 vssd1 vssd1 vccd1 vccd1 net3877 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_96_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_96_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout475_X net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout854_A _03203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1331 top.I2C.data_out\[9\] vssd1 vssd1 vccd1 vccd1 net3888 sky130_fd_sc_hd__dlygate4sd3_1
X_08848_ top.CPU.registers.data\[75\] net1369 net967 top.CPU.registers.data\[107\]
+ net901 vssd1 vssd1 vccd1 vccd1 _04487_ sky130_fd_sc_hd__o221a_1
Xhold1342 top.CPU.registers.data\[40\] vssd1 vssd1 vccd1 vccd1 net3899 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1353 top.CPU.addressnew\[16\] vssd1 vssd1 vccd1 vccd1 net3910 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1364 top.mmio.mem_data_i\[5\] vssd1 vssd1 vccd1 vccd1 net3921 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1375 top.mmio.mem_data_i\[1\] vssd1 vssd1 vccd1 vccd1 net3932 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07902__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1386 top.SPI.timem\[19\] vssd1 vssd1 vccd1 vccd1 net3943 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12239__A1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1397 top.CPU.registers.data\[450\] vssd1 vssd1 vccd1 vccd1 net3954 sky130_fd_sc_hd__dlygate4sd3_1
X_08779_ top.CPU.registers.data\[300\] top.CPU.registers.data\[268\] net814 vssd1
+ vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout642_X net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1384_X net1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13315__S net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09104__A1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10810_ _05127_ _05550_ vssd1 vssd1 vccd1 vccd1 _06420_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ _06637_ net243 net162 net3550 vssd1 vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08312__C1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11998__B1 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07666__A1 _03262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10741_ net659 _06354_ vssd1 vssd1 vccd1 vccd1 _06355_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout907_X net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10670__B1 _06284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13460_ top.CPU.handler.toreg\[19\] _02951_ net120 vssd1 vssd1 vccd1 vccd1 _02485_
+ sky130_fd_sc_hd__mux2_1
X_10672_ top.CPU.fetch.current_ra\[9\] net1040 net633 top.CPU.handler.toreg\[9\] vssd1
+ vssd1 vccd1 vccd1 _06289_ sky130_fd_sc_hd__a22o_1
X_12411_ top.CPU.addressnew\[3\] top.CPU.addressnew\[2\] top.CPU.addressnew\[5\] top.CPU.addressnew\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06937_ sky130_fd_sc_hd__nand4_1
X_13391_ top.mmio.mem_data_i\[23\] net593 net1345 vssd1 vssd1 vccd1 vccd1 _02911_
+ sky130_fd_sc_hd__a21o_1
XFILLER_139_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_20_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_8
X_15130_ clknet_leaf_53_clk _01340_ net1136 vssd1 vssd1 vccd1 vccd1 top.I2C.sda_out
+ sky130_fd_sc_hd__dfstp_1
X_12342_ net37 top.I2C.output_state\[24\] vssd1 vssd1 vccd1 vccd1 _06892_ sky130_fd_sc_hd__and2b_1
XFILLER_127_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08091__A1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07549__A top.CPU.control_unit.instruction\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_138_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15061_ clknet_leaf_55_clk _00015_ net1134 vssd1 vssd1 vccd1 vccd1 top.I2C.output_state\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12273_ _06887_ vssd1 vssd1 vccd1 vccd1 top.CPU.fetch.nrst sky130_fd_sc_hd__inv_2
XFILLER_153_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08918__A1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10406__C _06033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_12_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11224_ net529 net441 net136 net546 vssd1 vssd1 vccd1 vccd1 _06667_ sky130_fd_sc_hd__and4_1
XANTENNA__11517__A3 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10725__A1 _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12902__B top.CPU.alu.program_counter\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11922__B1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13286__A top.CPU.handler.readout vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07555__Y _03194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09483__B net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11155_ net3670 net303 _06637_ net489 vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__a22o_1
X_13923__93 clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 net1562 sky130_fd_sc_hd__inv_2
XFILLER_110_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10106_ _05743_ vssd1 vssd1 vccd1 vccd1 _05744_ sky130_fd_sc_hd__inv_2
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11086_ net3514 net366 _06597_ net324 vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__a22o_1
X_15963_ net2297 _02173_ net1208 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[763\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13675__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_87_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_49_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10037_ _03309_ _03313_ net547 vssd1 vssd1 vccd1 vccd1 _05676_ sky130_fd_sc_hd__and3_1
X_15894_ net2228 _02104_ net1228 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[694\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_76_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11150__A1 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13427__A0 top.CPU.handler.toreg\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11093__X _06604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_86_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11988_ _06550_ net350 net181 net2728 vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__a22o_1
XANTENNA__08303__C1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11989__B1 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13727_ top.SPI.timem\[13\] _03071_ vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__nor2_1
X_16515_ clknet_leaf_49_clk _02677_ net1129 vssd1 vssd1 vccd1 vccd1 top.mmio.mem_data_i\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11253__B _06213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10939_ net3827 net222 _06516_ net316 vssd1 vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__a22o_1
XFILLER_56_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10661__A0 _04567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16446_ clknet_leaf_85_clk _02609_ net1263 vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__dfrtp_1
X_13658_ net2710 _07391_ net663 vssd1 vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12609_ top.SPI.timem\[9\] top.SPI.timem\[8\] top.SPI.timem\[11\] top.SPI.timem\[10\]
+ vssd1 vssd1 vccd1 vccd1 _07109_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_30_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14555__725 clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 net2194 sky130_fd_sc_hd__inv_2
X_16377_ clknet_leaf_73_clk _02586_ net1152 vssd1 vssd1 vccd1 vccd1 top.CPU.fetch.current_ra\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_13589_ net3910 _03019_ net580 vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__mux2_1
XANTENNA__09803__C1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_11_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_8
X_15328_ net1662 _01538_ net1093 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[128\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11756__A3 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10964__B2 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15259_ net1593 _01469_ net1216 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12166__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07893__S net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15505__RESET_B net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09031__B1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10716__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12812__B _04123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11913__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout407 _05023_ vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__buf_2
X_09820_ top.CPU.registers.data\[250\] net1394 net838 top.CPU.registers.data\[218\]
+ net733 vssd1 vssd1 vccd1 vccd1 _05459_ sky130_fd_sc_hd__a221o_1
XFILLER_99_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_165_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout418 _02938_ vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10613__A net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout429 _06642_ vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__buf_4
XFILLER_140_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_129_Left_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09751_ top.CPU.registers.data\[987\] net1328 net862 top.CPU.registers.data\[1019\]
+ net775 vssd1 vssd1 vccd1 vccd1 _05390_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_126_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_78_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_clk sky130_fd_sc_hd__clkbuf_8
X_08702_ net738 _04333_ _04334_ net762 vssd1 vssd1 vccd1 vccd1 _04341_ sky130_fd_sc_hd__o211a_1
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09682_ net710 _05317_ _05318_ net642 vssd1 vssd1 vccd1 vccd1 _05321_ sky130_fd_sc_hd__a31o_1
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08633_ net744 _04270_ _04271_ net694 vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__a31o_1
XANTENNA__07896__A1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout170_A net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11444__A net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout268_A net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08564_ top.CPU.registers.data\[655\] net1314 net845 top.CPU.registers.data\[687\]
+ net716 vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__a221o_1
XANTENNA__09098__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07515_ top.CPU.control_unit.instruction\[6\] net1409 vssd1 vssd1 vccd1 vccd1 _03154_
+ sky130_fd_sc_hd__nand2b_2
XFILLER_120_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09193__S0 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08495_ net793 _04128_ _04129_ net721 vssd1 vssd1 vccd1 vccd1 _04134_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout435_A _06467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_138_Left_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1177_A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout602_A net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout223_X net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14298__468 clknet_leaf_161_clk vssd1 vssd1 vccd1 vccd1 net1937 sky130_fd_sc_hd__inv_2
XFILLER_148_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09116_ top.CPU.registers.data\[551\] top.CPU.registers.data\[519\] net832 vssd1
+ vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__mux2_1
XFILLER_136_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09047_ top.CPU.registers.data\[40\] top.CPU.registers.data\[8\] net808 vssd1 vssd1
+ vccd1 vccd1 _04686_ sky130_fd_sc_hd__mux2_1
XFILLER_164_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15246__RESET_B net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold450 top.CPU.registers.data\[608\] vssd1 vssd1 vccd1 vccd1 net3007 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout592_X net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout971_A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold461 top.CPU.registers.data\[567\] vssd1 vssd1 vccd1 vccd1 net3018 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11904__B1 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold472 top.CPU.registers.data\[216\] vssd1 vssd1 vccd1 vccd1 net3029 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_147_Left_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09573__A1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold483 top.CPU.registers.data\[465\] vssd1 vssd1 vccd1 vccd1 net3040 sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 _01212_ vssd1 vssd1 vccd1 vccd1 net3051 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08781__C1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout930 net935 vssd1 vssd1 vccd1 vccd1 net930 sky130_fd_sc_hd__clkbuf_4
Xfanout941 net942 vssd1 vssd1 vccd1 vccd1 net941 sky130_fd_sc_hd__clkbuf_2
X_09949_ _03959_ _03987_ _05587_ vssd1 vssd1 vccd1 vccd1 _05588_ sky130_fd_sc_hd__o21a_1
Xfanout952 net953 vssd1 vssd1 vccd1 vccd1 net952 sky130_fd_sc_hd__clkbuf_4
Xfanout963 _03337_ vssd1 vssd1 vccd1 vccd1 net963 sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_69_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout857_X net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09325__A1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout974 net975 vssd1 vssd1 vccd1 vccd1 net974 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout985 net1003 vssd1 vssd1 vccd1 vccd1 net985 sky130_fd_sc_hd__clkbuf_4
X_12960_ top.CPU.alu.program_counter\[31\] _07389_ vssd1 vssd1 vccd1 vccd1 _07399_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_5_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout996 net997 vssd1 vssd1 vccd1 vccd1 net996 sky130_fd_sc_hd__clkbuf_4
Xhold1150 top.CPU.registers.data\[228\] vssd1 vssd1 vccd1 vccd1 net3707 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08533__C1 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1161 top.CPU.registers.data\[233\] vssd1 vssd1 vccd1 vccd1 net3718 sky130_fd_sc_hd__dlygate4sd3_1
X_11911_ net3752 net185 net349 _06036_ vssd1 vssd1 vccd1 vccd1 _01655_ sky130_fd_sc_hd__a22o_1
XANTENNA__13553__B _06426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13409__A0 top.CPU.control_unit.instruction\[27\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold1172 top.CPU.registers.data\[865\] vssd1 vssd1 vccd1 vccd1 net3729 sky130_fd_sc_hd__dlygate4sd3_1
X_12891_ top.CPU.alu.program_counter\[24\] _07322_ top.CPU.alu.program_counter\[25\]
+ vssd1 vssd1 vccd1 vccd1 _07336_ sky130_fd_sc_hd__a21oi_1
Xhold1183 top.CPU.registers.data\[951\] vssd1 vssd1 vccd1 vccd1 net3740 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1194 top.CPU.registers.data\[946\] vssd1 vssd1 vccd1 vccd1 net3751 sky130_fd_sc_hd__dlygate4sd3_1
X_11842_ _06673_ net203 net154 net2908 vssd1 vssd1 vccd1 vccd1 _01719_ sky130_fd_sc_hd__a22o_1
XFILLER_166_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_156_Left_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14242__412 clknet_leaf_143_clk vssd1 vssd1 vccd1 vccd1 net1881 sky130_fd_sc_hd__inv_2
XANTENNA__11073__B _06575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08836__B1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11773_ _06616_ net201 net161 net3421 vssd1 vssd1 vccd1 vccd1 _01782_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_64_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10643__A0 _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14539__709 clknet_leaf_164_clk vssd1 vssd1 vccd1 vccd1 net2178 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_101_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16300_ clknet_leaf_107_clk _02509_ net1248 vssd1 vssd1 vccd1 vccd1 top.CPU.data_out\[11\]
+ sky130_fd_sc_hd__dfrtp_2
X_13512_ _04254_ _02966_ vssd1 vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_64_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09759__A top.CPU.alu.program_counter\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10724_ _04862_ _05559_ _06337_ vssd1 vssd1 vccd1 vccd1 _06338_ sky130_fd_sc_hd__a21bo_1
XFILLER_41_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16231_ clknet_leaf_33_clk _02441_ net1123 vssd1 vssd1 vccd1 vccd1 top.CPU.control_unit.instruction\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_13443_ _02881_ _02937_ _02939_ vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__a21o_1
X_10655_ net3388 net225 net312 _06272_ vssd1 vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__a22o_1
XFILLER_173_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16162_ net2496 _02372_ net1173 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[962\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_139_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13374_ top.I2C.data_out\[18\] net556 _02898_ vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__a21oi_1
Xclkload17 clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 clkload17/Y sky130_fd_sc_hd__clkinv_8
XFILLER_154_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10586_ net550 _04397_ net503 _04395_ _06206_ vssd1 vssd1 vccd1 vccd1 _06207_ sky130_fd_sc_hd__o221a_1
Xclkload28 clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 clkload28/Y sky130_fd_sc_hd__inv_16
XFILLER_166_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload39 clknet_leaf_180_clk vssd1 vssd1 vccd1 vccd1 clkload39/Y sky130_fd_sc_hd__inv_4
XFILLER_86_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15113_ net1495 _01326_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r2_prev\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_12325_ net2590 _04255_ net1156 vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__mux2_1
XFILLER_5_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16093_ net2427 _02303_ net1113 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[893\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12913__A top.CPU.alu.program_counter\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12148__B1 _06749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_165_Left_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15044_ clknet_leaf_93_clk _01289_ net1268 vssd1 vssd1 vccd1 vccd1 top.SPI.command\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07566__X _03205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13287__Y _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09013__B1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12256_ net2902 net143 net431 vssd1 vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__mux2_1
XANTENNA__12699__A1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11207_ net3478 net297 _06659_ net479 vssd1 vssd1 vccd1 vccd1 _02247_ sky130_fd_sc_hd__a22o_1
X_12187_ net3871 net656 _06860_ vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__o21a_1
XANTENNA__11371__A1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11138_ net572 net525 net438 _06271_ vssd1 vssd1 vccd1 vccd1 _06628_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_143_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09316__A1 top.CPU.control_unit.instruction\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13112__A2 net1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15946_ net2280 _02156_ net1084 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[746\]
+ sky130_fd_sc_hd__dfrtp_1
X_11069_ net144 net534 vssd1 vssd1 vccd1 vccd1 _06590_ sky130_fd_sc_hd__and2_1
XFILLER_77_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_160_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11123__A1 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_0_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08838__A net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08524__C1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07878__A1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15877_ net2211 _02087_ net1062 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[677\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11264__A net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09619__A2 net1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14864__1034 clknet_leaf_199_clk vssd1 vssd1 vccd1 vccd1 net2503 sky130_fd_sc_hd__inv_2
XANTENNA__11426__A2 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10634__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08280_ _03889_ _03917_ vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_158_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16429_ clknet_leaf_56_clk _00011_ net1142 vssd1 vssd1 vccd1 vccd1 top.I2C.I2C_state\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14026__196 clknet_leaf_150_clk vssd1 vssd1 vccd1 vccd1 net1665 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_119_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11729__A3 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09252__A0 top.CPU.alu.program_counter\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11430__C _06575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10937__B2 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_wire658_X net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08358__A2 net1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13351__A2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout204 net211 vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__clkbuf_4
Xfanout215 _06752_ vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07566__B1 top.CPU.control_unit.instruction\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout226 net227 vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__clkbuf_8
XFILLER_87_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08763__C1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout237 net243 vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__clkbuf_4
X_09803_ top.CPU.registers.data\[666\] net1335 net867 top.CPU.registers.data\[698\]
+ net710 vssd1 vssd1 vccd1 vccd1 _05442_ sky130_fd_sc_hd__a221o_1
Xfanout248 net249 vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__clkbuf_8
Xfanout259 net262 vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__clkbuf_8
XFILLER_87_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14683__853 clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 net2322 sky130_fd_sc_hd__inv_2
X_07995_ net933 _03632_ _03633_ net953 vssd1 vssd1 vccd1 vccd1 _03634_ sky130_fd_sc_hd__o211a_1
XFILLER_75_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09307__A1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09734_ net797 _05371_ _05372_ net751 vssd1 vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__o211a_1
XFILLER_74_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09665_ top.CPU.registers.data\[537\] net869 net698 _05303_ vssd1 vssd1 vccd1 vccd1
+ _05304_ sky130_fd_sc_hd__o211a_1
XANTENNA__10489__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout552_A _03172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14724__894 clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 net2363 sky130_fd_sc_hd__inv_2
XANTENNA_fanout173_X net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1294_A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08616_ net689 _04254_ _04227_ vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__o21ai_2
XFILLER_83_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08530__A2 net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10873__B1 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09596_ _05227_ _05232_ net452 vssd1 vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_46_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11417__A2 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08547_ net953 _04171_ _04170_ net933 vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_46_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout817_A net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout438_X net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08478_ net678 _04101_ _04102_ vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__and3_1
XANTENNA__12090__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout605_X net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1347_X net1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10440_ _05295_ _06065_ _06066_ _06063_ vssd1 vssd1 vccd1 vccd1 _06067_ sky130_fd_sc_hd__a31o_1
XANTENNA__08046__A1 net1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09243__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08597__A2 net1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10371_ net404 _05739_ vssd1 vssd1 vccd1 vccd1 _06001_ sky130_fd_sc_hd__nor2_1
XFILLER_152_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12110_ _06640_ net244 net179 top.CPU.registers.data\[97\] vssd1 vssd1 vccd1 vccd1
+ _06823_ sky130_fd_sc_hd__a22o_1
XFILLER_124_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09518__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13090_ top.CPU.data_out\[25\] net2830 net561 vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__mux2_1
XFILLER_124_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08422__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12041_ _06591_ _06779_ _06781_ net2834 vssd1 vssd1 vccd1 vccd1 _01546_ sky130_fd_sc_hd__a22o_1
XANTENNA__12145__A3 net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold280 net59 vssd1 vssd1 vccd1 vccd1 net2837 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07546__B net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold291 top.SPI.parameters\[27\] vssd1 vssd1 vccd1 vccd1 net2848 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12879__S net1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout760 _03208_ vssd1 vssd1 vccd1 vccd1 net760 sky130_fd_sc_hd__clkbuf_4
X_15800_ net2134 _02010_ net1148 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[600\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout771 net772 vssd1 vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__buf_2
Xfanout782 _03206_ vssd1 vssd1 vccd1 vccd1 net782 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11105__A1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_184_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout793 net794 vssd1 vssd1 vccd1 vccd1 net793 sky130_fd_sc_hd__clkbuf_4
X_12943_ top.CPU.alu.program_counter\[29\] _07383_ net1361 vssd1 vssd1 vccd1 vccd1
+ _01192_ sky130_fd_sc_hd__mux2_1
X_15731_ net2065 _01941_ net1185 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[531\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11656__A2 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_64_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12874_ _07319_ _07320_ vssd1 vssd1 vccd1 vccd1 _07321_ sky130_fd_sc_hd__xnor2_1
X_15662_ net1996 _01872_ net1104 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[462\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11825_ _06659_ net234 net156 net3199 vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__a22o_1
X_15593_ net1927 _01803_ net1060 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[393\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11408__A2 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_199_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11756_ net147 net538 net500 net194 net3003 vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__a32o_1
XFILLER_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12081__A2 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10092__A1 _03684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10707_ _05625_ _05634_ vssd1 vssd1 vccd1 vccd1 _06322_ sky130_fd_sc_hd__nor2_1
XFILLER_140_1008 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11687_ net519 _06510_ net206 net167 net2752 vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__a32o_1
XANTENNA_clkbuf_leaf_122_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13426_ net3897 _02849_ net122 vssd1 vssd1 vccd1 vccd1 _02466_ sky130_fd_sc_hd__mux2_1
X_16214_ net2548 _02424_ net1221 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[1014\]
+ sky130_fd_sc_hd__dfrtp_1
X_10638_ _04603_ _05280_ vssd1 vssd1 vccd1 vccd1 _06256_ sky130_fd_sc_hd__nand2_1
XANTENNA__09234__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload106 clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 clkload106/Y sky130_fd_sc_hd__clkinv_8
XFILLER_155_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload117 clknet_leaf_167_clk vssd1 vssd1 vccd1 vccd1 clkload117/Y sky130_fd_sc_hd__inv_6
Xclkload128 clknet_leaf_170_clk vssd1 vssd1 vccd1 vccd1 clkload128/Y sky130_fd_sc_hd__inv_2
Xclkload139 clknet_leaf_147_clk vssd1 vssd1 vccd1 vccd1 clkload139/Y sky130_fd_sc_hd__inv_16
XANTENNA__09785__A1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11041__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16145_ net2479 _02355_ net1190 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[945\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13581__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13357_ net888 _02886_ vssd1 vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__and2_1
X_10569_ _06190_ vssd1 vssd1 vccd1 vccd1 _06191_ sky130_fd_sc_hd__inv_2
XFILLER_155_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07796__B1 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07737__A top.CPU.alu.program_counter\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12308_ net2561 _05265_ net1175 vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__mux2_1
X_16076_ net2410 _02286_ net1071 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[876\]
+ sky130_fd_sc_hd__dfrtp_1
X_13288_ top.mmio.mem_data_i\[5\] top.mmio.mem_data_i\[4\] top.mmio.mem_data_i\[6\]
+ top.mmio.mem_data_i\[7\] vssd1 vssd1 vccd1 vccd1 _02831_ sky130_fd_sc_hd__and4b_1
XFILLER_170_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14370__540 clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 net2009 sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_137_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15027_ clknet_leaf_95_clk _01272_ net1260 vssd1 vssd1 vccd1 vccd1 top.SPI.parameters\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11259__A net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14667__837 clknet_leaf_164_clk vssd1 vssd1 vccd1 vccd1 net2306 sky130_fd_sc_hd__inv_2
X_12239_ net3158 net138 net433 vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__mux2_1
XANTENNA__12136__A3 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_17_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08745__C1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09952__A _03889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14411__581 clknet_leaf_122_clk vssd1 vssd1 vccd1 vccd1 net2050 sky130_fd_sc_hd__inv_2
X_07780_ top.CPU.registers.data\[798\] net996 vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__and2_1
X_14708__878 clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 net2347 sky130_fd_sc_hd__inv_2
XFILLER_77_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput4 DAT_I[11] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07472__A top.CPU.control_unit.instruction\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09163__S net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11647__A2 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15929_ net2263 _02139_ net1245 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[729\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10855__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09450_ _05084_ _05087_ net454 vssd1 vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__mux2_1
XFILLER_64_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08401_ net618 _04038_ _04039_ net610 vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__a31o_1
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09381_ top.CPU.control_unit.instruction\[23\] _04595_ vssd1 vssd1 vccd1 vccd1 _05020_
+ sky130_fd_sc_hd__or2_1
XFILLER_52_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13413__S net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09399__A net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08332_ top.CPU.registers.data\[755\] net1383 net987 top.CPU.registers.data\[723\]
+ net912 vssd1 vssd1 vccd1 vccd1 _03971_ sky130_fd_sc_hd__a221o_1
XANTENNA__08276__A1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12072__A2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16293__Q top.CPU.data_out\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08263_ net957 _03892_ _03901_ net613 vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__a211o_1
XANTENNA__11441__B net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_0_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout133_A _05990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09225__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08194_ top.CPU.registers.data\[599\] net1295 net1014 top.CPU.registers.data\[631\]
+ net936 vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__a221o_1
XANTENNA__08579__A2 net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11868__S net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout300_A _06645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12553__A net1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1042_A _03165_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11169__A net1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1307_A _03113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08736__C1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout290_X net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout767_A net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07978_ top.CPU.registers.data\[152\] net983 _03616_ vssd1 vssd1 vccd1 vccd1 _03617_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__08478__A net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09717_ net682 _05339_ _05340_ vssd1 vssd1 vccd1 vccd1 _05356_ sky130_fd_sc_hd__and3_1
XANTENNA__11638__A2 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout934_A net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1297_X net1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09161__C1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08503__A2 net1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10012__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09648_ _04470_ _05282_ _05285_ _04331_ _05286_ vssd1 vssd1 vccd1 vccd1 _05287_ sky130_fd_sc_hd__o221a_1
XFILLER_71_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09579_ top.CPU.registers.data\[352\] top.CPU.registers.data\[320\] net976 vssd1
+ vssd1 vccd1 vccd1 _05218_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout722_X net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12728__A top.CPU.alu.program_counter\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13323__S net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11610_ net140 net3453 net214 vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__mux2_1
XFILLER_169_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ net3841 top.wm.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1 _07092_ sky130_fd_sc_hd__o21ai_1
XFILLER_70_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12063__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11541_ _06373_ net354 vssd1 vssd1 vccd1 vccd1 _06738_ sky130_fd_sc_hd__and2_1
XFILLER_168_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10248__A net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11472_ net130 net3582 net264 vssd1 vssd1 vccd1 vccd1 _02050_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_98_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13211_ net3797 _02779_ _02786_ _02773_ vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__a22o_1
X_10423_ net406 _05827_ _06042_ _05664_ vssd1 vssd1 vccd1 vccd1 _06051_ sky130_fd_sc_hd__a211o_1
XANTENNA__13563__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14354__524 clknet_leaf_201_clk vssd1 vssd1 vccd1 vccd1 net1993 sky130_fd_sc_hd__inv_2
X_13142_ top.SPI.command\[4\] top.CPU.data_out\[4\] net557 vssd1 vssd1 vccd1 vccd1
+ _01293_ sky130_fd_sc_hd__mux2_1
XFILLER_109_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10354_ _05640_ _05733_ _05753_ _05650_ vssd1 vssd1 vccd1 vccd1 _05985_ sky130_fd_sc_hd__a22oi_1
XFILLER_152_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13073_ top.CPU.data_out\[8\] net2775 net560 vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__mux2_1
X_14863__1033 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 net2502 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_76_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10285_ net394 _05775_ vssd1 vssd1 vccd1 vccd1 _05918_ sky130_fd_sc_hd__nor2_1
X_12024_ top.CPU.registers.data\[149\] net653 net363 vssd1 vssd1 vccd1 vccd1 _06789_
+ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_168_Right_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10711__A _06141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout590 net591 vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07950__B1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10430__B net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10837__B1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15714_ net2048 _01924_ net1171 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[514\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkload9_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12926_ _07366_ _07367_ vssd1 vssd1 vccd1 vccd1 _07368_ sky130_fd_sc_hd__or2_1
XFILLER_62_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09711__S net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15645_ net1979 _01855_ net1122 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[445\]
+ sky130_fd_sc_hd__dfrtp_1
X_12857_ _07305_ _07304_ net126 vssd1 vssd1 vccd1 vccd1 _07306_ sky130_fd_sc_hd__mux2_1
XFILLER_22_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12638__A top.I2C.output_state\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11808_ _06034_ net3785 net157 vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__mux2_1
X_12788_ top.CPU.alu.program_counter\[14\] _07243_ net1361 vssd1 vssd1 vccd1 vccd1
+ _01177_ sky130_fd_sc_hd__mux2_1
XANTENNA__09455__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08327__S net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15576_ net1910 _01786_ net1101 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[376\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_155_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11262__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13962__132 clknet_leaf_147_clk vssd1 vssd1 vccd1 vccd1 net1601 sky130_fd_sc_hd__inv_2
X_11739_ _06584_ net203 net194 net3089 vssd1 vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__a22o_1
XFILLER_159_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09207__B1 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13554__A2 _03137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13409_ top.CPU.control_unit.instruction\[27\] _02924_ net670 vssd1 vssd1 vccd1 vccd1
+ _02461_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_133_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07769__B1 net1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14097__267 clknet_leaf_190_clk vssd1 vssd1 vccd1 vccd1 net1736 sky130_fd_sc_hd__inv_2
X_16128_ net2462 _02338_ net1092 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[928\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08430__A1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08981__A2 net1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08950_ top.CPU.registers.data\[810\] top.CPU.registers.data\[778\] net971 vssd1
+ vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__mux2_1
X_16059_ net2393 _02269_ net1208 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[859\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11317__B2 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08718__C1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07901_ _03536_ _03539_ net638 vssd1 vssd1 vccd1 vccd1 _03540_ sky130_fd_sc_hd__a21o_1
XFILLER_116_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08881_ top.CPU.registers.data\[811\] top.CPU.registers.data\[779\] net806 vssd1
+ vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_135_Right_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08194__B1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_102_Left_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09391__C1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07473__Y _03113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07832_ net791 _03465_ _03466_ net743 vssd1 vssd1 vccd1 vccd1 _03471_ sky130_fd_sc_hd__o211a_1
XFILLER_99_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13884__54 clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 net1523 sky130_fd_sc_hd__inv_2
XANTENNA__09369__S0 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07763_ net800 _03398_ _03399_ net730 vssd1 vssd1 vccd1 vccd1 _03402_ sky130_fd_sc_hd__o211a_1
XANTENNA__09143__C1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09502_ top.CPU.registers.data\[833\] net1305 net1028 top.CPU.registers.data\[865\]
+ net945 vssd1 vssd1 vccd1 vccd1 _05141_ sky130_fd_sc_hd__a221o_1
X_07694_ _03103_ _03153_ net1279 net1380 net1408 vssd1 vssd1 vccd1 vccd1 _03333_ sky130_fd_sc_hd__o2111a_1
XANTENNA__13490__A1 _04951_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09433_ top.CPU.registers.data\[322\] net1294 net1015 top.CPU.registers.data\[354\]
+ net936 vssd1 vssd1 vccd1 vccd1 _05072_ sky130_fd_sc_hd__a221o_1
XANTENNA__15772__RESET_B net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10546__A1_N net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12561__B_N _06210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout250_A _06733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14795__965 clknet_leaf_164_clk vssd1 vssd1 vccd1 vccd1 net2434 sky130_fd_sc_hd__inv_2
XANTENNA__10994__C net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout348_A net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09364_ top.CPU.registers.data\[195\] net990 net956 _05002_ vssd1 vssd1 vccd1 vccd1
+ _05003_ sky130_fd_sc_hd__a211o_1
XANTENNA__13242__A1 _02803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12045__A2 _06779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_111_Left_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08315_ net796 _03946_ _03953_ net643 vssd1 vssd1 vccd1 vccd1 _03954_ sky130_fd_sc_hd__a211o_1
XANTENNA__11171__B _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13793__A2 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09295_ top.CPU.registers.data\[228\] net1381 net992 top.CPU.registers.data\[196\]
+ net918 vssd1 vssd1 vccd1 vccd1 _04934_ sky130_fd_sc_hd__a221o_1
XFILLER_123_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10068__A _04891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout515_A net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14041__211 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 net1680 sky130_fd_sc_hd__inv_2
XFILLER_165_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14338__508 clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 net1977 sky130_fd_sc_hd__inv_2
X_08246_ _03882_ _03884_ net699 vssd1 vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__mux2_1
XFILLER_138_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09749__A1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11598__S net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13379__A _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08177_ net749 _03814_ _03815_ net707 vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__o211a_1
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout303_X net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10359__A2 _05988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11556__A1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12753__B1 _03118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09068__S net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10515__B _05672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout884_A _03095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13666__X _03048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10007__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1212_X net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_120_Left_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08709__C1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11308__B2 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10070_ _04987_ net377 vssd1 vssd1 vccd1 vccd1 _05708_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout672_X net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11859__A2 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08185__B1 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_102_Right_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08724__A2 _04361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07932__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09134__C1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13760_ top.I2C.which_data_address\[2\] _03090_ _03089_ vssd1 vssd1 vccd1 vccd1 _02645_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_46_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10972_ net3694 net218 _06537_ net318 vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__a22o_1
XFILLER_56_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13481__A1 net1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09685__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10295__A1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09531__S net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10295__B2 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12711_ top.CPU.alu.program_counter\[8\] _07164_ vssd1 vssd1 vccd1 vccd1 _07173_
+ sky130_fd_sc_hd__and2_1
XANTENNA__13561__B _06371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11492__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13691_ net1354 top.SPI.state\[4\] top.SPI.timem\[0\] vssd1 vssd1 vccd1 vccd1 _03049_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12458__A _03541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12642_ top.I2C.byte_manager_done net3779 vssd1 vssd1 vccd1 vccd1 _00005_ sky130_fd_sc_hd__and2_1
X_13946__116 clknet_leaf_160_clk vssd1 vssd1 vccd1 vccd1 net1585 sky130_fd_sc_hd__inv_2
X_15430_ net1764 _01640_ net1072 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[230\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12036__A2 _06779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11081__B _06428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15361_ net1695 _01571_ net1231 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[161\]
+ sky130_fd_sc_hd__dfrtp_1
X_12573_ _06171_ _06188_ vssd1 vssd1 vccd1 vccd1 _07078_ sky130_fd_sc_hd__nor2_1
XFILLER_30_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07999__B1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11524_ _06650_ net260 net252 net3414 vssd1 vssd1 vccd1 vccd1 _02007_ sky130_fd_sc_hd__a22o_1
X_15292_ net1626 _01502_ net1195 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[92\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_168_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12905__B _05499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13536__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09486__B _05123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11455_ net562 net480 vssd1 vssd1 vccd1 vccd1 _06726_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_150_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11547__A1 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10406_ net661 net441 _06033_ vssd1 vssd1 vccd1 vccd1 _06035_ sky130_fd_sc_hd__and3_2
XFILLER_152_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11386_ _06505_ net276 net271 net3656 vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__a22o_1
XANTENNA__10755__C1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13125_ top.SPI.command\[4\] _02727_ top.SPI.command\[3\] top.SPI.command\[2\] vssd1
+ vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_111_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10337_ _03919_ _05967_ vssd1 vssd1 vccd1 vccd1 _05968_ sky130_fd_sc_hd__nand2_1
XFILLER_152_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16230__RESET_B net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13056_ net3617 _07453_ net894 vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__mux2_1
X_10268_ net224 _05901_ _05897_ _05893_ vssd1 vssd1 vccd1 vccd1 _05902_ sky130_fd_sc_hd__o211ai_2
XFILLER_97_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08176__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09373__C1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1330 net1331 vssd1 vssd1 vccd1 vccd1 net1330 sky130_fd_sc_hd__buf_2
X_12007_ _06718_ net239 net151 net3446 vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__a22o_1
Xfanout1341 net1342 vssd1 vssd1 vccd1 vccd1 net1341 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07734__B _03371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1352 net1353 vssd1 vssd1 vccd1 vccd1 net1352 sky130_fd_sc_hd__buf_2
X_10199_ _05728_ _05746_ net309 vssd1 vssd1 vccd1 vccd1 _05835_ sky130_fd_sc_hd__mux2_1
Xfanout1363 top.CPU.alu.immediate\[31\] vssd1 vssd1 vccd1 vccd1 net1363 sky130_fd_sc_hd__clkbuf_4
Xfanout1374 net1377 vssd1 vssd1 vccd1 vccd1 net1374 sky130_fd_sc_hd__clkbuf_4
XFILLER_78_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1385 top.CPU.control_unit.instruction\[20\] vssd1 vssd1 vccd1 vccd1 net1385
+ sky130_fd_sc_hd__buf_4
Xfanout1396 net1399 vssd1 vssd1 vccd1 vccd1 net1396 sky130_fd_sc_hd__clkbuf_4
XFILLER_94_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14482__652 clknet_leaf_201_clk vssd1 vssd1 vccd1 vccd1 net2121 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_109_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08479__A1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09676__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14779__949 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 net2418 sky130_fd_sc_hd__inv_2
XFILLER_47_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09441__S net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12909_ _07351_ _07352_ vssd1 vssd1 vccd1 vccd1 _07353_ sky130_fd_sc_hd__nor2_1
XANTENNA__11483__B1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14523__693 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 net2162 sky130_fd_sc_hd__inv_2
X_15628_ net1962 _01838_ net1079 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[428\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_146_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09428__B1 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08057__S net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15559_ net1893 _01769_ net1197 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[359\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_170_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08100__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08100_ top.CPU.registers.data_out_r1_prev\[21\] net875 net696 _03731_ _03738_ vssd1
+ vssd1 vccd1 vccd1 _03739_ sky130_fd_sc_hd__o2111a_1
XANTENNA__11786__A1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09080_ top.CPU.registers.data\[680\] top.CPU.registers.data\[648\] net975 vssd1
+ vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__mux2_1
XFILLER_147_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08031_ top.CPU.registers.data\[980\] net1318 net849 top.CPU.registers.data\[1012\]
+ net719 vssd1 vssd1 vccd1 vccd1 _03670_ sky130_fd_sc_hd__a221o_1
XANTENNA__13199__A top.I2C.output_state\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold802 top.CPU.registers.data\[285\] vssd1 vssd1 vccd1 vccd1 net3359 sky130_fd_sc_hd__dlygate4sd3_1
Xhold813 top.CPU.registers.data\[380\] vssd1 vssd1 vccd1 vccd1 net3370 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold824 top.CPU.registers.data\[829\] vssd1 vssd1 vccd1 vccd1 net3381 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09600__B1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold835 top.CPU.registers.data\[902\] vssd1 vssd1 vccd1 vccd1 net3392 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10746__C1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold846 top.CPU.registers.data\[632\] vssd1 vssd1 vccd1 vccd1 net3403 sky130_fd_sc_hd__dlygate4sd3_1
Xhold857 top.CPU.registers.data\[597\] vssd1 vssd1 vccd1 vccd1 net3414 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09982_ _05619_ _05620_ vssd1 vssd1 vccd1 vccd1 _05621_ sky130_fd_sc_hd__nor2_1
XFILLER_115_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold868 top.CPU.registers.data\[836\] vssd1 vssd1 vccd1 vccd1 net3425 sky130_fd_sc_hd__dlygate4sd3_1
Xhold879 top.CPU.registers.data\[151\] vssd1 vssd1 vccd1 vccd1 net3436 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_168_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09616__S net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08933_ net1284 _04568_ _04571_ net617 vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__a211o_1
XFILLER_88_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08167__B1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13138__S _07418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout298_A _06645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10989__C net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08864_ top.CPU.registers.data\[587\] net1309 net840 top.CPU.registers.data\[619\]
+ net761 vssd1 vssd1 vccd1 vccd1 _04503_ sky130_fd_sc_hd__a221o_1
XANTENNA__10351__A net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1005_A net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07914__B1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07815_ net743 _03448_ _03449_ vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__and3_1
X_08795_ top.CPU.registers.data\[460\] net1372 net977 top.CPU.registers.data\[492\]
+ net1364 vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__o221a_1
XFILLER_84_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout465_A net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11881__S net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07746_ _03383_ _03384_ net712 vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__a21o_1
XANTENNA__13463__A1 net1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08756__A _04363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11474__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07677_ _03271_ _03284_ _03314_ vssd1 vssd1 vccd1 vccd1 _03316_ sky130_fd_sc_hd__or3_2
XANTENNA_fanout632_A _03291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout253_X net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1374_A net1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09416_ top.CPU.alu.program_counter\[3\] _05054_ net1035 vssd1 vssd1 vccd1 vccd1
+ _05055_ sky130_fd_sc_hd__mux2_2
XFILLER_53_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14862__1032 clknet_leaf_164_clk vssd1 vssd1 vccd1 vccd1 net2501 sky130_fd_sc_hd__inv_2
X_09347_ net776 _04965_ _04972_ _04985_ vssd1 vssd1 vccd1 vccd1 _04986_ sky130_fd_sc_hd__a31o_2
XANTENNA_fanout420_X net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout518_X net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11777__A1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09278_ _04915_ _04916_ net624 _04914_ vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__o211a_1
XANTENNA__08642__A1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13518__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08229_ net802 _03862_ _03863_ net731 vssd1 vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_95_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07850__C1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_839 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10526__A net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11240_ net528 net441 net132 net546 vssd1 vssd1 vccd1 vccd1 _06675_ sky130_fd_sc_hd__and4_1
XFILLER_4_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10245__B net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout887_X net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08945__A2 net1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09593__Y _05232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11171_ net662 _05847_ net430 vssd1 vssd1 vccd1 vccd1 _06647_ sky130_fd_sc_hd__and3_1
X_10122_ _05740_ _05757_ _05759_ vssd1 vssd1 vccd1 vccd1 _05760_ sky130_fd_sc_hd__and3_1
XFILLER_161_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12460__B _05428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08158__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10899__C net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10053_ _05688_ net601 _05691_ vssd1 vssd1 vccd1 vccd1 _05692_ sky130_fd_sc_hd__a21o_2
X_14930_ clknet_leaf_60_clk _01176_ net1160 vssd1 vssd1 vccd1 vccd1 top.CPU.alu.program_counter\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08253__S0 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14466__636 clknet_leaf_140_clk vssd1 vssd1 vccd1 vccd1 net2105 sky130_fd_sc_hd__inv_2
XANTENNA_input26_A DAT_I[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09107__C1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13812_ net3354 net333 net326 top.CPU.data_out\[14\] vssd1 vssd1 vccd1 vccd1 _02692_
+ sky130_fd_sc_hd__a22o_1
XFILLER_29_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14210__380 clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 net1849 sky130_fd_sc_hd__inv_2
XFILLER_29_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10268__A1 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09261__S net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14507__677 clknet_leaf_149_clk vssd1 vssd1 vccd1 vccd1 net2146 sky130_fd_sc_hd__inv_2
X_16531_ clknet_leaf_99_clk _02693_ net1257 vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__dfrtp_1
XFILLER_16_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11465__B1 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13743_ top.SPI.timem\[19\] _03080_ vssd1 vssd1 vccd1 vccd1 _03082_ sky130_fd_sc_hd__and2_1
X_10955_ net659 _05697_ _05808_ net544 vssd1 vssd1 vccd1 vccd1 _06528_ sky130_fd_sc_hd__and4_1
XANTENNA__08330__B1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11092__A net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16462_ clknet_leaf_86_clk _02624_ net1265 vssd1 vssd1 vccd1 vccd1 top.SPI.timem\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12009__A2 _06779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13674_ net3606 net331 net330 top.CPU.addressnew\[7\] vssd1 vssd1 vccd1 vccd1 _02602_
+ sky130_fd_sc_hd__a22o_1
X_10886_ net484 net459 _06485_ net220 net2942 vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__a32o_1
XFILLER_19_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15413_ net1747 _01623_ net1215 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[213\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11217__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12625_ top.I2C.which_data_address\[0\] top.I2C.which_data_address\[1\] top.I2C.which_data_address\[2\]
+ vssd1 vssd1 vccd1 vccd1 _07118_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_14_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16393_ clknet_leaf_51_clk _00067_ net1134 vssd1 vssd1 vccd1 vccd1 top.I2C.reader_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__11768__A1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09497__A net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12556_ net2617 top.CPU.busy _07061_ net2558 vssd1 vssd1 vccd1 vccd1 _00023_ sky130_fd_sc_hd__a211o_1
XFILLER_129_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08633__A1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15344_ net1678 _01554_ net1156 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[144\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_129_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11507_ net481 net472 _06641_ net254 net3007 vssd1 vssd1 vccd1 vccd1 _02018_ sky130_fd_sc_hd__a32o_1
XFILLER_156_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12487_ _04566_ _04594_ _04499_ _04531_ vssd1 vssd1 vccd1 vccd1 _06996_ sky130_fd_sc_hd__o2bb2a_1
X_15275_ net1609 _01485_ net1058 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[75\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_172_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold109 top.CPU.addressnew\[30\] vssd1 vssd1 vccd1 vccd1 net2666 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09189__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11438_ net567 net495 _06580_ net265 net3147 vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__a32o_1
XANTENNA__13390__A0 net1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08397__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12193__B2 _06741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11369_ net474 _06477_ net273 net3325 vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__a22o_1
XANTENNA__12651__A top.CPU.done vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13108_ top.SPI.command\[0\] top.SPI.state\[0\] top.SPI.paroutput\[24\] net1358 vssd1
+ vssd1 vccd1 vccd1 _02719_ sky130_fd_sc_hd__a22o_1
XANTENNA__11267__A net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13039_ top.SPI.parameters\[21\] top.SPI.paroutput\[13\] net1356 vssd1 vssd1 vccd1
+ vccd1 _07445_ sky130_fd_sc_hd__mux2_1
XFILLER_21_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1160 net1164 vssd1 vssd1 vccd1 vccd1 net1160 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_128_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_163_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1171 net1179 vssd1 vssd1 vccd1 vccd1 net1171 sky130_fd_sc_hd__clkbuf_4
Xfanout1182 net1188 vssd1 vssd1 vccd1 vccd1 net1182 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_163_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1193 net1196 vssd1 vssd1 vccd1 vccd1 net1193 sky130_fd_sc_hd__clkbuf_4
X_13854__24 clknet_leaf_150_clk vssd1 vssd1 vccd1 vccd1 net1493 sky130_fd_sc_hd__inv_2
XFILLER_54_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07600_ net802 _03234_ _03235_ _03238_ net699 vssd1 vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__o311a_1
X_08580_ net740 _04217_ _04218_ net766 vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__o211a_1
XANTENNA__07480__A top.I2C.output_state\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10259__A1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09113__A2 net1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07531_ top.CPU.control_unit.instruction\[7\] net659 vssd1 vssd1 vccd1 vccd1 _03170_
+ sky130_fd_sc_hd__nand2_8
XFILLER_35_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11456__B1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07462_ top.I2C.bit_timer_state\[0\] vssd1 vssd1 vccd1 vccd1 _03102_ sky130_fd_sc_hd__inv_2
XFILLER_90_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09201_ net930 _04830_ _04831_ net625 vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__o211a_1
XFILLER_22_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09132_ top.CPU.registers.data\[167\] net1382 net995 top.CPU.registers.data\[135\]
+ net683 vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__a221o_1
XFILLER_33_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09063_ top.CPU.registers.data\[456\] net1373 net970 top.CPU.registers.data\[488\]
+ net1364 vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__o221a_1
XFILLER_135_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12037__S net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07832__C1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout213_A _06752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08014_ top.CPU.registers.data\[340\] net1318 net849 top.CPU.registers.data\[372\]
+ net768 vssd1 vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__a221o_1
XFILLER_151_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold610 top.CPU.registers.data\[29\] vssd1 vssd1 vccd1 vccd1 net3167 sky130_fd_sc_hd__dlygate4sd3_1
Xhold621 top.CPU.registers.data\[404\] vssd1 vssd1 vccd1 vccd1 net3178 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10065__B _05266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold632 top.CPU.registers.data\[452\] vssd1 vssd1 vccd1 vccd1 net3189 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11876__S net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold643 top.CPU.handler.toreg\[3\] vssd1 vssd1 vccd1 vccd1 net3200 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09585__C1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold654 top.CPU.registers.data\[152\] vssd1 vssd1 vccd1 vccd1 net3211 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10195__B1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold665 _01211_ vssd1 vssd1 vccd1 vccd1 net3222 sky130_fd_sc_hd__dlygate4sd3_1
Xhold676 top.CPU.registers.data\[631\] vssd1 vssd1 vccd1 vccd1 net3233 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10734__A2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14153__323 clknet_leaf_157_clk vssd1 vssd1 vccd1 vccd1 net1792 sky130_fd_sc_hd__inv_2
XFILLER_143_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07655__A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold687 top.CPU.registers.data\[26\] vssd1 vssd1 vccd1 vccd1 net3244 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_34_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold698 top.CPU.registers.data\[217\] vssd1 vssd1 vccd1 vccd1 net3255 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10352__Y _05983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09965_ _03243_ _03371_ vssd1 vssd1 vccd1 vccd1 _05604_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout582_A net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09337__C1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08916_ top.CPU.registers.data\[298\] top.CPU.registers.data\[266\] net811 vssd1
+ vssd1 vccd1 vccd1 _04555_ sky130_fd_sc_hd__mux2_1
XFILLER_76_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09896_ _04501_ _04532_ vssd1 vssd1 vccd1 vccd1 _05535_ sky130_fd_sc_hd__and2b_1
XFILLER_112_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1310 top.SPI.command\[7\] vssd1 vssd1 vccd1 vccd1 net3867 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1321 top.I2C.data_out\[8\] vssd1 vssd1 vccd1 vccd1 net3878 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10498__B2 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1332 top.CPU.registers.data\[503\] vssd1 vssd1 vccd1 vccd1 net3889 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout370_X net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1343 top.I2C.data_out\[13\] vssd1 vssd1 vccd1 vccd1 net3900 sky130_fd_sc_hd__dlygate4sd3_1
X_08847_ _04484_ _04485_ net927 vssd1 vssd1 vccd1 vccd1 _04486_ sky130_fd_sc_hd__mux2_1
XANTENNA__07899__C1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1354 top.CPU.registers.data\[751\] vssd1 vssd1 vccd1 vccd1 net3911 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08560__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout847_A net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout468_X net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1365 top.mmio.mem_data_i\[20\] vssd1 vssd1 vccd1 vccd1 net3922 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1376 top.CPU.registers.data\[247\] vssd1 vssd1 vccd1 vccd1 net3933 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13436__A1 _03200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08778_ top.CPU.registers.data\[76\] net1311 net842 top.CPU.registers.data\[108\]
+ net763 vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__a221o_1
Xhold1387 top.CPU.registers.data\[86\] vssd1 vssd1 vccd1 vccd1 net3944 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1398 top.CPU.registers.data\[78\] vssd1 vssd1 vccd1 vccd1 net3955 sky130_fd_sc_hd__dlygate4sd3_1
X_07729_ _03364_ _03367_ _03342_ vssd1 vssd1 vccd1 vccd1 _03368_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_0_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout635_X net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08312__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1377_X net1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10740_ net603 _06352_ _06353_ vssd1 vssd1 vccd1 vccd1 _06354_ sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_0_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10671_ _06273_ _06274_ _06287_ vssd1 vssd1 vccd1 vccd1 _06288_ sky130_fd_sc_hd__o21bai_4
XANTENNA_fanout802_X net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12410_ _06935_ vssd1 vssd1 vccd1 vccd1 _06936_ sky130_fd_sc_hd__inv_2
XANTENNA__13331__S net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13390_ net1365 _02910_ net667 vssd1 vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__mux2_1
XANTENNA__08615__A1 _03342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12341_ net1411 top.I2C.bit_timer_state\[0\] vssd1 vssd1 vccd1 vccd1 _06891_ sky130_fd_sc_hd__or2_2
XANTENNA__07549__B net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07823__C1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15060_ clknet_leaf_49_clk _00064_ net1128 vssd1 vssd1 vccd1 vccd1 top.I2C.output_state\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_126_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12272_ net34 net38 vssd1 vssd1 vccd1 vccd1 _06887_ sky130_fd_sc_hd__nand2_8
XFILLER_5_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13372__A0 top.CPU.control_unit.instruction\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11223_ net493 net468 _06666_ net296 net2647 vssd1 vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__a32o_1
XFILLER_141_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12902__C top.CPU.alu.program_counter\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13286__B _03126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11154_ net474 _06636_ vssd1 vssd1 vccd1 vccd1 _06637_ sky130_fd_sc_hd__nor2_1
XFILLER_1_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10105_ _05332_ _05467_ net374 vssd1 vssd1 vccd1 vccd1 _05743_ sky130_fd_sc_hd__mux2_1
XFILLER_110_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09328__C1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11087__A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15962_ net2296 _02172_ net1253 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[762\]
+ sky130_fd_sc_hd__dfrtp_1
X_11085_ net130 net534 vssd1 vssd1 vccd1 vccd1 _06597_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_145_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10036_ net510 _05674_ _03373_ vssd1 vssd1 vccd1 vccd1 _05675_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09343__A2 net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11686__B1 net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15893_ net2227 _02103_ net1216 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[693\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08551__A0 _04188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11150__A2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16386__Q top.SPI.state\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11438__B1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08303__B1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11987_ _06548_ net342 net180 net2803 vssd1 vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__a22o_1
XFILLER_91_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16514_ clknet_leaf_57_clk _02676_ net1144 vssd1 vssd1 vccd1 vccd1 top.mmio.mem_data_i\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_13726_ _03070_ _03071_ vssd1 vssd1 vccd1 vccd1 _02631_ sky130_fd_sc_hd__nor2_1
XFILLER_90_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10938_ net440 _06428_ net437 vssd1 vssd1 vccd1 vccd1 _06516_ sky130_fd_sc_hd__and3_1
XANTENNA__11253__C net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10661__A1 _04634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16445_ clknet_leaf_86_clk _02608_ net1265 vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__dfrtp_1
X_13657_ net2854 _07382_ net665 vssd1 vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__mux2_1
X_10869_ net493 net468 _06474_ net223 net3098 vssd1 vssd1 vccd1 vccd1 _02400_ sky130_fd_sc_hd__a32o_1
XFILLER_158_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14594__764 clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 net2233 sky130_fd_sc_hd__inv_2
XFILLER_13_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12608_ top.SPI.timem\[1\] top.SPI.timem\[0\] top.SPI.timem\[3\] top.SPI.timem\[2\]
+ vssd1 vssd1 vccd1 vccd1 _07108_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_30_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08067__C1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16376_ clknet_leaf_72_clk _02585_ net1158 vssd1 vssd1 vccd1 vccd1 top.CPU.fetch.current_ra\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08335__S net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13588_ top.CPU.alu.program_counter\[16\] _06147_ net1352 vssd1 vssd1 vccd1 vccd1
+ _03019_ sky130_fd_sc_hd__mux2_1
XFILLER_173_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15327_ net1661 _01537_ net1224 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[127\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07814__C1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12539_ _03322_ _03323_ _07047_ vssd1 vssd1 vccd1 vccd1 _07048_ sky130_fd_sc_hd__mux2_1
XFILLER_69_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10964__A2 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15258_ net1592 _01468_ net1255 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[58\]
+ sky130_fd_sc_hd__dfrtp_1
X_14137__307 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 net1776 sky130_fd_sc_hd__inv_2
XANTENNA__09567__C1 net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08909__A2 net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12381__A top.CPU.handler.readout vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15189_ net1526 _01399_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r1_prev\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_165_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07475__A net1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout408 _05023_ vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__buf_2
Xfanout419 _02938_ vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__clkbuf_2
XFILLER_99_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10613__B net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07593__A1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14861__1031 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 net2500 sky130_fd_sc_hd__inv_2
XANTENNA__13764__X _03095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09750_ top.CPU.registers.data\[955\] top.CPU.registers.data\[923\] net827 vssd1
+ vssd1 vccd1 vccd1 _05389_ sky130_fd_sc_hd__mux2_1
XFILLER_100_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09334__A2 net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08701_ top.CPU.registers.data\[973\] net1311 net842 top.CPU.registers.data\[1005\]
+ net714 vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__a221o_1
XANTENNA__09690__A net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11677__B1 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09681_ top.CPU.registers.data\[761\] net1394 net837 top.CPU.registers.data\[729\]
+ net732 vssd1 vssd1 vccd1 vccd1 _05320_ sky130_fd_sc_hd__a221o_1
XFILLER_66_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13416__S net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08632_ top.CPU.registers.data\[974\] net1320 net851 top.CPU.registers.data\[1006\]
+ net769 vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__a221o_1
XANTENNA__12320__S net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16296__Q top.CPU.data_out\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11429__B1 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08563_ top.CPU.registers.data\[559\] top.CPU.registers.data\[527\] net811 vssd1
+ vssd1 vccd1 vccd1 _04202_ sky130_fd_sc_hd__mux2_1
XANTENNA__11444__B net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout163_A _06760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07514_ top.CPU.control_unit.instruction\[6\] net1409 vssd1 vssd1 vccd1 vccd1 _03153_
+ sky130_fd_sc_hd__and2b_2
XFILLER_63_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07648__A2 net1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09193__S1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08494_ top.CPU.registers.data\[464\] net1322 net852 top.CPU.registers.data\[496\]
+ net771 vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__a221o_1
XFILLER_120_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10652__A1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout330_A _03048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout428_A _06701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1072_A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08058__C1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10404__A1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09115_ net707 _04752_ _04753_ _04751_ vssd1 vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__a31o_1
XFILLER_148_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11601__B1 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10076__A _04698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09270__A1 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout216_X net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1337_A net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07937__X _03576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09046_ top.CPU.registers.data\[456\] net1312 net843 top.CPU.registers.data\[488\]
+ net763 vssd1 vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__a221o_1
XFILLER_117_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout797_A net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09558__C1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold440 top.CPU.registers.data\[717\] vssd1 vssd1 vccd1 vccd1 net2997 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold451 top.CPU.registers.data\[345\] vssd1 vssd1 vccd1 vccd1 net3008 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold462 top.CPU.registers.data\[647\] vssd1 vssd1 vccd1 vccd1 net3019 sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 top.CPU.registers.data\[141\] vssd1 vssd1 vccd1 vccd1 net3030 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08230__C1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold484 top.CPU.registers.data\[582\] vssd1 vssd1 vccd1 vccd1 net3041 sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 top.CPU.registers.data\[392\] vssd1 vssd1 vccd1 vccd1 net3052 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout964_A net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07584__A1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout920 net924 vssd1 vssd1 vccd1 vccd1 net920 sky130_fd_sc_hd__clkbuf_4
Xfanout931 net932 vssd1 vssd1 vccd1 vccd1 net931 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11380__A2 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09948_ _05576_ _05583_ _05586_ _05295_ vssd1 vssd1 vccd1 vccd1 _05587_ sky130_fd_sc_hd__o22a_1
Xfanout942 net949 vssd1 vssd1 vccd1 vccd1 net942 sky130_fd_sc_hd__clkbuf_4
Xfanout953 net963 vssd1 vssd1 vccd1 vccd1 net953 sky130_fd_sc_hd__buf_4
Xfanout964 net965 vssd1 vssd1 vccd1 vccd1 net964 sky130_fd_sc_hd__clkbuf_4
Xfanout975 net976 vssd1 vssd1 vccd1 vccd1 net975 sky130_fd_sc_hd__clkbuf_4
Xfanout986 net989 vssd1 vssd1 vccd1 vccd1 net986 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11668__B1 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09879_ net447 vssd1 vssd1 vccd1 vccd1 _05518_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_5_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout752_X net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout997 net1003 vssd1 vssd1 vccd1 vccd1 net997 sky130_fd_sc_hd__buf_2
Xhold1140 top.CPU.registers.data\[901\] vssd1 vssd1 vccd1 vccd1 net3697 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1151 top.SPI.timem\[1\] vssd1 vssd1 vccd1 vccd1 net3708 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1162 top.CPU.registers.data\[410\] vssd1 vssd1 vccd1 vccd1 net3719 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09730__C1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11910_ net3631 net186 net351 _06011_ vssd1 vssd1 vccd1 vccd1 _01656_ sky130_fd_sc_hd__a22o_1
XFILLER_45_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1173 top.CPU.registers.data\[852\] vssd1 vssd1 vccd1 vccd1 net3730 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12890_ top.CPU.alu.program_counter\[24\] _03118_ _07333_ _07335_ vssd1 vssd1 vccd1
+ vccd1 _01187_ sky130_fd_sc_hd__a22o_1
XANTENNA__11683__A3 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1184 top.CPU.registers.data\[856\] vssd1 vssd1 vccd1 vccd1 net3741 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1195 top.CPU.registers.data\[245\] vssd1 vssd1 vccd1 vccd1 net3752 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09105__A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11841_ _06672_ net210 net154 net2708 vssd1 vssd1 vccd1 vccd1 _01720_ sky130_fd_sc_hd__a22o_1
XANTENNA__12093__B1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14281__451 clknet_leaf_157_clk vssd1 vssd1 vccd1 vccd1 net1920 sky130_fd_sc_hd__inv_2
X_11772_ _06615_ net203 net162 net3519 vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_101_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14578__748 clknet_leaf_193_clk vssd1 vssd1 vccd1 vccd1 net2217 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10643__A1 _04567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13511_ top.CPU.data_out\[14\] net588 _02969_ _02975_ vssd1 vssd1 vccd1 vccd1 _02512_
+ sky130_fd_sc_hd__o22a_1
X_10723_ _04862_ _05559_ net511 vssd1 vssd1 vccd1 vccd1 _06337_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_64_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11840__B1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09759__B net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16230_ clknet_leaf_72_clk _02440_ net1152 vssd1 vssd1 vccd1 vccd1 top.CPU.control_unit.instruction\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_81_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13442_ net3798 _02942_ net121 vssd1 vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__mux2_1
X_10654_ net572 net513 net438 _06271_ vssd1 vssd1 vccd1 vccd1 _06272_ sky130_fd_sc_hd__and4_1
XFILLER_174_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_750 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08155__S net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14322__492 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 net1961 sky130_fd_sc_hd__inv_2
X_14619__789 clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 net2258 sky130_fd_sc_hd__inv_2
XFILLER_154_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13373_ net1345 top.mmio.mem_data_i\[18\] net597 vssd1 vssd1 vccd1 vccd1 _02898_
+ sky130_fd_sc_hd__o21a_1
X_16161_ net2495 _02371_ net1224 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[961\]
+ sky130_fd_sc_hd__dfrtp_1
X_10585_ _04392_ net506 net508 _04394_ vssd1 vssd1 vccd1 vccd1 _06206_ sky130_fd_sc_hd__o2bb2a_1
Xclkload18 clknet_leaf_193_clk vssd1 vssd1 vccd1 vccd1 clkload18/Y sky130_fd_sc_hd__inv_4
Xclkload29 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 clkload29/Y sky130_fd_sc_hd__inv_4
X_15112_ net1494 _01325_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r2_prev\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09775__A net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12324_ net2568 _04188_ net1156 vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__mux2_1
X_16092_ net2426 _02302_ net1193 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[892\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12913__B _05429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15043_ clknet_leaf_91_clk _01288_ vssd1 vssd1 vccd1 vccd1 top.SPI.percount\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_12255_ net3166 _06149_ net432 vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__mux2_1
XANTENNA__10159__B1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_147_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11206_ net456 _06374_ net429 vssd1 vssd1 vccd1 vccd1 _06659_ sky130_fd_sc_hd__and3_1
XANTENNA__09564__A2 net1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12186_ net568 net364 _06668_ net170 top.CPU.registers.data\[58\] vssd1 vssd1 vccd1
+ vccd1 _06860_ sky130_fd_sc_hd__a32o_1
XFILLER_122_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11371__A2 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11137_ net478 net456 _06627_ net301 net3575 vssd1 vssd1 vccd1 vccd1 _02285_ sky130_fd_sc_hd__a32o_1
XFILLER_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13648__A1 _07300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11248__C net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11659__B1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11068_ net323 net145 net535 net366 net2688 vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__a32o_1
X_15945_ net2279 _02155_ net1056 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[745\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_160_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11123__A2 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12320__A1 _03716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08524__B1 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10019_ _03613_ _05332_ net374 vssd1 vssd1 vccd1 vccd1 _05658_ sky130_fd_sc_hd__mux2_1
X_15876_ net2210 _02086_ net1198 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[676\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11674__A3 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08288__C1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13709_ top.SPI.timem\[7\] _03058_ vssd1 vssd1 vccd1 vccd1 _03060_ sky130_fd_sc_hd__and2_1
XFILLER_32_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_158_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16428_ clknet_leaf_56_clk _00010_ net1135 vssd1 vssd1 vccd1 vccd1 top.I2C.I2C_state\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13584__A0 top.CPU.alu.program_counter\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16359_ clknet_leaf_32_clk _02568_ net1125 vssd1 vssd1 vccd1 vccd1 top.CPU.fetch.current_ra\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09252__A1 _04889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08055__A2 net1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10937__A2 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08460__C1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07476__Y _03116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11439__B net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout205 net211 vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__buf_4
XANTENNA__11362__A2 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout216 net219 vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08763__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10635__C_N net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout227 net228 vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__clkbuf_8
X_09802_ top.CPU.registers.data\[922\] net1337 net867 top.CPU.registers.data\[954\]
+ net698 vssd1 vssd1 vccd1 vccd1 _05441_ sky130_fd_sc_hd__a221o_1
Xfanout238 net239 vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09691__Y _05330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout249 _06739_ vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__clkbuf_8
XFILLER_87_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07994_ top.CPU.registers.data\[920\] net1290 net1010 top.CPU.registers.data\[952\]
+ net907 vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__a221o_1
XFILLER_140_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09733_ top.CPU.registers.data\[763\] net1391 net827 top.CPU.registers.data\[731\]
+ net777 vssd1 vssd1 vccd1 vccd1 _05372_ sky130_fd_sc_hd__a221o_1
XFILLER_68_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10630__Y _06249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout280_A net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12311__A1 _03508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08515__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout378_A net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11455__A net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09664_ top.CPU.registers.data\[569\] net837 vssd1 vssd1 vccd1 vccd1 _05303_ sky130_fd_sc_hd__or2_1
XANTENNA__12862__A2 _03756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11665__A3 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14265__435 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 net1904 sky130_fd_sc_hd__inv_2
X_08615_ _03342_ _04240_ _04253_ vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__o21ai_4
XANTENNA__11174__B net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10873__A1 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09595_ _05226_ _05233_ net455 vssd1 vssd1 vccd1 vccd1 _05234_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout166_X net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout545_A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1287_A net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08818__A1 net1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08546_ net676 _04168_ _04169_ net909 vssd1 vssd1 vccd1 vccd1 _04185_ sky130_fd_sc_hd__o211a_1
XFILLER_35_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13811__B2 top.CPU.data_out\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14306__476 clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 net1945 sky130_fd_sc_hd__inv_2
XANTENNA__11822__B1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08477_ top.CPU.registers.data_out_r2_prev\[17\] net687 net620 _04115_ vssd1 vssd1
+ vccd1 vccd1 _04116_ sky130_fd_sc_hd__o211a_1
XFILLER_168_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08294__A2 net1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout712_A _03212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13834__4 clknet_leaf_146_clk vssd1 vssd1 vccd1 vccd1 net1473 sky130_fd_sc_hd__inv_2
XANTENNA_fanout1075_X net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11190__A net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13575__B1 _03011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09779__C1 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout500_X net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1242_X net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_149_Right_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10370_ net407 _05999_ vssd1 vssd1 vccd1 vccd1 _06000_ sky130_fd_sc_hd__nor2_1
XANTENNA__11050__B2 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13327__A0 top.CPU.control_unit.instruction\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_156_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09029_ top.CPU.registers.data\[808\] top.CPU.registers.data\[776\] net811 vssd1
+ vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__mux2_1
X_12040_ _06590_ _06779_ _06781_ net3251 vssd1 vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__a22o_1
XANTENNA__11889__A0 _06311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold270 top.CPU.addressnew\[25\] vssd1 vssd1 vccd1 vccd1 net2827 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08203__C1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08754__A0 _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07557__A1 net1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold281 top.CPU.registers.data\[178\] vssd1 vssd1 vccd1 vccd1 net2838 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_160_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11353__A2 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold292 top.CPU.registers.data\[880\] vssd1 vssd1 vccd1 vccd1 net2849 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_160_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout750 net760 vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__clkbuf_2
Xfanout761 net764 vssd1 vssd1 vccd1 vccd1 net761 sky130_fd_sc_hd__clkbuf_4
Xfanout772 net782 vssd1 vssd1 vccd1 vccd1 net772 sky130_fd_sc_hd__buf_2
Xfanout783 net786 vssd1 vssd1 vccd1 vccd1 net783 sky130_fd_sc_hd__buf_2
XANTENNA__12302__A1 _04828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout794 _03205_ vssd1 vssd1 vccd1 vccd1 net794 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11105__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13056__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15730_ net2064 _01940_ net1102 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[530\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09703__C1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12942_ _07382_ _07379_ net129 vssd1 vssd1 vccd1 vccd1 _07383_ sky130_fd_sc_hd__mux2_1
XFILLER_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15661_ net1995 _01871_ net1059 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[461\]
+ sky130_fd_sc_hd__dfrtp_1
X_12873_ top.CPU.alu.program_counter\[22\] _03916_ _07310_ vssd1 vssd1 vccd1 vccd1
+ _07320_ sky130_fd_sc_hd__a21o_1
XFILLER_65_86 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_83_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11824_ _06355_ net3563 net156 vssd1 vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__mux2_1
XANTENNA__12066__B1 _03185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15592_ net1926 _01802_ net1089 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[392\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_159_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13802__B2 top.CPU.data_out\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11755_ _06594_ net197 net192 net2963 vssd1 vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__a22o_1
X_14860__1030 clknet_leaf_189_clk vssd1 vssd1 vccd1 vccd1 net2499 sky130_fd_sc_hd__inv_2
X_10706_ net397 _06243_ vssd1 vssd1 vccd1 vccd1 _06321_ sky130_fd_sc_hd__nand2_1
XANTENNA__10092__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11686_ _06507_ net196 net164 net3152 vssd1 vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__a22o_1
XANTENNA__13566__A0 top.CPU.alu.program_counter\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16213_ net2547 _02423_ net1210 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[1013\]
+ sky130_fd_sc_hd__dfrtp_1
X_13425_ _07062_ _07065_ _07077_ _07080_ vssd1 vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__and4bb_1
XFILLER_174_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10637_ net3680 net225 net311 _06255_ vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__a22o_1
Xclkload107 clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 clkload107/Y sky130_fd_sc_hd__clkinv_8
Xclkload118 clknet_leaf_182_clk vssd1 vssd1 vccd1 vccd1 clkload118/Y sky130_fd_sc_hd__inv_8
XANTENNA__11041__A1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15890__RESET_B net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload129 clknet_leaf_171_clk vssd1 vssd1 vccd1 vccd1 clkload129/Y sky130_fd_sc_hd__inv_2
X_16144_ net2478 _02354_ net1155 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[944\]
+ sky130_fd_sc_hd__dfrtp_1
X_10568_ net602 _06188_ _06189_ vssd1 vssd1 vccd1 vccd1 _06190_ sky130_fd_sc_hd__a21oi_4
X_13356_ top.I2C.data_out\[13\] net553 _02885_ net596 vssd1 vssd1 vccd1 vccd1 _02886_
+ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_116_Right_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08993__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12307_ net3825 _05191_ net1253 vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__mux2_1
XANTENNA__07737__B net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16075_ net2409 _02285_ net1058 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[875\]
+ sky130_fd_sc_hd__dfrtp_1
X_13287_ top.CPU.handler.readout _03126_ vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__nand2_4
X_10499_ _06115_ _06121_ _06123_ vssd1 vssd1 vccd1 vccd1 _06124_ sky130_fd_sc_hd__and3_2
XFILLER_154_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_15_Left_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15026_ clknet_leaf_98_clk _01271_ net1254 vssd1 vssd1 vccd1 vccd1 top.SPI.parameters\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09537__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12238_ _06572_ _06796_ _06885_ net168 net3179 vssd1 vssd1 vccd1 vccd1 _01442_ sky130_fd_sc_hd__a32o_1
XFILLER_96_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11344__A2 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12169_ net4009 net174 _06852_ _06660_ vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__a22o_1
XFILLER_96_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07753__A net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14249__419 clknet_leaf_158_clk vssd1 vssd1 vccd1 vccd1 net1888 sky130_fd_sc_hd__inv_2
Xinput5 DAT_I[12] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11275__A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15928_ net2262 _02138_ net1148 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[728\]
+ sky130_fd_sc_hd__dfrtp_1
X_15859_ net2193 _02069_ net1186 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[659\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07720__A1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08400_ top.CPU.registers.data\[754\] net1379 net978 top.CPU.registers.data\[722\]
+ net909 vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__a221o_1
X_09380_ _05018_ vssd1 vssd1 vccd1 vccd1 _05019_ sky130_fd_sc_hd__inv_2
XANTENNA__12057__B1 _03185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08584__A _04222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08331_ top.CPU.registers.data\[595\] net1294 net1015 top.CPU.registers.data\[627\]
+ net936 vssd1 vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__a221o_1
XFILLER_51_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11804__B1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11214__S net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08262_ net680 _03893_ _03894_ vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_173_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11280__B2 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08193_ top.CPU.registers.data\[759\] net1381 net987 top.CPU.registers.data\[727\]
+ net912 vssd1 vssd1 vccd1 vccd1 _03832_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout126_A net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14650__820 clknet_leaf_162_clk vssd1 vssd1 vccd1 vccd1 net2289 sky130_fd_sc_hd__inv_2
XANTENNA__08523__S net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12553__B top.SPI.busy vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08984__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11583__A2 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1035_A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11335__A2 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11884__S net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout495_A net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08200__A2 net1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout283_X net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07977_ top.CPU.registers.data\[184\] net1010 net907 vssd1 vssd1 vccd1 vccd1 _03616_
+ sky130_fd_sc_hd__a21o_1
XFILLER_68_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09716_ top.CPU.registers.data_out_r2_prev\[25\] net688 _05353_ _05354_ net622 vssd1
+ vssd1 vccd1 vccd1 _05355_ sky130_fd_sc_hd__o221a_1
XANTENNA__11099__B2 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09161__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10846__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09700__A2 net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09647_ _04259_ _04327_ _04258_ vssd1 vssd1 vccd1 vccd1 _05286_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout548_X net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout927_A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13604__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12048__B1 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09578_ top.CPU.registers.data\[288\] top.CPU.registers.data\[256\] net976 vssd1
+ vssd1 vccd1 vccd1 _05217_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13796__B1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08529_ top.CPU.registers.data\[48\] top.CPU.registers.data\[16\] net984 vssd1 vssd1
+ vccd1 vccd1 _04168_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout715_X net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09464__A1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08267__A2 net1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11540_ net483 _06355_ net355 net251 net3041 vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__a32o_1
XANTENNA__08672__C1 net1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11810__A3 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11471_ net567 net494 _06596_ net266 net2733 vssd1 vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__a32o_1
XANTENNA__10816__X _06426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09216__A1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12744__A top.CPU.alu.program_counter\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13012__A2 _07429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13210_ net892 top.I2C.data_out\[21\] _02785_ vssd1 vssd1 vccd1 vccd1 _02786_ sky130_fd_sc_hd__mux2_1
X_10422_ _05817_ _05982_ _06048_ _06049_ vssd1 vssd1 vccd1 vccd1 _06050_ sky130_fd_sc_hd__o211a_1
XANTENNA__09529__S net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12220__B1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14393__563 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 net2032 sky130_fd_sc_hd__inv_2
XFILLER_152_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13141_ top.SPI.command\[3\] top.CPU.data_out\[3\] net557 vssd1 vssd1 vccd1 vccd1
+ _01292_ sky130_fd_sc_hd__mux2_1
X_10353_ _03315_ _03859_ _05632_ _05981_ _05980_ vssd1 vssd1 vccd1 vccd1 _05984_ sky130_fd_sc_hd__a221o_1
XFILLER_3_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10782__B1 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13072_ top.CPU.data_out\[7\] net3064 net558 vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__mux2_1
XFILLER_152_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10284_ _05365_ net510 net505 _05366_ _05916_ vssd1 vssd1 vccd1 vccd1 _05917_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_76_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12023_ net365 _06722_ _06788_ _06787_ vssd1 vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__a31o_1
XFILLER_78_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout580 net582 vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__clkbuf_4
XFILLER_65_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09152__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10430__C net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15713_ net2047 _01923_ net1231 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[513\]
+ sky130_fd_sc_hd__dfrtp_1
X_12925_ top.CPU.alu.program_counter\[28\] _03576_ vssd1 vssd1 vccd1 vccd1 _07367_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__10837__B2 top.CPU.handler.toreg\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12919__A top.CPU.alu.program_counter\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12039__A0 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15644_ net1978 _01854_ net1234 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[444\]
+ sky130_fd_sc_hd__dfrtp_1
X_12856_ top.CPU.alu.program_counter\[21\] _07298_ vssd1 vssd1 vccd1 vccd1 _07305_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__13787__B1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11807_ _06488_ _06643_ net239 net158 net3371 vssd1 vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__a32o_1
XFILLER_92_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15575_ net1909 _01785_ net1180 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[375\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12787_ _07242_ _07239_ net128 vssd1 vssd1 vccd1 vccd1 _07243_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_155_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11262__A1 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11738_ _06583_ net500 net194 net2990 vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__a22o_1
XANTENNA__11801__A3 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14634__804 clknet_leaf_151_clk vssd1 vssd1 vccd1 vccd1 net2273 sky130_fd_sc_hd__inv_2
XFILLER_174_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_116_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11669_ _06484_ net209 net167 net3318 vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_116_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13408_ net890 _02923_ vssd1 vssd1 vccd1 vccd1 _02924_ sky130_fd_sc_hd__and2_1
XANTENNA__09758__A2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11014__B2 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_133_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08966__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11565__A2 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16127_ net2461 _02337_ net1219 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[927\]
+ sky130_fd_sc_hd__dfrtp_1
X_13339_ top.mmio.mem_data_i\[9\] net592 net1343 vssd1 vssd1 vccd1 vccd1 _02873_ sky130_fd_sc_hd__a21o_1
XFILLER_51_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10174__A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10773__B1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16058_ net2392 _02268_ net1243 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[858\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_103_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11317__A2 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13485__A _03137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15009_ clknet_leaf_96_clk _01254_ net1248 vssd1 vssd1 vccd1 vccd1 top.SPI.parameters\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_07900_ net700 _03537_ _03538_ vssd1 vssd1 vccd1 vccd1 _03539_ sky130_fd_sc_hd__or3_1
XFILLER_69_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08880_ net784 _04517_ _04518_ net713 vssd1 vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__o211a_1
XFILLER_116_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09391__B1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07831_ net791 _03459_ _03460_ net719 vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__o211a_1
XANTENNA__14953__RESET_B net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11436__C net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09369__S1 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07762_ net754 _03392_ _03393_ net712 vssd1 vssd1 vccd1 vccd1 _03401_ sky130_fd_sc_hd__a31o_1
XFILLER_38_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07770__X _03409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09501_ top.CPU.registers.data_out_r2_prev\[1\] net688 _05137_ _05139_ net960 vssd1
+ vssd1 vccd1 vccd1 _05140_ sky130_fd_sc_hd__o221a_1
X_07693_ net1047 _03262_ vssd1 vssd1 vccd1 vccd1 _03332_ sky130_fd_sc_hd__nand2_4
XFILLER_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_998 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13424__S net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09432_ top.CPU.registers.data_out_r2_prev\[2\] net687 net620 _05063_ vssd1 vssd1
+ vccd1 vccd1 _05071_ sky130_fd_sc_hd__o211a_1
XFILLER_169_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09363_ top.CPU.registers.data\[227\] net1381 vssd1 vssd1 vccd1 vccd1 _05002_ sky130_fd_sc_hd__and2_1
XFILLER_36_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08314_ _03949_ _03952_ net1308 vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__o21a_1
XANTENNA__12450__B1 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09294_ _04930_ _04931_ _04932_ net918 net957 vssd1 vssd1 vccd1 vccd1 _04933_ sky130_fd_sc_hd__o221a_1
XANTENNA__11171__C net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10068__B net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14080__250 clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 net1719 sky130_fd_sc_hd__inv_2
XFILLER_20_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08245_ net802 _03873_ _03874_ _03883_ vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__a31o_1
XANTENNA__11879__S net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14377__547 clknet_leaf_157_clk vssd1 vssd1 vccd1 vccd1 net2016 sky130_fd_sc_hd__inv_2
XANTENNA_fanout410_A net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1152_A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout129_X net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout508_A net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_183_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08176_ top.CPU.registers.data\[919\] net1325 net856 top.CPU.registers.data\[951\]
+ net724 vssd1 vssd1 vccd1 vccd1 _03815_ sky130_fd_sc_hd__a221o_1
XANTENNA__08406__C1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12753__A1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14121__291 clknet_leaf_155_clk vssd1 vssd1 vccd1 vccd1 net1760 sky130_fd_sc_hd__inv_2
XFILLER_4_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11556__A2 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_63_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14418__588 clknet_leaf_193_clk vssd1 vssd1 vccd1 vccd1 net2057 sky130_fd_sc_hd__inv_2
XFILLER_173_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1038_X net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08709__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11308__A2 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_198_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout498_X net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1205_X net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_78_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout665_X net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_121_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10971_ net520 _06010_ _06523_ vssd1 vssd1 vccd1 vccd1 _06537_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout832_X net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08488__A2 net1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13481__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12710_ top.CPU.alu.program_counter\[7\] _07172_ net1360 vssd1 vssd1 vccd1 vccd1
+ _01170_ sky130_fd_sc_hd__mux2_1
XANTENNA__10295__A2 _05367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13690_ net2636 net337 vssd1 vssd1 vccd1 vccd1 _02618_ sky130_fd_sc_hd__and2_1
XANTENNA__08428__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12458__B _03575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_136_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13985__155 clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 net1624 sky130_fd_sc_hd__inv_2
X_12641_ net2780 top.I2C.read_byte_done vssd1 vssd1 vccd1 vccd1 _00006_ sky130_fd_sc_hd__and2_1
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09437__A1 net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11081__C net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15360_ net1694 _01570_ net1092 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[160\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_16_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12572_ top.CPU.done _06462_ _07075_ _07068_ vssd1 vssd1 vccd1 vccd1 _07077_ sky130_fd_sc_hd__a31o_1
XANTENNA__08645__C1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11523_ net3502 net252 _06734_ _06488_ vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__a22o_1
X_15291_ net1625 _01501_ net1210 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[91\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08660__A2 net1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11454_ net570 _03189_ vssd1 vssd1 vccd1 vccd1 _06725_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_150_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10405_ net661 _06033_ vssd1 vssd1 vccd1 vccd1 _06034_ sky130_fd_sc_hd__and2_1
XFILLER_137_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11385_ _06504_ net275 net271 net3281 vssd1 vssd1 vccd1 vccd1 _02125_ sky130_fd_sc_hd__a22o_1
XANTENNA__09070__C1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10755__B1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13124_ top.SPI.command\[0\] top.SPI.command\[5\] _07093_ vssd1 vssd1 vccd1 vccd1
+ _02727_ sky130_fd_sc_hd__and3b_1
XFILLER_11_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10336_ _04057_ _05966_ _03922_ vssd1 vssd1 vccd1 vccd1 _05967_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_111_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_9_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_9_0_clk sky130_fd_sc_hd__clkbuf_8
X_10267_ _05900_ _05793_ vssd1 vssd1 vccd1 vccd1 _05901_ sky130_fd_sc_hd__and2b_1
X_13055_ top.SPI.parameters\[29\] top.SPI.paroutput\[21\] net1355 vssd1 vssd1 vccd1
+ vccd1 _07453_ sky130_fd_sc_hd__mux2_1
XANTENNA__10507__B1 _05643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1320 net1322 vssd1 vssd1 vccd1 vccd1 net1320 sky130_fd_sc_hd__clkbuf_4
X_12006_ net1401 _06575_ _06751_ vssd1 vssd1 vccd1 vccd1 _06781_ sky130_fd_sc_hd__or3_4
XFILLER_121_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1331 _03109_ vssd1 vssd1 vccd1 vccd1 net1331 sky130_fd_sc_hd__buf_2
Xfanout1342 _03102_ vssd1 vssd1 vccd1 vccd1 net1342 sky130_fd_sc_hd__clkbuf_2
X_10198_ net384 _05743_ net395 vssd1 vssd1 vccd1 vccd1 _05834_ sky130_fd_sc_hd__a21oi_1
Xfanout1353 top.CPU.handler.state\[3\] vssd1 vssd1 vccd1 vccd1 net1353 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11180__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1364 net1365 vssd1 vssd1 vccd1 vccd1 net1364 sky130_fd_sc_hd__buf_4
XFILLER_93_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1375 net1376 vssd1 vssd1 vccd1 vccd1 net1375 sky130_fd_sc_hd__buf_2
XANTENNA__08686__X _04325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1386 net1388 vssd1 vssd1 vccd1 vccd1 net1386 sky130_fd_sc_hd__clkbuf_4
Xfanout1397 net1399 vssd1 vssd1 vccd1 vccd1 net1397 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09676__A1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12908_ _07340_ _07342_ _07350_ _07339_ vssd1 vssd1 vccd1 vccd1 _07352_ sky130_fd_sc_hd__a211oi_1
XANTENNA__12680__B1 _03118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09023__A net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10691__C1 _06301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15627_ net1961 _01837_ net1064 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[427\]
+ sky130_fd_sc_hd__dfrtp_1
X_12839_ _07289_ _07286_ net127 vssd1 vssd1 vccd1 vccd1 _07290_ sky130_fd_sc_hd__mux2_1
X_14064__234 clknet_leaf_194_clk vssd1 vssd1 vccd1 vccd1 net1703 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_174_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11235__B2 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15558_ net1892 _01768_ net1073 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[358\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_170_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12384__A _06918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15489_ net1823 _01699_ net1232 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[289\]
+ sky130_fd_sc_hd__dfrtp_1
X_14105__275 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 net1744 sky130_fd_sc_hd__inv_2
X_08030_ net693 _03667_ _03668_ vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__and3_1
XANTENNA__07478__A net1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput30 DAT_I[6] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08939__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold803 top.CPU.registers.data\[261\] vssd1 vssd1 vccd1 vccd1 net3360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold814 top.CPU.registers.data\[342\] vssd1 vssd1 vccd1 vccd1 net3371 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08403__A2 net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold825 top.CPU.registers.data\[198\] vssd1 vssd1 vccd1 vccd1 net3382 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold836 top.CPU.registers.data\[39\] vssd1 vssd1 vccd1 vccd1 net3393 sky130_fd_sc_hd__dlygate4sd3_1
Xhold847 top.CPU.registers.data\[649\] vssd1 vssd1 vccd1 vccd1 net3404 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold858 top.CPU.registers.data\[365\] vssd1 vssd1 vccd1 vccd1 net3415 sky130_fd_sc_hd__dlygate4sd3_1
X_09981_ _05123_ net372 vssd1 vssd1 vccd1 vccd1 _05620_ sky130_fd_sc_hd__nor2_1
Xhold869 top.CPU.registers.data\[845\] vssd1 vssd1 vccd1 vccd1 net3426 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08801__S net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_168_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08932_ _04569_ _04570_ net1367 vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__o21a_1
XANTENNA__11728__A net1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12323__S net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09364__B1 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16299__Q top.CPU.data_out\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10989__D net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14762__932 clknet_leaf_145_clk vssd1 vssd1 vccd1 vccd1 net2401 sky130_fd_sc_hd__inv_2
X_08863_ top.CPU.registers.data\[555\] top.CPU.registers.data\[523\] net806 vssd1
+ vssd1 vccd1 vccd1 _04502_ sky130_fd_sc_hd__mux2_1
XFILLER_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout193_A net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11710__A2 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07814_ top.CPU.registers.data\[861\] net1318 net850 top.CPU.registers.data\[893\]
+ net693 vssd1 vssd1 vccd1 vccd1 _03453_ sky130_fd_sc_hd__a221o_1
X_08794_ top.CPU.registers.data\[428\] top.CPU.registers.data\[396\] top.CPU.registers.data\[300\]
+ top.CPU.registers.data\[268\] net977 net1280 vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__mux4_1
XFILLER_38_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07745_ top.CPU.registers.data\[766\] net1394 net833 top.CPU.registers.data\[734\]
+ net730 vssd1 vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout360_A net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14803__973 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 net2442 sky130_fd_sc_hd__inv_2
XFILLER_72_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12559__A _05806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13463__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13969__139 clknet_leaf_190_clk vssd1 vssd1 vccd1 vccd1 net1608 sky130_fd_sc_hd__inv_2
XANTENNA_fanout458_A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07676_ _03298_ _03310_ _03313_ vssd1 vssd1 vccd1 vccd1 _03315_ sky130_fd_sc_hd__and3_4
XANTENNA__12278__B _06887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09415_ top.CPU.registers.data_out_r1_prev\[3\] net875 _05039_ _05053_ vssd1 vssd1
+ vccd1 vccd1 _05054_ sky130_fd_sc_hd__o211a_2
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout246_X net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout625_A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1367_A net1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09346_ net798 _04978_ _04984_ vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__and3_1
XANTENNA__08627__C1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout413_X net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09277_ net672 _04898_ _04899_ net611 vssd1 vssd1 vccd1 vccd1 _04916_ sky130_fd_sc_hd__a31o_1
XFILLER_166_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08228_ top.CPU.registers.data\[470\] net1330 net861 top.CPU.registers.data\[502\]
+ net776 vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_95_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07850__B1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout994_A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10526__B net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11529__A2 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10018__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08159_ net795 _03792_ _03793_ net723 vssd1 vssd1 vccd1 vccd1 _03798_ sky130_fd_sc_hd__o211a_1
XFILLER_10_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09052__C1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1322_X net1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10245__C net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09807__S net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07602__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11170_ net3800 net297 _06646_ net484 vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__a22o_1
XFILLER_164_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout782_X net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10121_ net396 net385 net417 vssd1 vssd1 vccd1 vccd1 _05759_ sky130_fd_sc_hd__o21ai_2
XFILLER_122_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10542__A net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10052_ top.CPU.fetch.current_ra\[31\] net1043 net634 top.CPU.handler.toreg\[31\]
+ vssd1 vssd1 vccd1 vccd1 _05691_ sky130_fd_sc_hd__a22o_1
XANTENNA__09108__A net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07905__A1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11162__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08253__S1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11701__A2 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08947__A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13811_ net3692 net333 net326 top.CPU.data_out\[13\] vssd1 vssd1 vccd1 vccd1 _02691_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_input19_A DAT_I[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12469__A _03754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16530_ clknet_leaf_99_clk _02692_ net1255 vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__dfrtp_1
X_13742_ net3943 _03080_ vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__nor2_1
X_14048__218 clknet_leaf_110_clk vssd1 vssd1 vccd1 vccd1 net1687 sky130_fd_sc_hd__inv_2
XANTENNA__11465__A1 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10954_ net3491 net218 _06527_ net321 vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__a22o_1
XFILLER_73_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16461_ clknet_leaf_87_clk _02623_ net1272 vssd1 vssd1 vccd1 vccd1 top.SPI.timem\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13673_ net3313 net332 net330 top.CPU.addressnew\[6\] vssd1 vssd1 vccd1 vccd1 _02601_
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_191_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_191_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10885_ _05961_ net436 vssd1 vssd1 vccd1 vccd1 _06485_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_104_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11217__A1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15412_ net1746 _01622_ net1113 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[212\]
+ sky130_fd_sc_hd__dfrtp_1
X_12624_ _03125_ top.I2C.I2C_state\[2\] net3657 vssd1 vssd1 vccd1 vccd1 _00032_ sky130_fd_sc_hd__a21o_1
XANTENNA__09778__A net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16392_ clknet_leaf_86_clk _00020_ net1264 vssd1 vssd1 vccd1 vccd1 top.SPI.register\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_157_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15343_ net1677 _01553_ net1099 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[143\]
+ sky130_fd_sc_hd__dfrtp_1
X_12555_ top.CPU.done _07060_ vssd1 vssd1 vccd1 vccd1 _07061_ sky130_fd_sc_hd__nor2_1
XFILLER_106_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11506_ _06640_ net261 net257 net3647 vssd1 vssd1 vccd1 vccd1 _02019_ sky130_fd_sc_hd__a22o_1
XFILLER_129_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15274_ net1608 _01484_ net1088 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[74\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07841__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12486_ _06974_ _06975_ _06994_ _06972_ vssd1 vssd1 vccd1 vccd1 _06995_ sky130_fd_sc_hd__o211a_1
XFILLER_8_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09269__S0 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11437_ net3422 net265 _06719_ net489 vssd1 vssd1 vccd1 vccd1 _02077_ sky130_fd_sc_hd__a22o_1
XFILLER_7_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12193__A2 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11368_ _06476_ net283 net274 net3135 vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__a22o_1
XFILLER_98_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16451__RESET_B net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13107_ _03140_ top.SPI.count\[2\] _02716_ _02718_ vssd1 vssd1 vccd1 vccd1 _01277_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__14920__Q top.CPU.alu.program_counter\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14746__916 clknet_leaf_158_clk vssd1 vssd1 vccd1 vccd1 net2385 sky130_fd_sc_hd__inv_2
XFILLER_3_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11940__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10319_ _03650_ _05594_ net512 vssd1 vssd1 vccd1 vccd1 _05951_ sky130_fd_sc_hd__o21a_1
XFILLER_112_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11299_ net3588 net291 _06707_ net494 vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__a22o_1
XANTENNA__13142__A1 top.CPU.data_out\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13038_ net3967 _07444_ net894 vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__mux2_1
XFILLER_26_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09018__A _03331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1150 net1151 vssd1 vssd1 vccd1 vccd1 net1150 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_128_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1161 net1164 vssd1 vssd1 vccd1 vccd1 net1161 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_128_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1172 net1179 vssd1 vssd1 vccd1 vccd1 net1172 sky130_fd_sc_hd__clkbuf_2
XFILLER_66_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_163_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1183 net1188 vssd1 vssd1 vccd1 vccd1 net1183 sky130_fd_sc_hd__clkbuf_2
XFILLER_67_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10900__B1 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1194 net1196 vssd1 vssd1 vccd1 vccd1 net1194 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09452__S net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14989_ clknet_leaf_90_clk _01234_ net1267 vssd1 vssd1 vccd1 vccd1 top.SPI.paroutput\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_81_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11283__A net1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07530_ top.CPU.control_unit.instruction\[7\] net662 vssd1 vssd1 vccd1 vccd1 _03169_
+ sky130_fd_sc_hd__and2_2
XANTENNA__08857__C1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07461_ top.CPU.handler.state\[5\] vssd1 vssd1 vccd1 vccd1 _03101_ sky130_fd_sc_hd__inv_2
XANTENNA__10664__C1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_182_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_182_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_90_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09200_ net625 _04832_ _04838_ net610 vssd1 vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__a211o_1
XFILLER_50_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08609__C1 net1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11759__A2 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09131_ net958 _04769_ _04768_ net614 vssd1 vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__a211o_1
XFILLER_120_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09062_ top.CPU.registers.data\[328\] net1376 net970 top.CPU.registers.data\[360\]
+ net1281 vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__o221a_1
XFILLER_148_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10431__A2 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Left_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08013_ top.CPU.registers.data\[308\] top.CPU.registers.data\[276\] net816 vssd1
+ vssd1 vccd1 vccd1 _03652_ sky130_fd_sc_hd__mux2_1
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09034__C1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold600 top.CPU.registers.data\[785\] vssd1 vssd1 vccd1 vccd1 net3157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold611 top.CPU.registers.data\[983\] vssd1 vssd1 vccd1 vccd1 net3168 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout206_A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold622 top.CPU.registers.data\[32\] vssd1 vssd1 vccd1 vccd1 net3179 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08388__A1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold633 top.CPU.registers.data\[719\] vssd1 vssd1 vccd1 vccd1 net3190 sky130_fd_sc_hd__dlygate4sd3_1
Xhold644 top.CPU.registers.data\[700\] vssd1 vssd1 vccd1 vccd1 net3201 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold655 top.I2C.I2C_state\[25\] vssd1 vssd1 vccd1 vccd1 net3212 sky130_fd_sc_hd__dlygate4sd3_1
X_14192__362 clknet_leaf_197_clk vssd1 vssd1 vccd1 vccd1 net1831 sky130_fd_sc_hd__inv_2
XANTENNA__11392__B1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold666 top.CPU.registers.data\[932\] vssd1 vssd1 vccd1 vccd1 net3223 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07596__C1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold677 top.I2C.output_state\[9\] vssd1 vssd1 vccd1 vccd1 net3234 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11931__A2 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold688 top.CPU.registers.data\[278\] vssd1 vssd1 vccd1 vccd1 net3245 sky130_fd_sc_hd__dlygate4sd3_1
X_09964_ _05601_ _05594_ _05367_ _03650_ vssd1 vssd1 vccd1 vccd1 _05603_ sky130_fd_sc_hd__nand4b_2
Xhold699 top.CPU.registers.data\[130\] vssd1 vssd1 vccd1 vccd1 net3256 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_34_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14489__659 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 net2128 sky130_fd_sc_hd__inv_2
XANTENNA__09337__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08915_ net787 _04552_ _04553_ net741 vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_51_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09895_ _05283_ _05533_ vssd1 vssd1 vccd1 vccd1 _05534_ sky130_fd_sc_hd__and2_1
XANTENNA__11144__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11892__S net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout196_X net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1300 top.CPU.registers.data\[230\] vssd1 vssd1 vccd1 vccd1 net3857 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1311 top.CPU.fetch.current_ra\[8\] vssd1 vssd1 vccd1 vccd1 net3868 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1322 top.I2C.data_out\[2\] vssd1 vssd1 vccd1 vccd1 net3879 sky130_fd_sc_hd__dlygate4sd3_1
X_08846_ top.CPU.registers.data\[171\] top.CPU.registers.data\[139\] net969 vssd1
+ vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__mux2_1
Xhold1333 top.CPU.registers.data\[954\] vssd1 vssd1 vccd1 vccd1 net3890 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1344 top.CPU.registers.data\[282\] vssd1 vssd1 vccd1 vccd1 net3901 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07671__A _03291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1355 top.CPU.registers.data\[103\] vssd1 vssd1 vccd1 vccd1 net3912 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1366 top.I2C.I2C_state\[8\] vssd1 vssd1 vccd1 vccd1 net3923 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1377 top.CPU.registers.data\[77\] vssd1 vssd1 vccd1 vccd1 net3934 sky130_fd_sc_hd__dlygate4sd3_1
X_08777_ top.CPU.registers.data\[44\] top.CPU.registers.data\[12\] net815 vssd1 vssd1
+ vccd1 vccd1 _04416_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout742_A net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout363_X net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1388 top.CPU.registers.data\[92\] vssd1 vssd1 vccd1 vccd1 net3945 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1399 top.CPU.registers.data\[107\] vssd1 vssd1 vccd1 vccd1 net3956 sky130_fd_sc_hd__dlygate4sd3_1
X_07728_ net923 _03366_ _03365_ net628 vssd1 vssd1 vccd1 vccd1 _03367_ sky130_fd_sc_hd__o211a_1
XANTENNA__11447__B2 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08848__C1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11998__A2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07659_ net1044 _03252_ _03292_ _03296_ vssd1 vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__or4bb_2
XFILLER_14_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_173_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_173_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout530_X net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout628_X net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10670_ _06285_ _06286_ _06284_ vssd1 vssd1 vccd1 vccd1 _06287_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09499__S0 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09329_ net752 _04966_ _04967_ net696 vssd1 vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__o211a_1
XANTENNA__08076__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09273__C1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12340_ net2631 _05226_ net1096 vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__mux2_1
XFILLER_126_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout997_X net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12271_ net3027 net131 net431 vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__mux2_1
X_14433__603 clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 net2072 sky130_fd_sc_hd__inv_2
XANTENNA__12752__A net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08379__A1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12175__A2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11222_ net532 net442 _05848_ net545 vssd1 vssd1 vccd1 vccd1 _06666_ sky130_fd_sc_hd__and4_1
XANTENNA__11383__B1 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12471__B _04048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13059__S net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11922__A2 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12902__D _07322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11153_ net552 net517 net502 net149 vssd1 vssd1 vccd1 vccd1 _06636_ sky130_fd_sc_hd__or4b_1
XFILLER_1_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09328__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10104_ net411 _05665_ vssd1 vssd1 vccd1 vccd1 _05742_ sky130_fd_sc_hd__nand2_2
XFILLER_122_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11087__B _03185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11084_ net3435 net369 _06596_ net319 vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__a22o_1
X_15961_ net2295 _02171_ net1245 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[761\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09423__S0 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10035_ _05673_ vssd1 vssd1 vccd1 vccd1 _05674_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_145_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12883__B1 _03916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15892_ net2226 _02102_ net1082 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[692\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08551__A1 _04189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11438__A1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_86_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11986_ _06547_ net345 net181 net3002 vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_86_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16513_ clknet_leaf_47_clk _02675_ net1137 vssd1 vssd1 vccd1 vccd1 top.mmio.mem_data_i\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11989__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09500__B1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13725_ top.SPI.timem\[12\] _07109_ _03060_ vssd1 vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__and3_1
XFILLER_17_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10937_ net3714 net222 _06515_ net317 vssd1 vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_164_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_164_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_56_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11831__A net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16444_ clknet_leaf_81_clk _02607_ net1242 vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__dfrtp_1
XFILLER_143_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13656_ net3129 _07365_ net665 vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__mux2_1
X_10868_ net137 _06467_ vssd1 vssd1 vccd1 vccd1 _06474_ sky130_fd_sc_hd__and2_1
XANTENNA__10718__Y _06333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12607_ top.SPI.timem\[5\] top.SPI.timem\[4\] top.SPI.timem\[6\] top.SPI.timem\[7\]
+ vssd1 vssd1 vccd1 vccd1 _07107_ sky130_fd_sc_hd__or4b_1
X_16375_ clknet_leaf_73_clk _02584_ net1158 vssd1 vssd1 vccd1 vccd1 top.CPU.fetch.current_ra\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13587_ net3949 _03018_ net580 vssd1 vssd1 vccd1 vccd1 _02545_ sky130_fd_sc_hd__mux2_1
XFILLER_13_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10799_ net444 _06408_ _06409_ _06401_ vssd1 vssd1 vccd1 vccd1 _06410_ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_30_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15326_ net1660 _01536_ net1201 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[126\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_173_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12538_ _05580_ _07046_ vssd1 vssd1 vccd1 vccd1 _07047_ sky130_fd_sc_hd__or2_1
XANTENNA__07814__B1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09016__C1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15257_ net1591 _01467_ net1245 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[57\]
+ sky130_fd_sc_hd__dfrtp_1
X_12469_ _03754_ _03783_ vssd1 vssd1 vccd1 vccd1 _06978_ sky130_fd_sc_hd__nand2_1
X_14176__346 clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 net1815 sky130_fd_sc_hd__inv_2
XANTENNA__12166__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15188_ net1525 _01398_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r1_prev\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12381__B _03126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09031__A2 net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11374__B1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11913__A2 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_165_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout409 _05023_ vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_165_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09319__A0 _04952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13914__84 clknet_leaf_159_clk vssd1 vssd1 vccd1 vccd1 net1553 sky130_fd_sc_hd__inv_2
XFILLER_113_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14217__387 clknet_leaf_157_clk vssd1 vssd1 vccd1 vccd1 net1856 sky130_fd_sc_hd__inv_2
XANTENNA__10613__C net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13666__A2 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08858__Y _04497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08700_ top.CPU.registers.data\[845\] net1311 net842 top.CPU.registers.data\[877\]
+ net738 vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__a221o_1
XANTENNA__11677__A1 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09680_ top.CPU.registers.data\[601\] net1336 net869 top.CPU.registers.data\[633\]
+ net757 vssd1 vssd1 vccd1 vccd1 _05319_ sky130_fd_sc_hd__a221o_1
XANTENNA__10910__A _05694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08631_ net792 _04269_ vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__or2_1
XFILLER_39_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08562_ net788 _04195_ _04196_ _04200_ net636 vssd1 vssd1 vccd1 vccd1 _04201_ sky130_fd_sc_hd__a311o_1
XANTENNA__09098__A2 net1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11444__C _05694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07513_ _03149_ _03105_ _03145_ vssd1 vssd1 vccd1 vccd1 _03152_ sky130_fd_sc_hd__and3b_2
XFILLER_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_155_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_155_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_63_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08493_ top.CPU.registers.data\[432\] top.CPU.registers.data\[400\] net821 vssd1
+ vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout156_A net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13004__Y _07431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08058__B1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09255__C1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout323_A net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09114_ top.CPU.registers.data\[967\] net1326 net857 top.CPU.registers.data\[999\]
+ net724 vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__a221o_1
XFILLER_148_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10076__B net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11887__S net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09045_ net785 _04683_ vssd1 vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__or2_1
XFILLER_164_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1232_A net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout209_X net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12157__A2 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09558__B1 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold430 top.CPU.registers.data\[937\] vssd1 vssd1 vccd1 vccd1 net2987 sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 top.CPU.registers.data\[636\] vssd1 vssd1 vccd1 vccd1 net2998 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold452 top.CPU.registers.data\[416\] vssd1 vssd1 vccd1 vccd1 net3009 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout692_A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold463 top.CPU.registers.data\[517\] vssd1 vssd1 vccd1 vccd1 net3020 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11188__A net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11904__A2 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold474 top.CPU.registers.data\[477\] vssd1 vssd1 vccd1 vccd1 net3031 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1020_X net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold485 top.CPU.registers.data\[423\] vssd1 vssd1 vccd1 vccd1 net3042 sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 top.I2C.output_state\[18\] vssd1 vssd1 vccd1 vccd1 net3053 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08781__A1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout910 _03353_ vssd1 vssd1 vccd1 vccd1 net910 sky130_fd_sc_hd__buf_2
Xfanout921 net922 vssd1 vssd1 vccd1 vccd1 net921 sky130_fd_sc_hd__clkbuf_4
X_09947_ _05297_ _05584_ _05585_ vssd1 vssd1 vccd1 vccd1 _05586_ sky130_fd_sc_hd__a21boi_1
Xfanout932 net935 vssd1 vssd1 vccd1 vccd1 net932 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout480_X net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout943 net944 vssd1 vssd1 vccd1 vccd1 net943 sky130_fd_sc_hd__clkbuf_4
Xfanout954 net962 vssd1 vssd1 vccd1 vccd1 net954 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout578_X net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout957_A net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout965 net966 vssd1 vssd1 vccd1 vccd1 net965 sky130_fd_sc_hd__clkbuf_4
Xfanout976 net1003 vssd1 vssd1 vccd1 vccd1 net976 sky130_fd_sc_hd__buf_2
XFILLER_58_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09878_ _03273_ _03312_ _03325_ _05516_ vssd1 vssd1 vccd1 vccd1 _05517_ sky130_fd_sc_hd__or4_1
XANTENNA__10820__A net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout987 net989 vssd1 vssd1 vccd1 vccd1 net987 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout998 net1002 vssd1 vssd1 vccd1 vccd1 net998 sky130_fd_sc_hd__clkbuf_4
Xhold1130 top.CPU.registers.data\[761\] vssd1 vssd1 vccd1 vccd1 net3687 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08497__A net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1141 top.I2C.I2C_state\[9\] vssd1 vssd1 vccd1 vccd1 net3698 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08533__A1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09730__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1152 top.SPI.timem\[6\] vssd1 vssd1 vccd1 vccd1 net3709 sky130_fd_sc_hd__dlygate4sd3_1
X_08829_ _04466_ _04467_ vssd1 vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__nor2_1
Xhold1163 top.CPU.registers.data\[955\] vssd1 vssd1 vccd1 vccd1 net3720 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1174 top.CPU.registers.data\[67\] vssd1 vssd1 vccd1 vccd1 net3731 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout745_X net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1185 top.CPU.registers.data\[866\] vssd1 vssd1 vccd1 vccd1 net3742 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07741__C1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1196 top.CPU.registers.data\[239\] vssd1 vssd1 vccd1 vccd1 net3753 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11840_ _06671_ net238 net154 net3125 vssd1 vssd1 vccd1 vccd1 _01721_ sky130_fd_sc_hd__a22o_1
XFILLER_166_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_146_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_146_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout912_X net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11771_ _06614_ net210 net162 net3705 vssd1 vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__a22o_1
XANTENNA__09494__C1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13510_ _04323_ _02966_ vssd1 vssd1 vccd1 vccd1 _02975_ sky130_fd_sc_hd__nor2_2
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10722_ net3644 net227 net316 _06336_ vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_64_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13441_ _02878_ _02937_ _02939_ vssd1 vssd1 vccd1 vccd1 _02942_ sky130_fd_sc_hd__a21o_1
XFILLER_9_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08049__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10653_ net660 net145 vssd1 vssd1 vccd1 vccd1 _06271_ sky130_fd_sc_hd__and2_1
XANTENNA__09246__C1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16160_ net2494 _02370_ net1092 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[960\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_70_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13372_ top.CPU.control_unit.instruction\[17\] _02897_ net670 vssd1 vssd1 vccd1 vccd1
+ _02451_ sky130_fd_sc_hd__mux2_1
X_10584_ net410 _06196_ _06200_ _06204_ vssd1 vssd1 vccd1 vccd1 _06205_ sky130_fd_sc_hd__a31o_1
XFILLER_167_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload19 clknet_leaf_194_clk vssd1 vssd1 vccd1 vccd1 clkload19/Y sky130_fd_sc_hd__clkinv_8
XFILLER_5_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15111_ net1493 _01324_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r2_prev\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12323_ net2600 _04122_ net1191 vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__mux2_1
X_16091_ net2425 _02301_ net1209 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[891\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12482__A _03610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12148__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09549__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15042_ clknet_leaf_91_clk _01287_ vssd1 vssd1 vccd1 vccd1 top.SPI.percount\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_119_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12254_ net2866 net139 net433 vssd1 vssd1 vccd1 vccd1 _01427_ sky130_fd_sc_hd__mux2_1
XFILLER_123_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11356__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11205_ _06355_ net3570 net298 vssd1 vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__mux2_1
XANTENNA__11098__A net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12185_ net566 net363 _06667_ _06859_ _06858_ vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__a41o_1
XFILLER_150_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08959__X _04598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08772__A1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11136_ net514 _06254_ vssd1 vssd1 vccd1 vccd1 _06627_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_79_Left_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07980__C1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11067_ net323 _06253_ net534 net366 net2761 vssd1 vssd1 vccd1 vccd1 _02317_ sky130_fd_sc_hd__a32o_1
XFILLER_48_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15944_ net2278 _02154_ net1077 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[744\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_160_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10018_ _05399_ _05467_ net379 vssd1 vssd1 vccd1 vccd1 _05657_ sky130_fd_sc_hd__mux2_1
XFILLER_23_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15875_ net2209 _02085_ net1206 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[675\]
+ sky130_fd_sc_hd__dfrtp_1
X_14561__731 clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 net2200 sky130_fd_sc_hd__inv_2
XFILLER_63_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08288__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12657__A top.CPU.alu.program_counter\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11969_ _06522_ net342 net231 net3127 vssd1 vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_137_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_137_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_17_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14602__772 clknet_leaf_151_clk vssd1 vssd1 vccd1 vccd1 net2241 sky130_fd_sc_hd__inv_2
X_13708_ _03058_ net3710 vssd1 vssd1 vccd1 vccd1 _02625_ sky130_fd_sc_hd__nor2_1
XFILLER_44_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08383__S0 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_88_Left_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_158_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16427_ clknet_leaf_54_clk _00009_ net1135 vssd1 vssd1 vccd1 vccd1 top.I2C.I2C_state\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13639_ net3831 _07210_ net665 vssd1 vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__mux2_1
XANTENNA__09237__C1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16358_ clknet_leaf_32_clk _02567_ net1125 vssd1 vssd1 vccd1 vccd1 top.CPU.fetch.current_ra\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_158_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15309_ net1643 _01519_ net1058 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[109\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16289_ clknet_leaf_109_clk _02498_ net1240 vssd1 vssd1 vccd1 vccd1 top.CPU.data_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08460__B1 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12139__A2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11347__B1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13000__B net1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08212__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_97_Left_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout206 net211 vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__clkbuf_4
XFILLER_113_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout217 net219 vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__buf_4
X_09801_ _05437_ _05439_ net733 vssd1 vssd1 vccd1 vccd1 _05440_ sky130_fd_sc_hd__o21a_1
Xfanout228 _03191_ vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__buf_4
Xfanout239 net243 vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__buf_4
XANTENNA_clkload10_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07993_ top.CPU.registers.data\[824\] top.CPU.registers.data\[792\] net983 vssd1
+ vssd1 vccd1 vccd1 _03632_ sky130_fd_sc_hd__mux2_1
X_09732_ top.CPU.registers.data\[699\] top.CPU.registers.data\[667\] net827 vssd1
+ vssd1 vccd1 vccd1 _05371_ sky130_fd_sc_hd__mux2_1
XFILLER_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11455__B net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09663_ top.CPU.registers.data\[825\] net1336 net869 top.CPU.registers.data\[793\]
+ net710 vssd1 vssd1 vccd1 vccd1 _05302_ sky130_fd_sc_hd__o221a_1
XFILLER_28_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout273_A net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08614_ _03116_ _04248_ _04251_ _04252_ net611 vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__a311o_1
XFILLER_131_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09594_ _05232_ vssd1 vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__inv_2
XANTENNA__10873__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08545_ top.CPU.registers.data_out_r2_prev\[16\] net685 net619 _04183_ vssd1 vssd1
+ vccd1 vccd1 _04184_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout440_A net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_128_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_128_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1182_A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10086__A0 _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout159_X net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout538_A net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08476_ net913 _04103_ _04114_ net606 vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__a211o_1
XANTENNA__11190__B net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09228__C1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout705_A net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1068_X net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10389__A1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11586__B1 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11050__A2 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09028_ top.CPU.alu.program_counter\[8\] net1034 vssd1 vssd1 vccd1 vccd1 _04667_
+ sky130_fd_sc_hd__nor2_1
XFILLER_152_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout695_X net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11338__B1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08203__B1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold260 top.CPU.registers.data\[538\] vssd1 vssd1 vccd1 vccd1 net2817 sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 net60 vssd1 vssd1 vccd1 vccd1 net2828 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1402_X net1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold282 top.CPU.registers.data\[179\] vssd1 vssd1 vccd1 vccd1 net2839 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08754__A1 _04392_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07557__A2 _03180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold293 top.CPU.registers.data\[618\] vssd1 vssd1 vccd1 vccd1 net2850 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout862_X net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout740 net747 vssd1 vssd1 vccd1 vccd1 net740 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07962__C1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout751 net753 vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__clkbuf_4
Xfanout762 net763 vssd1 vssd1 vccd1 vccd1 net762 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12241__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14545__715 clknet_leaf_186_clk vssd1 vssd1 vccd1 vccd1 net2184 sky130_fd_sc_hd__inv_2
Xfanout773 net782 vssd1 vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_142_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout784 net786 vssd1 vssd1 vccd1 vccd1 net784 sky130_fd_sc_hd__buf_2
Xfanout795 net804 vssd1 vssd1 vccd1 vccd1 net795 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09703__B1 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12941_ _07380_ _07381_ vssd1 vssd1 vccd1 vccd1 _07382_ sky130_fd_sc_hd__nor2_1
XANTENNA__07714__C1 net1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15660_ net1994 _01870_ net1069 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[460\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12872_ _07317_ _07318_ vssd1 vssd1 vccd1 vccd1 _07319_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_83_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ _06510_ _06648_ net240 net158 net2893 vssd1 vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__a32o_1
X_15591_ net1925 _01801_ net1201 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[391\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_119_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_119_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_27_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09467__C1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11754_ _06593_ net499 net193 net3193 vssd1 vssd1 vccd1 vccd1 _01800_ sky130_fd_sc_hd__a22o_1
XFILLER_53_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10705_ net548 _05541_ _06318_ _06319_ vssd1 vssd1 vccd1 vccd1 _06320_ sky130_fd_sc_hd__o211a_1
XFILLER_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11685_ net456 _06506_ net234 net164 net3287 vssd1 vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__a32o_1
XANTENNA__16224__RESET_B net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16212_ net2546 _02422_ net1112 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[1012\]
+ sky130_fd_sc_hd__dfrtp_1
X_13424_ net1363 _02935_ net670 vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__mux2_1
X_10636_ net524 _06254_ vssd1 vssd1 vccd1 vccd1 _06255_ sky130_fd_sc_hd__nor2_1
XANTENNA__08690__A _04294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09234__A2 net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12924__B _03576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload108 clknet_leaf_153_clk vssd1 vssd1 vccd1 vccd1 clkload108/Y sky130_fd_sc_hd__inv_6
Xclkload119 clknet_leaf_184_clk vssd1 vssd1 vccd1 vccd1 clkload119/Y sky130_fd_sc_hd__inv_4
X_16143_ net2477 _02353_ net1095 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[943\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_128_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13355_ top.mmio.mem_data_i\[13\] net592 net1343 vssd1 vssd1 vccd1 vccd1 _02885_
+ sky130_fd_sc_hd__a21o_1
XFILLER_154_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10567_ top.CPU.fetch.current_ra\[14\] net1043 net634 top.CPU.handler.toreg\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06189_ sky130_fd_sc_hd__a22o_1
XFILLER_127_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08993__A1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07796__A2 net1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12306_ net4021 _05121_ net1235 vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__mux2_1
X_16074_ net2408 _02284_ net1085 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[874\]
+ sky130_fd_sc_hd__dfrtp_1
X_13286_ top.CPU.handler.readout _03126_ vssd1 vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__and2_1
X_10498_ _05521_ _06061_ _06122_ _06109_ net371 vssd1 vssd1 vccd1 vccd1 _06123_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_114_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15025_ clknet_leaf_83_clk net2786 net1261 vssd1 vssd1 vccd1 vccd1 top.SPI.parameters\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_114_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12237_ top.CPU.registers.data\[32\] net647 vssd1 vssd1 vccd1 vccd1 _06885_ sky130_fd_sc_hd__or2_1
XFILLER_46_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12940__A top.CPU.alu.program_counter\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12168_ top.CPU.registers.data\[68\] net651 net245 vssd1 vssd1 vccd1 vccd1 _06852_
+ sky130_fd_sc_hd__o21a_1
XFILLER_111_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07953__C1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11119_ net488 net464 _06617_ net303 net3537 vssd1 vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__a32o_1
XFILLER_7_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12099_ net3912 net652 _06817_ vssd1 vssd1 vccd1 vccd1 _01513_ sky130_fd_sc_hd__o21a_1
X_14288__458 clknet_leaf_196_clk vssd1 vssd1 vccd1 vccd1 net1927 sky130_fd_sc_hd__inv_2
XANTENNA__09026__A _04634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput6 DAT_I[13] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
X_15927_ net2261 _02137_ net1182 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[727\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11501__B1 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15858_ net2192 _02068_ net1106 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[658\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_92_774 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09313__X _04952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14329__499 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 net1968 sky130_fd_sc_hd__inv_2
X_15789_ net2123 _01999_ net1071 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[589\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_51_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11291__A net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08330_ top.CPU.registers.data\[243\] net1383 net988 top.CPU.registers.data\[211\]
+ net955 vssd1 vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__a221o_1
XANTENNA__08130__C1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13006__B1 _07431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08261_ top.CPU.registers.data\[246\] net1382 net998 top.CPU.registers.data\[214\]
+ net959 vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_138_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11280__A2 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13557__A1 _03000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08192_ net954 _03825_ _03827_ _03830_ vssd1 vssd1 vccd1 vccd1 _03831_ sky130_fd_sc_hd__a31o_1
XANTENNA__09225__A2 net1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10635__A net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11169__C net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08197__C1 net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14232__402 clknet_leaf_174_clk vssd1 vssd1 vccd1 vccd1 net1871 sky130_fd_sc_hd__inv_2
XFILLER_160_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1028_A net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout390_A net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10543__B2 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout488_A net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08759__B net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07944__C1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11740__B1 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10370__A net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07976_ top.CPU.registers.data\[24\] net983 _03614_ vssd1 vssd1 vccd1 vccd1 _03615_
+ sky130_fd_sc_hd__a21o_1
XFILLER_75_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09715_ net946 _05344_ _05345_ net609 vssd1 vssd1 vccd1 vccd1 _05354_ sky130_fd_sc_hd__a31o_1
XANTENNA__13493__A0 top.CPU.data_out\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12296__A1 _04531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11099__A2 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout655_A net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09697__C1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout276_X net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1397_A net1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09646_ _04394_ _04465_ _04395_ vssd1 vssd1 vccd1 vccd1 _05285_ sky130_fd_sc_hd__o21a_1
XFILLER_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09577_ net929 _05215_ _05212_ net624 vssd1 vssd1 vccd1 vccd1 _05216_ sky130_fd_sc_hd__a211o_1
XFILLER_82_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout443_X net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout822_A _03204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08528_ top.CPU.registers.data\[336\] net1290 net1011 top.CPU.registers.data\[368\]
+ net933 vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_61_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08121__C1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_5 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08459_ top.CPU.registers.data\[913\] net1302 net1023 top.CPU.registers.data\[945\]
+ net919 vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__a221o_1
XANTENNA__08672__B1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout610_X net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout708_X net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11470_ net3432 net264 net259 _06595_ vssd1 vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__a22o_1
XANTENNA__11559__B1 _06741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire448 _05397_ vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_98_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10421_ _05733_ _05822_ _05840_ _05753_ vssd1 vssd1 vccd1 vccd1 _06049_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_98_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13140_ top.SPI.command\[2\] top.CPU.data_out\[2\] net557 vssd1 vssd1 vccd1 vccd1
+ _01291_ sky130_fd_sc_hd__mux2_1
X_10352_ _05793_ _05978_ _05762_ vssd1 vssd1 vccd1 vccd1 _05983_ sky130_fd_sc_hd__a21oi_1
XFILLER_125_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13071_ top.CPU.data_out\[6\] net3050 net559 vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__mux2_1
X_10283_ _05362_ net507 vssd1 vssd1 vccd1 vccd1 _05916_ sky130_fd_sc_hd__nand2_1
XFILLER_140_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12022_ top.CPU.registers.data\[150\] net654 vssd1 vssd1 vccd1 vccd1 _06788_ sky130_fd_sc_hd__or2_1
XFILLER_104_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10534__A1 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11731__B1 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15270__RESET_B net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout570 net571 vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__clkbuf_4
Xfanout581 net582 vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07950__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout592 _02843_ vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__buf_2
XFILLER_65_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14016__186 clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 net1655 sky130_fd_sc_hd__inv_2
XANTENNA__09152__A1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12924_ top.CPU.alu.program_counter\[28\] _03576_ vssd1 vssd1 vccd1 vccd1 _07366_
+ sky130_fd_sc_hd__and2_1
X_15712_ net2046 _01922_ net1091 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[512\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_62_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12919__B top.CPU.alu.program_counter\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12855_ _07302_ _07303_ vssd1 vssd1 vccd1 vccd1 _07304_ sky130_fd_sc_hd__xnor2_1
X_15643_ net1977 _01853_ net1214 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[443\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11806_ net134 net3754 net157 vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__mux2_1
X_15574_ net1908 _01784_ net1221 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[374\]
+ sky130_fd_sc_hd__dfrtp_1
X_12786_ _07240_ _07241_ vssd1 vssd1 vccd1 vccd1 _07242_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11798__A0 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09455__A2 net1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08112__C1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ net133 net538 net500 net194 net2743 vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__a32o_1
XANTENNA__11262__A2 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12935__A top.CPU.alu.program_counter\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14673__843 clknet_leaf_188_clk vssd1 vssd1 vccd1 vccd1 net2312 sky130_fd_sc_hd__inv_2
XFILLER_30_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09207__A2 net1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11668_ _06481_ net210 net167 net3149 vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_116_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12654__B _05087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13407_ top.I2C.data_out\[27\] net555 _02922_ net598 vssd1 vssd1 vccd1 vccd1 _02923_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_116_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14923__Q top.CPU.alu.program_counter\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10619_ _04600_ _05281_ net446 vssd1 vssd1 vccd1 vccd1 _06238_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11014__A2 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09612__C1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11599_ _05847_ net3369 net215 vssd1 vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_133_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10222__B1 _05680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16126_ net2460 _02336_ net1237 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[926\]
+ sky130_fd_sc_hd__dfrtp_1
X_13338_ net668 net889 _02871_ _02872_ vssd1 vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__a31o_1
X_14714__884 clknet_leaf_164_clk vssd1 vssd1 vccd1 vccd1 net2353 sky130_fd_sc_hd__inv_2
XFILLER_142_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16057_ net2391 _02267_ net1225 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[857\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_142_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13269_ net3879 _02814_ _02819_ net1053 vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08179__C1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15008_ clknet_leaf_98_clk _01253_ net1254 vssd1 vssd1 vccd1 vccd1 top.SPI.parameters\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10525__A1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11722__B1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07926__C1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08194__A2 net1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11286__A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07830_ net705 _03467_ _03468_ vssd1 vssd1 vccd1 vccd1 _03469_ sky130_fd_sc_hd__or3_1
XFILLER_69_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07761_ net800 _03396_ _03397_ net730 vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__o211a_1
XANTENNA__13475__B1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09679__C1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09500_ net629 _05138_ net614 vssd1 vssd1 vccd1 vccd1 _05139_ sky130_fd_sc_hd__a21o_1
X_07692_ net1047 _03262_ vssd1 vssd1 vccd1 vccd1 _03331_ sky130_fd_sc_hd__and2_1
XFILLER_112_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09431_ net606 _05066_ _05069_ vssd1 vssd1 vccd1 vccd1 _05070_ sky130_fd_sc_hd__or3_1
XANTENNA__14922__RESET_B net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09362_ top.CPU.registers.data\[67\] net1297 net1018 top.CPU.registers.data\[99\]
+ net956 vssd1 vssd1 vccd1 vccd1 _05001_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_23_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11789__B1 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08103__C1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08313_ net749 _03950_ _03951_ net707 vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__o211a_1
X_09293_ top.CPU.registers.data\[164\] top.CPU.registers.data\[132\] net992 vssd1
+ vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__mux2_1
XFILLER_36_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout236_A net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07939__A _03544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08244_ net756 _03877_ _03878_ net779 vssd1 vssd1 vccd1 vccd1 _03883_ sky130_fd_sc_hd__o211a_1
XANTENNA__12564__B _06426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08175_ top.CPU.registers.data\[823\] top.CPU.registers.data\[791\] net824 vssd1
+ vssd1 vccd1 vccd1 _03814_ sky130_fd_sc_hd__mux2_1
XANTENNA__08406__B1 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout403_A net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10365__A _03916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1145_A net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11895__S net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10652__X _06270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1312_A net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout393_X net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout772_A net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11713__B1 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07917__C1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09382__A1 net1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08185__A2 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07932__A2 net1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13466__A0 top.CPU.handler.toreg\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12269__A1 _06428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13875__45 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 net1514 sky130_fd_sc_hd__inv_2
X_07959_ top.CPU.registers.data\[984\] net1319 net850 top.CPU.registers.data\[1016\]
+ net693 vssd1 vssd1 vccd1 vccd1 _03598_ sky130_fd_sc_hd__a221o_1
XANTENNA__09134__A1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_45 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10970_ net3740 net218 _06536_ net316 vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__a22o_1
XANTENNA__09685__A2 net1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13481__A3 _02932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08893__A0 top.CPU.alu.program_counter\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09629_ _05267_ vssd1 vssd1 vccd1 vccd1 _05268_ sky130_fd_sc_hd__inv_2
XFILLER_15_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout825_X net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11492__A2 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12640_ top.I2C.output_state\[7\] net2627 vssd1 vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__and2_1
X_14360__530 clknet_leaf_167_clk vssd1 vssd1 vccd1 vccd1 net1999 sky130_fd_sc_hd__inv_2
X_14657__827 clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 net2296 sky130_fd_sc_hd__inv_2
X_12571_ _06462_ _07075_ vssd1 vssd1 vccd1 vccd1 _07076_ sky130_fd_sc_hd__nand2_1
XANTENNA__08645__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12755__A top.CPU.alu.program_counter\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_50_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09842__C1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11522_ net3958 net252 _06736_ net488 vssd1 vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__a22o_1
XANTENNA__07999__A2 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15290_ net1624 _01500_ net1252 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[90\]
+ sky130_fd_sc_hd__dfrtp_1
X_14401__571 clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 net2040 sky130_fd_sc_hd__inv_2
XFILLER_8_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11453_ net146 net3544 net264 vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10404_ net601 _06031_ _06032_ vssd1 vssd1 vccd1 vccd1 _06033_ sky130_fd_sc_hd__a21o_4
XANTENNA__11547__A3 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09070__B1 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11384_ _06503_ net277 net271 net3410 vssd1 vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__a22o_1
XANTENNA__11952__B1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13123_ net2687 _02726_ net897 vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__mux2_1
X_10335_ _03789_ _05965_ vssd1 vssd1 vccd1 vccd1 _05966_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_111_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12490__A net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13054_ net2961 _07452_ net895 vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__mux2_1
X_10266_ net403 _05899_ vssd1 vssd1 vccd1 vccd1 _05900_ sky130_fd_sc_hd__and2_1
XANTENNA__11704__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1310 net1323 vssd1 vssd1 vccd1 vccd1 net1310 sky130_fd_sc_hd__clkbuf_2
X_12005_ net534 _06779_ vssd1 vssd1 vccd1 vccd1 _06780_ sky130_fd_sc_hd__nand2_8
XANTENNA__08176__A2 net1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1321 net1322 vssd1 vssd1 vccd1 vccd1 net1321 sky130_fd_sc_hd__clkbuf_4
Xfanout1332 net1333 vssd1 vssd1 vccd1 vccd1 net1332 sky130_fd_sc_hd__clkbuf_4
X_10197_ net309 _05750_ vssd1 vssd1 vccd1 vccd1 _05833_ sky130_fd_sc_hd__nand2_1
Xfanout1343 net1344 vssd1 vssd1 vccd1 vccd1 net1343 sky130_fd_sc_hd__buf_2
XANTENNA__11180__A1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1354 top.SPI.register\[1\] vssd1 vssd1 vccd1 vccd1 net1354 sky130_fd_sc_hd__buf_2
Xfanout1365 top.CPU.control_unit.instruction\[22\] vssd1 vssd1 vccd1 vccd1 net1365
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_120_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1376 net1377 vssd1 vssd1 vccd1 vccd1 net1376 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13457__B1 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1387 net1388 vssd1 vssd1 vccd1 vccd1 net1387 sky130_fd_sc_hd__buf_4
Xfanout1398 net1399 vssd1 vssd1 vccd1 vccd1 net1398 sky130_fd_sc_hd__clkbuf_2
XFILLER_94_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12907_ _07326_ _07331_ _07339_ _07340_ _07350_ vssd1 vssd1 vccd1 vccd1 _07351_ sky130_fd_sc_hd__o311a_1
XFILLER_34_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1035 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12680__A1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11483__A2 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12838_ _07287_ _07288_ vssd1 vssd1 vccd1 vccd1 _07289_ sky130_fd_sc_hd__nor2_1
X_15626_ net1960 _01836_ net1094 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[426\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_174_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09428__A2 net1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12955__A_N top.CPU.alu.program_counter\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11235__A2 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12769_ _07213_ _07218_ vssd1 vssd1 vccd1 vccd1 _07226_ sky130_fd_sc_hd__nand2b_1
X_15557_ net1891 _01767_ net1083 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[357\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09833__C1 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_41_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08100__A2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11786__A3 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15488_ net1822 _01698_ net1094 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[288\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput20 DAT_I[26] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
Xinput31 DAT_I[7] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
XFILLER_174_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12196__B1 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold804 top.CPU.registers.data\[273\] vssd1 vssd1 vccd1 vccd1 net3361 sky130_fd_sc_hd__dlygate4sd3_1
Xhold815 top.CPU.fetch.current_ra\[3\] vssd1 vssd1 vccd1 vccd1 net3372 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09600__A2 net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold826 top.CPU.registers.data\[324\] vssd1 vssd1 vccd1 vccd1 net3383 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11943__B1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold837 top.CPU.registers.data\[376\] vssd1 vssd1 vccd1 vccd1 net3394 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07611__A1 net1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold848 top.CPU.registers.data\[730\] vssd1 vssd1 vccd1 vccd1 net3405 sky130_fd_sc_hd__dlygate4sd3_1
X_16109_ net2443 _02319_ net1076 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[909\]
+ sky130_fd_sc_hd__dfrtp_1
X_09980_ _05055_ net377 vssd1 vssd1 vccd1 vccd1 _05619_ sky130_fd_sc_hd__nor2_1
XFILLER_104_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10913__A _06213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold859 top.CPU.registers.data\[502\] vssd1 vssd1 vccd1 vccd1 net3416 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08931_ top.CPU.registers.data\[330\] net1374 net975 top.CPU.registers.data\[362\]
+ net1281 vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__o221a_1
XANTENNA__11728__B net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_941 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08167__A2 net1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08862_ _04500_ net1363 net452 vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__mux2_1
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07914__A2 net1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07813_ top.CPU.registers.data\[605\] net1319 net850 top.CPU.registers.data\[637\]
+ net705 vssd1 vssd1 vccd1 vccd1 _03452_ sky130_fd_sc_hd__a221o_1
X_08793_ top.CPU.registers.data_out_r2_prev\[12\] net689 vssd1 vssd1 vccd1 vccd1 _04432_
+ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout186_A net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07744_ top.CPU.registers.data\[606\] net1333 net864 top.CPU.registers.data\[638\]
+ net755 vssd1 vssd1 vccd1 vccd1 _03383_ sky130_fd_sc_hd__a221o_1
XANTENNA__08529__S net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09667__A2 net1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08324__C1 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12120__B1 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14344__514 clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 net1983 sky130_fd_sc_hd__inv_2
XFILLER_53_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10277__A3 _05367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07675_ net632 _03297_ _03309_ vssd1 vssd1 vccd1 vccd1 _03314_ sky130_fd_sc_hd__or3_1
XFILLER_52_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11474__A2 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout353_A _06771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09414_ net797 _05045_ _05052_ net643 vssd1 vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__a211o_1
XANTENNA__10682__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12959__C1 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09345_ net708 _04981_ _04982_ _04983_ vssd1 vssd1 vccd1 vccd1 _04984_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout520_A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08627__B1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12575__A _05988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout141_X net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1262_A net1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_32_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout239_X net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout618_A net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_33_Left_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11777__A3 net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09276_ net926 _04893_ _04894_ net950 vssd1 vssd1 vccd1 vccd1 _04915_ sky130_fd_sc_hd__o211a_1
XANTENNA__08117__X _03756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10985__B2 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08227_ top.CPU.registers.data\[438\] top.CPU.registers.data\[406\] net829 vssd1
+ vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1050_X net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08158_ top.CPU.registers.data\[471\] net1325 net856 top.CPU.registers.data\[503\]
+ net773 vssd1 vssd1 vccd1 vccd1 _03797_ sky130_fd_sc_hd__a221o_1
XANTENNA__09052__B1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout987_A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08089_ top.CPU.registers.data\[693\] top.CPU.registers.data\[661\] net827 vssd1
+ vssd1 vccd1 vccd1 _03728_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1315_X net1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09095__S net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10120_ net407 net395 net417 vssd1 vssd1 vccd1 vccd1 _05758_ sky130_fd_sc_hd__o21a_1
XFILLER_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout775_X net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_99_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_99_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08158__A2 net1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_42_Left_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10051_ _03148_ net1045 net881 vssd1 vssd1 vccd1 vccd1 _05690_ sky130_fd_sc_hd__a21o_1
XFILLER_103_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11162__A1 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13952__122 clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 net1591 sky130_fd_sc_hd__inv_2
XANTENNA__07905__A2 _03541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout942_X net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09107__A1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13810_ net3343 net333 net326 top.CPU.data_out\[12\] vssd1 vssd1 vccd1 vccd1 _02690_
+ sky130_fd_sc_hd__a22o_1
XFILLER_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08315__C1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12469__B _03783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13741_ _03079_ _03080_ vssd1 vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__nor2_1
X_14087__257 clknet_leaf_184_clk vssd1 vssd1 vccd1 vccd1 net1726 sky130_fd_sc_hd__inv_2
XANTENNA__11465__A2 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10953_ net519 net442 net137 net545 vssd1 vssd1 vccd1 vccd1 _06527_ sky130_fd_sc_hd__and4_1
XFILLER_71_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08330__A2 net1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13672_ net3133 net331 net330 top.CPU.addressnew\[5\] vssd1 vssd1 vccd1 vccd1 _02600_
+ sky130_fd_sc_hd__a22o_1
X_16460_ clknet_leaf_87_clk _02622_ net1271 vssd1 vssd1 vccd1 vccd1 top.SPI.timem\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10884_ net494 net469 _06484_ net223 net3006 vssd1 vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__a32o_1
XANTENNA__08963__A _04567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_51_Left_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12623_ _03121_ top.I2C.I2C_state\[3\] net2715 vssd1 vssd1 vccd1 vccd1 _00033_ sky130_fd_sc_hd__a21o_1
XANTENNA__08618__A0 _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15411_ net1745 _01621_ net1184 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[211\]
+ sky130_fd_sc_hd__dfrtp_1
X_16391_ clknet_leaf_84_clk net2611 net1264 vssd1 vssd1 vccd1 vccd1 top.SPI.register\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11217__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14128__298 clknet_leaf_200_clk vssd1 vssd1 vccd1 vccd1 net1767 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_14_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09815__C1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_23_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_8
X_15342_ net1676 _01552_ net1190 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[142\]
+ sky130_fd_sc_hd__dfrtp_1
X_12554_ top.CPU.handler.state\[2\] top.CPU.handler.state\[0\] vssd1 vssd1 vccd1 vccd1
+ _07060_ sky130_fd_sc_hd__nor2_1
XANTENNA__11768__A3 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09830__A2 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11505_ _06638_ net260 net256 net3214 vssd1 vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__a22o_1
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15273_ net1607 _01483_ net1056 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[73\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12485_ _06990_ _06993_ _06992_ vssd1 vssd1 vccd1 vccd1 _06994_ sky130_fd_sc_hd__or3b_1
XANTENNA__09269__S1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09794__A _05399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11436_ net565 net136 net539 vssd1 vssd1 vccd1 vccd1 _06719_ sky130_fd_sc_hd__and3_1
XFILLER_171_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11925__B1 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08397__A2 net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11367_ _06475_ net277 net271 net3185 vssd1 vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__a22o_1
XFILLER_152_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13106_ _07426_ _02717_ top.SPI.count\[3\] _06946_ vssd1 vssd1 vccd1 vccd1 _02718_
+ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_60_Left_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10318_ net399 _05946_ vssd1 vssd1 vccd1 vccd1 _05950_ sky130_fd_sc_hd__nor2_1
XFILLER_3_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14785__955 clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 net2424 sky130_fd_sc_hd__inv_2
XANTENNA__11548__B net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11298_ net475 _06482_ net428 vssd1 vssd1 vccd1 vccd1 _06707_ sky130_fd_sc_hd__and3_1
XFILLER_26_1001 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13037_ top.SPI.parameters\[20\] top.SPI.paroutput\[12\] net1355 vssd1 vssd1 vccd1
+ vccd1 _07444_ sky130_fd_sc_hd__mux2_1
X_10249_ _05499_ net507 net510 _05501_ vssd1 vssd1 vccd1 vccd1 _05883_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__09018__B _04656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1140 net1146 vssd1 vssd1 vccd1 vccd1 net1140 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_128_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14031__201 clknet_leaf_191_clk vssd1 vssd1 vccd1 vccd1 net1670 sky130_fd_sc_hd__inv_2
XFILLER_67_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1151 net1153 vssd1 vssd1 vccd1 vccd1 net1151 sky130_fd_sc_hd__clkbuf_2
Xfanout1162 net1164 vssd1 vssd1 vccd1 vccd1 net1162 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_128_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14826__996 clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 net2465 sky130_fd_sc_hd__inv_2
XFILLER_39_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_163_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1173 net1179 vssd1 vssd1 vccd1 vccd1 net1173 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10900__A1 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13255__S _06948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1184 net1187 vssd1 vssd1 vccd1 vccd1 net1184 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16420__RESET_B net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1195 net1196 vssd1 vssd1 vccd1 vccd1 net1195 sky130_fd_sc_hd__clkbuf_4
XFILLER_54_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14988_ clknet_leaf_93_clk _01233_ net1267 vssd1 vssd1 vccd1 vccd1 top.SPI.paroutput\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08306__C1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_182_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11283__B _03170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11456__A2 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_62_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07460_ top.CPU.alu.program_counter\[2\] vssd1 vssd1 vccd1 vccd1 _03100_ sky130_fd_sc_hd__inv_2
XANTENNA__08952__S0 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15609_ net1943 _01819_ net1246 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[409\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_197_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09806__C1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10908__A _06190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_14_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_8
X_09130_ top.CPU.registers.data\[679\] top.CPU.registers.data\[647\] top.CPU.registers.data\[551\]
+ top.CPU.registers.data\[519\] net995 net919 vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_33_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_77_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09821__A2 net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09061_ top.CPU.registers.data\[424\] top.CPU.registers.data\[392\] top.CPU.registers.data\[296\]
+ top.CPU.registers.data\[264\] net975 net1281 vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__mux4_1
XANTENNA__07832__A1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_120_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08012_ top.CPU.alu.program_counter\[20\] net1034 vssd1 vssd1 vccd1 vccd1 _03651_
+ sky130_fd_sc_hd__or2_1
XFILLER_116_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13497__Y _02968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09034__B1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15302__RESET_B net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold601 top.CPU.registers.data\[31\] vssd1 vssd1 vccd1 vccd1 net3158 sky130_fd_sc_hd__dlygate4sd3_1
Xhold612 top.CPU.registers.data\[905\] vssd1 vssd1 vccd1 vccd1 net3169 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11916__B1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold623 top.CPU.registers.data\[539\] vssd1 vssd1 vccd1 vccd1 net3180 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09585__A1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold634 top.CPU.fetch.current_ra\[22\] vssd1 vssd1 vccd1 vccd1 net3191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold645 top.CPU.registers.data\[710\] vssd1 vssd1 vccd1 vccd1 net3202 sky130_fd_sc_hd__dlygate4sd3_1
Xhold656 _00031_ vssd1 vssd1 vccd1 vccd1 net3213 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07596__B1 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12561__C _06228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold667 top.CPU.registers.data\[711\] vssd1 vssd1 vccd1 vccd1 net3224 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09963_ _05436_ _05503_ _05597_ _05600_ vssd1 vssd1 vccd1 vccd1 _05602_ sky130_fd_sc_hd__a31oi_2
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold678 top.CPU.registers.data\[44\] vssd1 vssd1 vccd1 vccd1 net3235 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13669__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_135_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold689 top.CPU.registers.data\[718\] vssd1 vssd1 vccd1 vccd1 net3246 sky130_fd_sc_hd__dlygate4sd3_1
X_13936__106 clknet_leaf_194_clk vssd1 vssd1 vccd1 vccd1 net1575 sky130_fd_sc_hd__inv_2
XFILLER_134_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08914_ top.CPU.registers.data\[458\] net1313 net844 top.CPU.registers.data\[490\]
+ net765 vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_51_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09894_ _04599_ _04567_ vssd1 vssd1 vccd1 vccd1 _05533_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_51_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1010_A net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11144__A1 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_15_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1108_A net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1301 top.CPU.registers.data\[1005\] vssd1 vssd1 vccd1 vccd1 net3858 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08845_ top.CPU.registers.data\[43\] top.CPU.registers.data\[11\] net969 vssd1 vssd1
+ vccd1 vccd1 _04484_ sky130_fd_sc_hd__mux2_1
XANTENNA__07899__A1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1312 top.CPU.registers.data\[888\] vssd1 vssd1 vccd1 vccd1 net3869 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1323 top.CPU.registers.data\[1000\] vssd1 vssd1 vccd1 vccd1 net3880 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1334 top.I2C.within_byte_counter_writing\[2\] vssd1 vssd1 vccd1 vccd1 net3891
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout470_A _03194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1345 top.CPU.registers.data\[84\] vssd1 vssd1 vccd1 vccd1 net3902 sky130_fd_sc_hd__dlygate4sd3_1
X_13845__15 clknet_leaf_76_clk vssd1 vssd1 vccd1 vccd1 net1484 sky130_fd_sc_hd__inv_2
XANTENNA__08560__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout189_X net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout568_A net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1356 top.CPU.registers.data\[925\] vssd1 vssd1 vccd1 vccd1 net3913 sky130_fd_sc_hd__dlygate4sd3_1
X_08776_ top.CPU.registers.data\[460\] net1316 net847 top.CPU.registers.data\[492\]
+ net767 vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__a221o_1
Xhold1367 top.CPU.registers.data\[1\] vssd1 vssd1 vccd1 vccd1 net3924 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1378 top.CPU.registers.data\[65\] vssd1 vssd1 vccd1 vccd1 net3935 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_108_Left_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1389 top.CPU.registers.data\[112\] vssd1 vssd1 vccd1 vccd1 net3946 sky130_fd_sc_hd__dlygate4sd3_1
X_07727_ top.CPU.registers.data\[1023\] top.CPU.registers.data\[991\] top.CPU.registers.data\[959\]
+ top.CPU.registers.data\[927\] net999 net959 vssd1 vssd1 vccd1 vccd1 _03366_ sky130_fd_sc_hd__mux4_1
XANTENNA__10981__D_N net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11447__A2 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout356_X net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout735_A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11761__X _06760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08312__A2 net1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09879__A net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10655__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07658_ net1044 _03252_ _03292_ _03296_ vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_0_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08783__A net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout902_A net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_8_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_8_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout523_X net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07589_ top.CPU.registers.data\[447\] net1334 net865 top.CPU.registers.data\[415\]
+ net756 vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__o221a_1
XANTENNA__09499__S1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09328_ top.CPU.registers.data\[644\] net1329 net860 top.CPU.registers.data\[676\]
+ net726 vssd1 vssd1 vccd1 vccd1 _04967_ sky130_fd_sc_hd__a221o_1
XFILLER_139_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09812__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11080__A0 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09259_ top.CPU.registers.data\[837\] net1286 net1004 top.CPU.registers.data\[869\]
+ net926 vssd1 vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_117_Left_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12270_ net3924 _06518_ net434 vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__mux2_1
X_14472__642 clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 net2111 sky130_fd_sc_hd__inv_2
XFILLER_135_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14769__939 clknet_leaf_190_clk vssd1 vssd1 vccd1 vccd1 net2408 sky130_fd_sc_hd__inv_2
XANTENNA__11907__B1 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11221_ net3381 net294 _06665_ net484 vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__a22o_1
XFILLER_49_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12244__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11383__A1 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08784__C1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11152_ net489 net466 _06635_ net303 net3034 vssd1 vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__a32o_1
X_14513__683 clknet_leaf_187_clk vssd1 vssd1 vccd1 vccd1 net2152 sky130_fd_sc_hd__inv_2
XANTENNA__08023__A net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10103_ net415 _05664_ vssd1 vssd1 vccd1 vccd1 _05741_ sky130_fd_sc_hd__nor2_1
XFILLER_1_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11083_ net531 _05694_ _06519_ vssd1 vssd1 vccd1 vccd1 _06596_ sky130_fd_sc_hd__and3_1
X_15960_ net2294 _02170_ net1148 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[760\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08958__A net1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09423__S1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11135__B2 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08536__C1 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input31_A DAT_I[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10034_ _03243_ _05671_ vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_145_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10986__C_N net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12883__A1 top.CPU.alu.program_counter\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15891_ net2225 _02101_ net1186 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[691\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11686__A2 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12883__B2 top.CPU.alu.program_counter\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11438__A2 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11985_ _06545_ net350 net182 net2978 vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_86_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08303__A2 net1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09500__A1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16512_ clknet_leaf_58_clk _02674_ net1144 vssd1 vssd1 vccd1 vccd1 top.mmio.mem_data_i\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_86_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13724_ net3985 _03068_ vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__nor2_1
X_10936_ net148 net437 vssd1 vssd1 vccd1 vccd1 _06515_ sky130_fd_sc_hd__and2_1
XFILLER_32_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08693__A top.CPU.alu.program_counter\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07801__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16443_ clknet_leaf_85_clk _02606_ net1263 vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11831__B net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13655_ net3112 _07363_ net666 vssd1 vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__mux2_1
X_10867_ net496 net469 net520 _06473_ _06470_ vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__a41o_1
XFILLER_20_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12646__C _06948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12606_ top.SPI.timem\[13\] top.SPI.timem\[12\] top.SPI.timem\[15\] top.SPI.timem\[14\]
+ vssd1 vssd1 vccd1 vccd1 _07106_ sky130_fd_sc_hd__or4b_1
XFILLER_157_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08067__A1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13586_ top.CPU.alu.program_counter\[15\] _06171_ net1352 vssd1 vssd1 vccd1 vccd1
+ _03018_ sky130_fd_sc_hd__mux2_1
X_16374_ clknet_leaf_75_clk _02583_ net1159 vssd1 vssd1 vccd1 vccd1 top.CPU.fetch.current_ra\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_169_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10798_ _06403_ _06404_ _06407_ vssd1 vssd1 vccd1 vccd1 _06409_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_30_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09803__A2 net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12537_ _05527_ _05573_ _07045_ vssd1 vssd1 vccd1 vccd1 _07046_ sky130_fd_sc_hd__nand3_1
X_15325_ net1659 _01535_ net1114 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[125\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15256_ net1590 _01466_ net1102 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[56\]
+ sky130_fd_sc_hd__dfrtp_1
X_12468_ _03754_ _03783_ _03887_ _03915_ vssd1 vssd1 vccd1 vccd1 _06977_ sky130_fd_sc_hd__o22ai_1
XANTENNA__14931__Q top.CPU.alu.program_counter\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09567__A1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11419_ _06556_ net276 net267 net3219 vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__a22o_1
X_15187_ net1524 _01397_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r1_prev\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_12399_ net2780 _03129_ top.I2C.I2C_state\[21\] vssd1 vssd1 vccd1 vccd1 _00035_ sky130_fd_sc_hd__a21o_1
XFILLER_141_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11374__A1 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_165_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_3_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_39_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08527__C1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09316__X _04955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07772__A net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08630_ top.CPU.registers.data\[942\] top.CPU.registers.data\[910\] net819 vssd1
+ vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__mux2_1
XFILLER_66_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08079__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07750__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08561_ net740 _04198_ _04199_ net766 vssd1 vssd1 vccd1 vccd1 _04200_ sky130_fd_sc_hd__o211a_1
XANTENNA__11429__A2 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13823__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07512_ net1278 _03149_ vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__or2_1
XANTENNA__10637__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08492_ top.CPU.registers.data\[240\] net1390 net820 top.CPU.registers.data\[208\]
+ net770 vssd1 vssd1 vccd1 vccd1 _04131_ sky130_fd_sc_hd__a221o_1
XANTENNA__12329__S net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout149_A _06412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09255__B1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10419__A2_N net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09113_ top.CPU.registers.data\[839\] net1332 net864 top.CPU.registers.data\[871\]
+ net749 vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_44_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14456__626 clknet_leaf_170_clk vssd1 vssd1 vccd1 vccd1 net2095 sky130_fd_sc_hd__inv_2
XFILLER_164_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11601__A2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout316_A net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09044_ top.CPU.registers.data\[424\] top.CPU.registers.data\[392\] net811 vssd1
+ vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__mux2_1
X_14200__370 clknet_leaf_168_clk vssd1 vssd1 vccd1 vccd1 net1839 sky130_fd_sc_hd__inv_2
Xhold420 top.CPU.registers.data\[889\] vssd1 vssd1 vccd1 vccd1 net2977 sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 top.CPU.registers.data\[208\] vssd1 vssd1 vccd1 vccd1 net2988 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07569__B1 top.CPU.control_unit.instruction\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11365__A1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold442 top.CPU.registers.data\[8\] vssd1 vssd1 vccd1 vccd1 net2999 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1225_A net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold453 top.CPU.registers.data\[550\] vssd1 vssd1 vccd1 vccd1 net3010 sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 top.CPU.registers.data\[979\] vssd1 vssd1 vccd1 vccd1 net3021 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11188__B net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08230__A1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold475 top.CPU.registers.data\[436\] vssd1 vssd1 vccd1 vccd1 net3032 sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 top.CPU.registers.data\[685\] vssd1 vssd1 vccd1 vccd1 net3043 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout685_A net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout900 net901 vssd1 vssd1 vccd1 vccd1 net900 sky130_fd_sc_hd__clkbuf_4
Xfanout911 net914 vssd1 vssd1 vccd1 vccd1 net911 sky130_fd_sc_hd__clkbuf_4
Xhold497 top.CPU.registers.data\[314\] vssd1 vssd1 vccd1 vccd1 net3054 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout922 net924 vssd1 vssd1 vccd1 vccd1 net922 sky130_fd_sc_hd__clkbuf_4
XFILLER_104_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09946_ _04021_ _04051_ vssd1 vssd1 vccd1 vccd1 _05585_ sky130_fd_sc_hd__or2_1
Xfanout933 net934 vssd1 vssd1 vccd1 vccd1 net933 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1013_X net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11117__B2 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout944 net948 vssd1 vssd1 vccd1 vccd1 net944 sky130_fd_sc_hd__clkbuf_4
XFILLER_98_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout955 net962 vssd1 vssd1 vccd1 vccd1 net955 sky130_fd_sc_hd__buf_2
Xfanout966 net1003 vssd1 vssd1 vccd1 vccd1 net966 sky130_fd_sc_hd__clkbuf_4
Xfanout977 net978 vssd1 vssd1 vccd1 vccd1 net977 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11668__A2 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1120 net105 vssd1 vssd1 vccd1 vccd1 net3677 sky130_fd_sc_hd__dlygate4sd3_1
X_09877_ _03310_ net547 _03323_ vssd1 vssd1 vccd1 vccd1 _05516_ sky130_fd_sc_hd__and3_1
XANTENNA__10820__B net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout473_X net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout852_A net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout988 net989 vssd1 vssd1 vccd1 vccd1 net988 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1131 top.CPU.registers.data\[644\] vssd1 vssd1 vccd1 vccd1 net3688 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout999 net1002 vssd1 vssd1 vccd1 vccd1 net999 sky130_fd_sc_hd__clkbuf_4
Xhold1142 top.CPU.registers.data\[500\] vssd1 vssd1 vccd1 vccd1 net3699 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1153 _03059_ vssd1 vssd1 vccd1 vccd1 net3710 sky130_fd_sc_hd__dlygate4sd3_1
X_08828_ _04431_ _04464_ vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__and2_1
XFILLER_57_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1164 top.CPU.registers.data\[253\] vssd1 vssd1 vccd1 vccd1 net3721 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07741__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1175 top.CPU.registers.data\[981\] vssd1 vssd1 vccd1 vccd1 net3732 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1186 top.CPU.registers.data\[778\] vssd1 vssd1 vccd1 vccd1 net3743 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1197 top.CPU.registers.data\[343\] vssd1 vssd1 vccd1 vccd1 net3754 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout640_X net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08759_ top.CPU.registers.data\[748\] net1386 vssd1 vssd1 vccd1 vccd1 _04398_ sky130_fd_sc_hd__and2_1
XANTENNA__13814__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout738_X net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1382_X net1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10628__B1 _06141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07719__S1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11770_ net464 _06613_ net238 net162 net3271 vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__a32o_1
XANTENNA__12093__A2 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10721_ net532 _06335_ vssd1 vssd1 vccd1 vccd1 _06336_ sky130_fd_sc_hd__nor2_1
XFILLER_41_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11840__A2 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12239__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout905_X net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13440_ net3552 _02941_ net121 vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__mux2_1
X_10652_ net603 _06268_ _06269_ vssd1 vssd1 vccd1 vccd1 _06270_ sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_81_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09246__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10267__B _05793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_125_Left_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13371_ net889 _02896_ vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__and2_1
X_10583_ _05667_ _05787_ _05792_ _05671_ _06203_ vssd1 vssd1 vccd1 vccd1 _06204_ sky130_fd_sc_hd__o221a_1
XFILLER_167_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14199__369 clknet_leaf_171_clk vssd1 vssd1 vccd1 vccd1 net1838 sky130_fd_sc_hd__inv_2
XANTENNA__12763__A top.CPU.alu.program_counter\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15110_ net1492 _01323_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r2_prev\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_12322_ net2567 _04048_ net1103 vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10800__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16090_ net2424 _02300_ net1244 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[890\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_103_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12482__B _03645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15041_ clknet_leaf_90_clk _01286_ vssd1 vssd1 vccd1 vccd1 top.SPI.percount\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_126_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09549__A1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12253_ net2934 net141 net431 vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__mux2_1
XANTENNA__10283__A _05362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11204_ net492 _06510_ _06648_ net300 net2856 vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__a32o_1
XFILLER_123_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11098__B net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12184_ top.CPU.registers.data\[59\] net654 vssd1 vssd1 vccd1 vccd1 _06859_ sky130_fd_sc_hd__or2_1
X_11135_ net3756 net301 _06626_ net479 vssd1 vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__a22o_1
XFILLER_1_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08688__A _04294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07980__B1 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15943_ net2277 _02153_ net1197 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[743\]
+ sky130_fd_sc_hd__dfrtp_1
X_11066_ net324 _06230_ net536 net367 net2691 vssd1 vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__a32o_1
XANTENNA__11659__A2 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09182__C1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10017_ net384 _05655_ _05653_ net391 vssd1 vssd1 vccd1 vccd1 _05656_ sky130_fd_sc_hd__o211a_1
XANTENNA__08524__A2 net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09721__A1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07732__A0 _03370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15874_ net2208 _02084_ net1171 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[674\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_36_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_121_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10619__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12084__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11968_ _06521_ net351 net232 net3308 vssd1 vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__a22o_1
XANTENNA__12657__B _05156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13707_ top.SPI.timem\[5\] _03056_ net3709 vssd1 vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__a21oi_1
XANTENNA__14926__Q top.CPU.alu.program_counter\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08383__S1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14143__313 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 net1782 sky130_fd_sc_hd__inv_2
X_10919_ net660 net145 net435 vssd1 vssd1 vccd1 vccd1 _06505_ sky130_fd_sc_hd__and3_1
XFILLER_149_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11899_ net475 _05695_ net239 net186 net2759 vssd1 vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__a32o_1
X_16426_ clknet_leaf_56_clk _00008_ net1141 vssd1 vssd1 vccd1 vccd1 top.I2C.I2C_state\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_158_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13638_ net2935 _07193_ net664 vssd1 vssd1 vccd1 vccd1 _02572_ sky130_fd_sc_hd__mux2_1
XANTENNA__09237__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10177__B net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16357_ clknet_leaf_28_clk _02566_ net1148 vssd1 vssd1 vccd1 vccd1 top.CPU.fetch.current_ra\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13569_ top.CPU.alu.program_counter\[8\] net1350 net582 vssd1 vssd1 vccd1 vccd1 _03008_
+ sky130_fd_sc_hd__o21a_1
XFILLER_74_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09458__S net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07767__A _03405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15308_ net1642 _01518_ net1071 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[108\]
+ sky130_fd_sc_hd__dfrtp_1
X_16288_ clknet_leaf_64_clk net2558 net1163 vssd1 vssd1 vccd1 vccd1 top.CPU.counter_on
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08215__X _03854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13336__A2 _07089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15239_ net1573 _01449_ net1195 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_172_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08212__A1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08763__A2 net1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout207 net211 vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__clkbuf_2
X_09800_ top.CPU.registers.data\[538\] net867 net698 _05438_ vssd1 vssd1 vccd1 vccd1
+ _05439_ sky130_fd_sc_hd__o211a_1
Xfanout218 net219 vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__buf_6
XANTENNA__10921__A net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout229 _06772_ vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__buf_6
XFILLER_86_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07992_ top.CPU.registers.data\[984\] net1289 net1009 top.CPU.registers.data\[1016\]
+ net906 vssd1 vssd1 vccd1 vccd1 _03631_ sky130_fd_sc_hd__a221o_1
XFILLER_101_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_163_Right_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09731_ net797 _05368_ _05369_ net727 vssd1 vssd1 vccd1 vccd1 _05370_ sky130_fd_sc_hd__o211a_1
XANTENNA__07658__B_N _03252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09662_ top.CPU.alu.program_counter\[25\] net1036 vssd1 vssd1 vccd1 vccd1 _05301_
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_2_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10858__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10322__A2 _05685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08613_ net1367 _04244_ _04243_ top.CPU.control_unit.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 _04252_ sky130_fd_sc_hd__o211a_1
XFILLER_55_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09593_ net1378 net1038 _05231_ vssd1 vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__o21ai_4
X_08544_ net676 _04177_ _04178_ _04182_ net616 vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__a311o_1
XANTENNA__12567__B _06288_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10086__A1 _04225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08475_ net955 _04105_ _04104_ net938 vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout433_A _06602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11822__A2 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1175_A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09228__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11035__B1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09779__A1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13575__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout221_X net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout319_X net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09027_ _04634_ _04663_ vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__or2_1
XANTENNA__11199__A net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10307__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold250 top.CPU.registers.data\[4\] vssd1 vssd1 vccd1 vccd1 net2807 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09400__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold261 top.CPU.registers.data\[432\] vssd1 vssd1 vccd1 vccd1 net2818 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_160_950 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout590_X net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold272 _02598_ vssd1 vssd1 vccd1 vccd1 net2829 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout688_X net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold283 top.CPU.registers.data\[166\] vssd1 vssd1 vccd1 vccd1 net2840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 top.CPU.registers.data\[676\] vssd1 vssd1 vccd1 vccd1 net2851 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10390__X _06019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout730 net734 vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__buf_2
Xfanout741 net747 vssd1 vssd1 vccd1 vccd1 net741 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07962__B1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09929_ _04468_ _05567_ _05538_ vssd1 vssd1 vccd1 vccd1 _05568_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_130_Right_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout752 net753 vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__clkbuf_4
XFILLER_77_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_142_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout763 net764 vssd1 vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__clkbuf_2
X_14584__754 clknet_leaf_169_clk vssd1 vssd1 vccd1 vccd1 net2223 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_142_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout855_X net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout774 net782 vssd1 vssd1 vccd1 vccd1 net774 sky130_fd_sc_hd__clkbuf_2
Xfanout785 net786 vssd1 vssd1 vccd1 vccd1 net785 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09164__C1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout796 net804 vssd1 vssd1 vccd1 vccd1 net796 sky130_fd_sc_hd__clkbuf_4
X_12940_ top.CPU.alu.program_counter\[29\] top.CPU.alu.program_counter\[28\] top.CPU.alu.program_counter\[27\]
+ _07346_ vssd1 vssd1 vccd1 vccd1 _07381_ sky130_fd_sc_hd__and4_1
XFILLER_18_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08911__C1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11933__Y _06772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12871_ top.CPU.alu.program_counter\[23\] _03823_ vssd1 vssd1 vccd1 vccd1 _07318_
+ sky130_fd_sc_hd__nand2_1
X_14625__795 clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 net2264 sky130_fd_sc_hd__inv_2
XANTENNA__11662__A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11822_ _06658_ net233 net156 net3377 vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_83_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09467__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15590_ net1924 _01800_ net1080 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[390\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12066__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13263__B2 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11753_ _06592_ net206 net195 net3025 vssd1 vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__a22o_1
XFILLER_92_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10704_ _04797_ net508 net503 _04796_ net443 vssd1 vssd1 vccd1 vccd1 _06319_ sky130_fd_sc_hd__o221a_1
X_11684_ net457 _06505_ net233 net164 net2910 vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__a32o_1
XANTENNA__08971__A net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16211_ net2545 _02421_ net1177 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[1011\]
+ sky130_fd_sc_hd__dfrtp_1
X_13423_ net889 _02934_ vssd1 vssd1 vccd1 vccd1 _02935_ sky130_fd_sc_hd__and2_1
XFILLER_14_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10635_ net551 net501 net142 vssd1 vssd1 vccd1 vccd1 _06254_ sky130_fd_sc_hd__or3b_1
XFILLER_14_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08978__C1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload109 clknet_leaf_154_clk vssd1 vssd1 vccd1 vccd1 clkload109/Y sky130_fd_sc_hd__inv_4
X_13354_ top.CPU.control_unit.instruction\[12\] _02884_ net671 vssd1 vssd1 vccd1 vccd1
+ _02446_ sky130_fd_sc_hd__mux2_1
X_16142_ net2476 _02352_ net1107 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[942\]
+ sky130_fd_sc_hd__dfrtp_1
X_10566_ net447 _06154_ _06176_ _06187_ vssd1 vssd1 vccd1 vccd1 _06188_ sky130_fd_sc_hd__a31o_1
XANTENNA__08442__A1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11041__A3 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10785__C1 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12305_ net2579 _05054_ net1185 vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__mux2_1
X_13285_ net1354 net1410 _06917_ vssd1 vssd1 vccd1 vccd1 _01409_ sky130_fd_sc_hd__o21a_1
XFILLER_127_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16073_ net2407 _02283_ net1055 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[873\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_170_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10497_ _05293_ _05583_ _06060_ vssd1 vssd1 vccd1 vccd1 _06122_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_114_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15024_ clknet_leaf_93_clk _01269_ net1267 vssd1 vssd1 vccd1 vccd1 top.SPI.parameters\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_142_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12236_ net475 _06698_ _06884_ net171 net3242 vssd1 vssd1 vccd1 vccd1 _01443_ sky130_fd_sc_hd__a32o_1
XFILLER_142_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12167_ net3950 net172 _06851_ _06738_ vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__a22o_1
XANTENNA__10741__A net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11118_ net574 net528 net440 net132 vssd1 vssd1 vccd1 vccd1 _06617_ sky130_fd_sc_hd__and4_1
X_12098_ net565 net362 _06632_ net178 top.CPU.registers.data\[103\] vssd1 vssd1 vccd1
+ vccd1 _06817_ sky130_fd_sc_hd__a32o_1
XANTENNA__12004__Y _06779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15926_ net2260 _02136_ net1227 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[726\]
+ sky130_fd_sc_hd__dfrtp_1
X_11049_ net530 _05694_ _06487_ vssd1 vssd1 vccd1 vccd1 _06583_ sky130_fd_sc_hd__and3_1
XFILLER_77_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput7 DAT_I[14] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11501__A1 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08902__C1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09741__S net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15857_ net2191 _02067_ net1192 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[657\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11572__A net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12057__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13254__B2 _02803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15788_ net2122 _01998_ net1071 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[588\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11804__A2 _06648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08260_ top.CPU.registers.data\[182\] net1382 net998 top.CPU.registers.data\[150\]
+ net681 vssd1 vssd1 vccd1 vccd1 _03899_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_138_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16409_ clknet_leaf_55_clk net2716 net1134 vssd1 vssd1 vccd1 vccd1 top.I2C.I2C_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07768__Y _03407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08191_ net679 _03828_ _03829_ net606 vssd1 vssd1 vccd1 vccd1 _03830_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_41_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12765__A0 top.CPU.alu.program_counter\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08433__A1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10635__B net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08984__A2 net1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14271__441 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 net1910 sky130_fd_sc_hd__inv_2
XANTENNA__09394__C1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14568__738 clknet_leaf_129_clk vssd1 vssd1 vccd1 vccd1 net2207 sky130_fd_sc_hd__inv_2
XFILLER_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10543__A2 _06141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07944__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15916__RESET_B net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07975_ top.CPU.registers.data\[56\] net1010 net934 vssd1 vssd1 vccd1 vccd1 _03614_
+ sky130_fd_sc_hd__a21o_1
X_14312__482 clknet_leaf_129_clk vssd1 vssd1 vccd1 vccd1 net1951 sky130_fd_sc_hd__inv_2
XFILLER_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09714_ net682 _05341_ _05342_ net922 vssd1 vssd1 vccd1 vccd1 _05353_ sky130_fd_sc_hd__o211a_1
XANTENNA__13493__A1 _04792_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14609__779 clknet_leaf_188_clk vssd1 vssd1 vccd1 vccd1 net2248 sky130_fd_sc_hd__inv_2
XFILLER_67_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09697__B1 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09161__A2 net1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09645_ _04603_ _05280_ _05283_ _05282_ vssd1 vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout171_X net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1292_A net1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout269_X net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout648_A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12048__A2 _06779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09576_ _05213_ _05214_ net951 vssd1 vssd1 vccd1 vccd1 _05215_ sky130_fd_sc_hd__mux2_1
XANTENNA__12297__B _06887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08527_ top.CPU.registers.data\[464\] net1290 net1011 top.CPU.registers.data\[496\]
+ net907 vssd1 vssd1 vccd1 vccd1 _04166_ sky130_fd_sc_hd__a221o_1
XANTENNA__13796__A2 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout815_A net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout436_X net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09887__A _03407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08458_ top.CPU.registers.data\[817\] top.CPU.registers.data\[785\] net995 vssd1
+ vssd1 vccd1 vccd1 _04097_ sky130_fd_sc_hd__mux2_1
XFILLER_168_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12584__Y _07088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout603_X net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07880__C1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08389_ top.CPU.registers.data\[562\] top.CPU.registers.data\[530\] net982 vssd1
+ vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__mux2_1
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10420_ net549 _03723_ net504 _03719_ _06047_ vssd1 vssd1 vccd1 vccd1 _06048_ sky130_fd_sc_hd__o221a_1
XANTENNA__11559__B2 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1036 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12220__A2 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09621__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10351_ net412 _05752_ vssd1 vssd1 vccd1 vccd1 _05982_ sky130_fd_sc_hd__or2_1
XFILLER_3_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12508__B1 _04291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10782__A2 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13070_ top.CPU.data_out\[5\] net3221 net558 vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__mux2_1
X_10282_ _05793_ _05914_ net224 vssd1 vssd1 vccd1 vccd1 _05915_ sky130_fd_sc_hd__a21oi_1
XFILLER_105_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12021_ top.CPU.registers.data\[150\] _06781_ vssd1 vssd1 vccd1 vccd1 _06787_ sky130_fd_sc_hd__and2_1
XANTENNA__12252__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout560 net561 vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__clkbuf_4
XFILLER_47_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09137__C1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout571 _03175_ vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__clkbuf_4
Xfanout582 net583 vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__clkbuf_2
Xfanout593 _02843_ vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09688__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10298__A1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15711_ net2045 _01921_ net1219 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[511\]
+ sky130_fd_sc_hd__dfrtp_1
X_12923_ top.CPU.alu.program_counter\[28\] _07362_ vssd1 vssd1 vccd1 vccd1 _07365_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__11495__B1 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07699__C1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08360__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15642_ net1976 _01852_ net1251 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[442\]
+ sky130_fd_sc_hd__dfrtp_1
X_12854_ top.CPU.alu.program_counter\[20\] _03685_ _07296_ vssd1 vssd1 vccd1 vccd1
+ _07303_ sky130_fd_sc_hd__a21oi_1
XFILLER_15_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13787__A2 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11805_ _05962_ net3744 net159 vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__mux2_1
XANTENNA__11247__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15573_ net1907 _01783_ net1215 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[373\]
+ sky130_fd_sc_hd__dfrtp_1
X_12785_ top.CPU.alu.program_counter\[14\] _07228_ vssd1 vssd1 vccd1 vccd1 _07241_
+ sky130_fd_sc_hd__nor2_1
XFILLER_15_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08112__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07869__X _03508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11736_ _06582_ net499 net193 net3428 vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_155_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09860__B1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08905__S net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12935__B _03477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11667_ net135 net3591 net166 vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__mux2_1
XFILLER_30_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13406_ top.mmio.mem_data_i\[27\] net593 net1346 vssd1 vssd1 vccd1 vccd1 _02922_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_116_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10618_ _04601_ _06234_ _06236_ net511 _05283_ vssd1 vssd1 vccd1 vccd1 _06237_ sky130_fd_sc_hd__a221o_1
XANTENNA__09612__B1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12211__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11598_ _05808_ net3249 net212 vssd1 vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__mux2_1
XFILLER_128_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10222__A1 _05429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08966__A2 net1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16125_ net2459 _02335_ net1119 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[925\]
+ sky130_fd_sc_hd__dfrtp_1
X_10549_ top.CPU.fetch.current_ra\[15\] net1043 net634 top.CPU.handler.toreg\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06172_ sky130_fd_sc_hd__a22o_1
XFILLER_127_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13337_ net668 net1407 vssd1 vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__and2b_1
X_14255__425 clknet_leaf_178_clk vssd1 vssd1 vccd1 vccd1 net1894 sky130_fd_sc_hd__inv_2
XANTENNA__10773__A2 _05685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16056_ net2390 _02266_ net1120 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[856\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_131_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13268_ top.I2C.data_out\[2\] net891 _02780_ vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__mux2_1
X_15007_ clknet_leaf_95_clk _01252_ net1260 vssd1 vssd1 vccd1 vccd1 top.SPI.parameters\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09915__A1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09376__C1 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12219_ net3289 net168 _06876_ vssd1 vssd1 vccd1 vccd1 _01452_ sky130_fd_sc_hd__a21o_1
X_13199_ top.I2C.output_state\[28\] _02773_ vssd1 vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__nand2_2
XFILLER_37_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10525__A2 _06147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09391__A2 net1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11286__B _05693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09128__C1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07760_ top.CPU.registers.data\[350\] net1333 net864 top.CPU.registers.data\[382\]
+ net781 vssd1 vssd1 vccd1 vccd1 _03399_ sky130_fd_sc_hd__a221o_1
XFILLER_38_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13475__A1 net1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09143__A2 net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15909_ net2243 _02119_ net1083 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[709\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11486__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07691_ net632 net547 _03328_ _03312_ _03317_ vssd1 vssd1 vccd1 vccd1 _03330_ sky130_fd_sc_hd__a2111o_1
XFILLER_64_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_200_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_200_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09430_ net954 _05068_ _05067_ net936 vssd1 vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__o211a_1
XFILLER_25_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09361_ top.CPU.registers.data\[35\] top.CPU.registers.data\[3\] net990 vssd1 vssd1
+ vccd1 vccd1 _05000_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11789__A1 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08312_ top.CPU.registers.data\[915\] net1327 net858 top.CPU.registers.data\[947\]
+ net724 vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__a221o_1
X_09292_ top.CPU.registers.data\[36\] net1020 net940 vssd1 vssd1 vccd1 vccd1 _04931_
+ sky130_fd_sc_hd__a21o_1
X_08243_ net799 _03875_ _03876_ _03881_ vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout131_A _06464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout229_A _06772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12564__C _06445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08174_ net748 _03811_ _03812_ net695 vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__o211a_1
XFILLER_119_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07658__C _03292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10365__B net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11410__B1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1040_A net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout598_A _07088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09367__C1 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08709__A2 net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10381__A net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1305_A net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07917__B1 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout386_X net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout765_A net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07958_ top.CPU.registers.data\[920\] net1321 net852 top.CPU.registers.data\[952\]
+ net694 vssd1 vssd1 vccd1 vccd1 _03597_ sky130_fd_sc_hd__a221o_1
XANTENNA__08786__A net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07889_ top.CPU.registers.data\[444\] top.CPU.registers.data\[412\] net833 vssd1
+ vssd1 vccd1 vccd1 _03528_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout932_A net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1295_X net1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09628_ net377 _05266_ vssd1 vssd1 vccd1 vccd1 _05267_ sky130_fd_sc_hd__and2_1
XFILLER_16_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08893__A1 _04531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09559_ top.CPU.registers.data\[576\] net1293 net1004 top.CPU.registers.data\[608\]
+ net928 vssd1 vssd1 vccd1 vccd1 _05198_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout720_X net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout818_X net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14696__866 clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 net2335 sky130_fd_sc_hd__inv_2
XANTENNA__13631__S net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12570_ _06067_ _06081_ _06103_ _07074_ vssd1 vssd1 vccd1 vccd1 _07075_ sky130_fd_sc_hd__a211oi_1
XFILLER_23_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11521_ net134 net356 vssd1 vssd1 vccd1 vccd1 _06736_ sky130_fd_sc_hd__and2_1
XFILLER_168_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12247__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11452_ net140 net3654 net263 vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__mux2_1
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14239__409 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 net1878 sky130_fd_sc_hd__inv_2
XANTENNA__08026__A net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10403_ top.CPU.fetch.current_ra\[21\] net1041 net883 top.CPU.handler.toreg\[21\]
+ vssd1 vssd1 vccd1 vccd1 _06032_ sky130_fd_sc_hd__a22o_1
XANTENNA__11401__B1 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11383_ net479 net471 _06502_ net271 net2997 vssd1 vssd1 vccd1 vccd1 _02127_ sky130_fd_sc_hd__a32o_1
XFILLER_152_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12771__A top.CPU.alu.program_counter\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10755__A2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13122_ top.SPI.command\[7\] net1410 top.SPI.paroutput\[31\] net1356 vssd1 vssd1
+ vccd1 vccd1 _02726_ sky130_fd_sc_hd__a22o_1
X_10334_ _04054_ _05964_ _03722_ _03988_ vssd1 vssd1 vccd1 vccd1 _05965_ sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_111_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09358__C1 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13053_ top.SPI.parameters\[28\] top.SPI.paroutput\[20\] net1357 vssd1 vssd1 vccd1
+ vccd1 _07452_ sky130_fd_sc_hd__mux2_1
XFILLER_127_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10265_ net396 _05886_ _05898_ _05738_ vssd1 vssd1 vccd1 vccd1 _05899_ sky130_fd_sc_hd__o22a_1
XFILLER_106_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10507__A2 _05937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07908__B1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1300 net1301 vssd1 vssd1 vccd1 vccd1 net1300 sky130_fd_sc_hd__clkbuf_2
X_12004_ net1401 _06751_ vssd1 vssd1 vccd1 vccd1 _06779_ sky130_fd_sc_hd__nor2_8
XFILLER_78_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1311 net1312 vssd1 vssd1 vccd1 vccd1 net1311 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09373__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10196_ _03316_ _03581_ net505 _03579_ _05831_ vssd1 vssd1 vccd1 vccd1 _05832_ sky130_fd_sc_hd__o221a_1
XFILLER_39_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1322 net1323 vssd1 vssd1 vccd1 vccd1 net1322 sky130_fd_sc_hd__buf_2
XFILLER_120_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1333 net1338 vssd1 vssd1 vccd1 vccd1 net1333 sky130_fd_sc_hd__clkbuf_4
Xfanout1344 net1345 vssd1 vssd1 vccd1 vccd1 net1344 sky130_fd_sc_hd__buf_1
XFILLER_120_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08581__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1355 top.SPI.state\[2\] vssd1 vssd1 vccd1 vccd1 net1355 sky130_fd_sc_hd__clkbuf_4
XFILLER_94_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1366 net1368 vssd1 vssd1 vccd1 vccd1 net1366 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13457__A1 net1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12710__S net1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1377 net1380 vssd1 vssd1 vccd1 vccd1 net1377 sky130_fd_sc_hd__clkbuf_4
Xfanout390 net392 vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__clkbuf_4
XFILLER_19_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1388 net1395 vssd1 vssd1 vccd1 vccd1 net1388 sky130_fd_sc_hd__clkbuf_4
XFILLER_94_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1399 top.CPU.control_unit.instruction\[13\] vssd1 vssd1 vccd1 vccd1 net1399
+ sky130_fd_sc_hd__buf_2
XANTENNA__11468__A0 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_109_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14640__810 clknet_leaf_199_clk vssd1 vssd1 vccd1 vccd1 net2279 sky130_fd_sc_hd__inv_2
XFILLER_47_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_109_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12906_ _07348_ _07349_ vssd1 vssd1 vccd1 vccd1 _07350_ sky130_fd_sc_hd__nor2_1
XFILLER_34_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkload7_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10691__A1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15625_ net1959 _01835_ net1061 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[425\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_174_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12837_ top.CPU.alu.program_counter\[18\] _07270_ top.CPU.alu.program_counter\[19\]
+ vssd1 vssd1 vccd1 vccd1 _07288_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_174_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15556_ net1890 _01766_ net1186 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[356\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08097__C1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08636__A1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12768_ _07223_ _07224_ vssd1 vssd1 vccd1 vccd1 _07225_ sky130_fd_sc_hd__or2_1
XFILLER_148_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_170_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11640__B1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11719_ _06559_ net198 net420 net2721 vssd1 vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__a22o_1
XANTENNA__07844__C1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15487_ net1821 _01697_ net1223 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[287\]
+ sky130_fd_sc_hd__dfrtp_1
X_12699_ net125 _07162_ net1360 vssd1 vssd1 vccd1 vccd1 _07163_ sky130_fd_sc_hd__o21a_1
XFILLER_174_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput10 DAT_I[17] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
Xinput21 DAT_I[27] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__buf_1
Xinput32 DAT_I[8] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12196__A1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold805 top.CPU.registers.data\[692\] vssd1 vssd1 vccd1 vccd1 net3362 sky130_fd_sc_hd__dlygate4sd3_1
Xhold816 top.SPI.parameters\[14\] vssd1 vssd1 vccd1 vccd1 net3373 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_max_cap449_X net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16108_ net2442 _02318_ net1076 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[908\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold827 top.CPU.registers.data\[156\] vssd1 vssd1 vccd1 vccd1 net3384 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold838 top.CPU.registers.data\[383\] vssd1 vssd1 vccd1 vccd1 net3395 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold849 top.CPU.registers.data\[346\] vssd1 vssd1 vccd1 vccd1 net3406 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10913__B net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08930_ top.CPU.registers.data\[458\] net1374 net972 top.CPU.registers.data\[490\]
+ net1365 vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__o221a_1
X_16039_ net2373 _02249_ net1199 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[839\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12499__A2 _05054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11728__C net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09364__A2 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08021__C1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08861_ net688 _04497_ _04498_ vssd1 vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__a21oi_1
XFILLER_96_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07812_ top.CPU.registers.data\[829\] net1389 net817 top.CPU.registers.data\[797\]
+ net692 vssd1 vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__a221o_1
X_08792_ net879 net450 _04429_ vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__o21a_1
XFILLER_42_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11459__A0 _06212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07743_ net700 _03381_ vssd1 vssd1 vccd1 vccd1 _03382_ sky130_fd_sc_hd__nand2_1
XFILLER_84_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08324__B1 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14383__553 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 net2022 sky130_fd_sc_hd__inv_2
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout179_A _06795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07674_ _03271_ _03284_ vssd1 vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__nor2_2
XFILLER_26_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08893__X _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10682__A1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09413_ _05048_ _05051_ net1308 vssd1 vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__o21a_1
XFILLER_53_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout346_A _06771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13304__X _02847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09344_ net697 _04979_ _04980_ net637 vssd1 vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__a31o_1
XANTENNA__08088__C1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14424__594 clknet_leaf_170_clk vssd1 vssd1 vccd1 vccd1 net2063 sky130_fd_sc_hd__inv_2
XFILLER_40_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09275_ net950 _04895_ _04913_ net605 vssd1 vssd1 vccd1 vccd1 _04914_ sky130_fd_sc_hd__a211o_1
XANTENNA__11631__B1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10376__A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout513_A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10985__A2 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08226_ top.CPU.registers.data\[246\] net1392 net835 top.CPU.registers.data\[214\]
+ net779 vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__a221o_1
XFILLER_119_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10095__B _05643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07850__A2 net1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08157_ top.CPU.registers.data\[439\] top.CPU.registers.data\[407\] net824 vssd1
+ vssd1 vccd1 vccd1 _03796_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout301_X net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1043_X net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_56_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08088_ net798 _03725_ _03726_ net726 vssd1 vssd1 vccd1 vccd1 _03727_ sky130_fd_sc_hd__o211a_1
XANTENNA__08260__C1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07602__A2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout882_A net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15249__RESET_B net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1308_X net1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10050_ _03148_ net1045 net881 vssd1 vssd1 vccd1 vccd1 _05689_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11698__B1 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout670_X net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13991__161 clknet_leaf_183_clk vssd1 vssd1 vccd1 vccd1 net1630 sky130_fd_sc_hd__inv_2
XFILLER_57_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11162__A2 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout768_X net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout935_X net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13740_ top.SPI.timem\[17\] top.SPI.timem\[18\] _03077_ vssd1 vssd1 vccd1 vccd1 _03080_
+ sky130_fd_sc_hd__and3_1
X_10952_ net3307 net218 _06526_ net320 vssd1 vssd1 vccd1 vccd1 _02369_ sky130_fd_sc_hd__a22o_1
XFILLER_84_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10673__A1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13671_ net2951 net331 net330 top.CPU.addressnew\[4\] vssd1 vssd1 vccd1 vccd1 _02599_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11870__B1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12766__A top.CPU.alu.program_counter\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10883_ net521 _06483_ vssd1 vssd1 vccd1 vccd1 _06484_ sky130_fd_sc_hd__and2_1
XFILLER_43_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15410_ net1744 _01620_ net1103 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[210\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_104_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12622_ _03125_ top.I2C.I2C_state\[1\] net3212 vssd1 vssd1 vccd1 vccd1 _00031_ sky130_fd_sc_hd__a21o_1
X_16390_ clknet_leaf_87_clk _07456_ net1264 vssd1 vssd1 vccd1 vccd1 top.SPI.register\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08618__A1 _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13611__A1 top.CPU.alu.program_counter\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11622__A0 _06373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15341_ net1675 _01551_ net1064 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[141\]
+ sky130_fd_sc_hd__dfrtp_1
X_12553_ net1346 top.SPI.busy top.CPU.done vssd1 vssd1 vccd1 vccd1 top.CPU.busy sky130_fd_sc_hd__or3b_1
XFILLER_156_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11504_ net3765 net256 _06730_ net489 vssd1 vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__a22o_1
XFILLER_145_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15272_ net1606 _01482_ net1066 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[72\]
+ sky130_fd_sc_hd__dfrtp_1
X_12484_ _06974_ _06991_ _06975_ vssd1 vssd1 vccd1 vccd1 _06993_ sky130_fd_sc_hd__or3b_1
XFILLER_138_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10189__A0 _03476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11435_ _05847_ net3661 net266 vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__mux2_1
XFILLER_7_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11366_ _06474_ net283 net274 net3526 vssd1 vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__a22o_1
X_13105_ top.SPI.count\[2\] _02716_ _02717_ _07426_ _06946_ vssd1 vssd1 vccd1 vccd1
+ _01276_ sky130_fd_sc_hd__o221a_1
X_10317_ net397 _05835_ _05948_ net404 vssd1 vssd1 vccd1 vccd1 _05949_ sky130_fd_sc_hd__o211a_1
XANTENNA__15601__RESET_B net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11548__C net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11297_ net3893 net292 _06706_ net494 vssd1 vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__a22o_1
XANTENNA__12006__A net1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10248_ net447 _05850_ _05881_ vssd1 vssd1 vccd1 vccd1 _05882_ sky130_fd_sc_hd__and3_1
X_13036_ net2742 _07443_ net896 vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__mux2_1
XANTENNA__11689__B1 net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1130 net1136 vssd1 vssd1 vccd1 vccd1 net1130 sky130_fd_sc_hd__clkbuf_4
Xfanout1141 net1143 vssd1 vssd1 vccd1 vccd1 net1141 sky130_fd_sc_hd__clkbuf_4
XFILLER_26_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14070__240 clknet_leaf_179_clk vssd1 vssd1 vccd1 vccd1 net1709 sky130_fd_sc_hd__inv_2
XFILLER_121_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09751__C1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1152 net1153 vssd1 vssd1 vccd1 vccd1 net1152 sky130_fd_sc_hd__clkbuf_4
X_10179_ net382 _05708_ _05709_ vssd1 vssd1 vccd1 vccd1 _05815_ sky130_fd_sc_hd__or3_1
XFILLER_93_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1163 net1164 vssd1 vssd1 vccd1 vccd1 net1163 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13763__C net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10361__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14367__537 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 net2006 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_163_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1174 net1179 vssd1 vssd1 vccd1 vccd1 net1174 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10900__A2 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1185 net1187 vssd1 vssd1 vccd1 vccd1 net1185 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14929__Q top.CPU.alu.program_counter\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09315__A top.CPU.control_unit.instruction\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1196 net1205 vssd1 vssd1 vccd1 vccd1 net1196 sky130_fd_sc_hd__clkbuf_2
X_14987_ clknet_leaf_93_clk _01232_ net1267 vssd1 vssd1 vccd1 vccd1 top.SPI.paroutput\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08306__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09503__C1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11283__C net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08857__A1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14111__281 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 net1750 sky130_fd_sc_hd__inv_2
XFILLER_19_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14408__578 clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 net2047 sky130_fd_sc_hd__inv_2
XFILLER_62_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_141_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11861__B1 net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08952__S1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15608_ net1942 _01818_ net1150 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[408\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08609__A1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09806__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12395__B net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10908__B _06472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15539_ net1873 _01749_ net1177 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[339\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11613__B1 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07817__C1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09060_ top.CPU.registers.data_out_r2_prev\[8\] net689 vssd1 vssd1 vccd1 vccd1 _04699_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__08490__C1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08011_ _03648_ _03649_ vssd1 vssd1 vccd1 vccd1 _03650_ sky130_fd_sc_hd__nand2b_4
XFILLER_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold602 top.SPI.parameters\[13\] vssd1 vssd1 vccd1 vccd1 net3159 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09196__S net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold613 top.CPU.registers.data\[319\] vssd1 vssd1 vccd1 vccd1 net3170 sky130_fd_sc_hd__dlygate4sd3_1
Xhold624 top.CPU.registers.data\[379\] vssd1 vssd1 vccd1 vccd1 net3181 sky130_fd_sc_hd__dlygate4sd3_1
Xhold635 top.CPU.registers.data\[362\] vssd1 vssd1 vccd1 vccd1 net3192 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08242__C1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold646 top.CPU.registers.data\[737\] vssd1 vssd1 vccd1 vccd1 net3203 sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 top.CPU.registers.data\[610\] vssd1 vssd1 vccd1 vccd1 net3214 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11392__A2 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12561__D _06251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold668 top.CPU.registers.data\[283\] vssd1 vssd1 vccd1 vccd1 net3225 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09962_ _05436_ _05503_ vssd1 vssd1 vccd1 vccd1 _05601_ sky130_fd_sc_hd__nand2_1
Xhold679 top.CPU.registers.data\[220\] vssd1 vssd1 vccd1 vccd1 net3236 sky130_fd_sc_hd__dlygate4sd3_1
X_13975__145 clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 net1614 sky130_fd_sc_hd__inv_2
X_08913_ top.CPU.registers.data\[426\] top.CPU.registers.data\[394\] net809 vssd1
+ vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__mux2_1
XANTENNA__09337__A2 net1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09893_ _04634_ _04661_ _04662_ _05279_ _05531_ vssd1 vssd1 vccd1 vccd1 _05532_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_51_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11144__A2 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13446__S net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout296_A _06662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08545__B1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1302 top.mmio.mem_data_i\[22\] vssd1 vssd1 vccd1 vccd1 net3859 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09742__C1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1313 top.I2C.data_out\[1\] vssd1 vssd1 vccd1 vccd1 net3870 sky130_fd_sc_hd__dlygate4sd3_1
X_08844_ net617 _04482_ _04477_ _03342_ vssd1 vssd1 vccd1 vccd1 _04483_ sky130_fd_sc_hd__o211a_1
XFILLER_84_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10352__B1 _05762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1324 top.CPU.registers.data\[998\] vssd1 vssd1 vccd1 vccd1 net3881 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1335 top.I2C.output_state\[24\] vssd1 vssd1 vccd1 vccd1 net3892 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1346 top.I2C.data_out\[11\] vssd1 vssd1 vccd1 vccd1 net3903 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1357 top.CPU.registers.data\[602\] vssd1 vssd1 vccd1 vccd1 net3914 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1368 top.mmio.mem_data_i\[12\] vssd1 vssd1 vccd1 vccd1 net3925 sky130_fd_sc_hd__dlygate4sd3_1
X_08775_ top.CPU.registers.data\[428\] top.CPU.registers.data\[396\] net814 vssd1
+ vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout463_A _03194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1379 top.I2C.output_state\[3\] vssd1 vssd1 vccd1 vccd1 net3936 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07726_ net681 _03346_ net947 _03345_ vssd1 vssd1 vccd1 vccd1 _03365_ sky130_fd_sc_hd__a211o_1
XFILLER_25_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07657_ top.CPU.control_unit.instruction\[4\] _03295_ _03293_ _03289_ net1038 vssd1
+ vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_0_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11852__B1 net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout251_X net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1372_A net1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout349_X net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout728_A net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07588_ top.CPU.registers.data\[319\] net836 net731 _03226_ vssd1 vssd1 vccd1 vccd1
+ _03227_ sky130_fd_sc_hd__o211a_1
XANTENNA__10377__Y _06007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09327_ top.CPU.registers.data\[548\] top.CPU.registers.data\[516\] net829 vssd1
+ vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__mux2_1
XANTENNA__07808__C1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout516_X net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09258_ top.CPU.registers.data\[453\] net1286 net1004 top.CPU.registers.data\[485\]
+ net900 vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__a221o_1
XFILLER_166_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07823__A2 net1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08209_ top.CPU.registers.data\[279\] net986 _03847_ vssd1 vssd1 vccd1 vccd1 _03848_
+ sky130_fd_sc_hd__a21o_1
X_09189_ top.CPU.registers.data_out_r1_prev\[6\] net871 _04813_ _04827_ vssd1 vssd1
+ vccd1 vccd1 _04828_ sky130_fd_sc_hd__o211a_2
XFILLER_119_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11220_ net460 net526 _06528_ vssd1 vssd1 vccd1 vccd1 _06665_ sky130_fd_sc_hd__and3_1
XANTENNA__08304__A net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout885_X net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_1035 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11383__A2 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11151_ net518 _06392_ vssd1 vssd1 vccd1 vccd1 _06635_ sky130_fd_sc_hd__nor2_1
XFILLER_150_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10102_ net404 _05739_ vssd1 vssd1 vccd1 vccd1 _05740_ sky130_fd_sc_hd__nand2_1
X_14054__224 clknet_leaf_122_clk vssd1 vssd1 vccd1 vccd1 net1693 sky130_fd_sc_hd__inv_2
XFILLER_150_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09328__A2 net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11082_ net3866 net366 _06595_ net324 vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__a22o_1
XFILLER_1_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11135__A2 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10033_ _03311_ _03322_ _03319_ vssd1 vssd1 vccd1 vccd1 _05672_ sky130_fd_sc_hd__a21o_4
XANTENNA__09733__C1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12260__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15890_ net2224 _02100_ net1105 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[690\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08000__A2 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12883__A2 _03823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input24_A DAT_I[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10159__A1_N _03477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10894__B2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_106_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11984_ _06544_ net345 net181 net2838 vssd1 vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_123_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16511_ clknet_leaf_59_clk _02673_ net1143 vssd1 vssd1 vccd1 vccd1 top.mmio.mem_data_i\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_86_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13723_ net3884 _03066_ _03069_ _07113_ vssd1 vssd1 vccd1 vccd1 _02630_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_123_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10935_ net490 net466 _06514_ net222 net3712 vssd1 vssd1 vccd1 vccd1 _02374_ sky130_fd_sc_hd__a32o_1
XANTENNA__11843__B1 net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12496__A _05154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08693__B net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11604__S net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16442_ clknet_leaf_67_clk _02605_ net1241 vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__dfrtp_1
X_13654_ net2841 _07347_ net665 vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__mux2_1
X_10866_ _05692_ _05693_ _06471_ vssd1 vssd1 vccd1 vccd1 _06473_ sky130_fd_sc_hd__and3_2
XFILLER_13_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12605_ top.SPI.timem\[16\] top.SPI.timem\[19\] top.SPI.timem\[18\] top.SPI.timem\[17\]
+ vssd1 vssd1 vccd1 vccd1 _07105_ sky130_fd_sc_hd__or4b_1
X_16373_ clknet_leaf_31_clk _02582_ net1126 vssd1 vssd1 vccd1 vccd1 top.CPU.fetch.current_ra\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13585_ net3977 _03017_ net580 vssd1 vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__mux2_1
XFILLER_13_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10797_ _05553_ _06402_ vssd1 vssd1 vccd1 vccd1 _06408_ sky130_fd_sc_hd__xor2_1
X_14752__922 clknet_leaf_125_clk vssd1 vssd1 vccd1 vccd1 net2391 sky130_fd_sc_hd__inv_2
XFILLER_157_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15324_ net1658 _01534_ net1195 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[124\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_158_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12536_ _04862_ _05543_ _07043_ _07044_ vssd1 vssd1 vccd1 vccd1 _07045_ sky130_fd_sc_hd__and4_1
XFILLER_12_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08913__S net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15255_ net1589 _01465_ net1184 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09016__A1 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12467_ _03819_ _03854_ _03887_ _03915_ vssd1 vssd1 vccd1 vccd1 _06976_ sky130_fd_sc_hd__a22o_1
XFILLER_126_831 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_144_Right_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11418_ _06554_ net275 net267 net3114 vssd1 vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__a22o_1
XANTENNA__08224__C1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13959__129 clknet_leaf_183_clk vssd1 vssd1 vccd1 vccd1 net1598 sky130_fd_sc_hd__inv_2
X_15186_ net1523 _01396_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r1_prev\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_12398_ _03122_ top.I2C.I2C_state\[12\] net2594 vssd1 vssd1 vccd1 vccd1 _00029_ sky130_fd_sc_hd__a21o_1
XANTENNA__08214__A net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11349_ net3826 net285 net275 _06214_ vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__a22o_1
XFILLER_4_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_165_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09744__S net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12323__A1 _04122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13520__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13266__S _02782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13019_ top.SPI.parameters\[11\] top.SPI.paroutput\[3\] net1356 vssd1 vssd1 vccd1
+ vccd1 _07435_ sky130_fd_sc_hd__mux2_1
XANTENNA__11677__A3 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07750__A1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12087__B1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08560_ top.CPU.registers.data\[143\] net811 net716 _04197_ vssd1 vssd1 vccd1 vccd1
+ _04199_ sky130_fd_sc_hd__a211o_1
XFILLER_81_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07511_ net1278 _03149_ vssd1 vssd1 vccd1 vccd1 _03150_ sky130_fd_sc_hd__nor2_1
XANTENNA__11834__B1 net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08491_ top.CPU.registers.data\[176\] top.CPU.registers.data\[144\] net820 vssd1
+ vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__mux2_1
XFILLER_81_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10919__A net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08058__A2 net1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09112_ net697 _04749_ _04750_ vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__and3_1
X_14495__665 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 net2134 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_44_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08463__C1 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11601__A3 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12853__B _03756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09043_ top.CPU.registers.data\[168\] top.CPU.registers.data\[136\] net808 vssd1
+ vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__mux2_1
XFILLER_136_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10654__A net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout211_A _06753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout309_A net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_111_Right_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09558__A2 net1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold410 top.CPU.registers.data\[812\] vssd1 vssd1 vccd1 vccd1 net2967 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_6_0_clk_X clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold421 top.CPU.registers.data\[177\] vssd1 vssd1 vccd1 vccd1 net2978 sky130_fd_sc_hd__dlygate4sd3_1
X_14038__208 clknet_leaf_178_clk vssd1 vssd1 vccd1 vccd1 net1677 sky130_fd_sc_hd__inv_2
Xhold432 top.CPU.registers.data\[807\] vssd1 vssd1 vccd1 vccd1 net2989 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10022__C1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11365__A2 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold443 top.CPU.registers.data\[846\] vssd1 vssd1 vccd1 vccd1 net3000 sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 top.CPU.registers.data\[970\] vssd1 vssd1 vccd1 vccd1 net3011 sky130_fd_sc_hd__dlygate4sd3_1
Xhold465 top.CPU.fetch.current_ra\[25\] vssd1 vssd1 vccd1 vccd1 net3022 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13905__75 clknet_leaf_180_clk vssd1 vssd1 vccd1 vccd1 net1544 sky130_fd_sc_hd__inv_2
Xhold476 top.CPU.registers.data\[697\] vssd1 vssd1 vccd1 vccd1 net3033 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1218_A net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold487 top.CPU.registers.data\[462\] vssd1 vssd1 vccd1 vccd1 net3044 sky130_fd_sc_hd__dlygate4sd3_1
Xhold498 top.CPU.registers.data\[403\] vssd1 vssd1 vccd1 vccd1 net3055 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout901 net910 vssd1 vssd1 vccd1 vccd1 net901 sky130_fd_sc_hd__buf_4
XANTENNA__13684__B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09945_ _04094_ _04124_ vssd1 vssd1 vccd1 vccd1 _05584_ sky130_fd_sc_hd__nor2_1
Xfanout912 net914 vssd1 vssd1 vccd1 vccd1 net912 sky130_fd_sc_hd__buf_2
Xfanout923 net924 vssd1 vssd1 vccd1 vccd1 net923 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12314__A1 _05498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11117__A2 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout934 net935 vssd1 vssd1 vccd1 vccd1 net934 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout299_X net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout678_A net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout945 net946 vssd1 vssd1 vccd1 vccd1 net945 sky130_fd_sc_hd__clkbuf_4
Xfanout956 net962 vssd1 vssd1 vccd1 vccd1 net956 sky130_fd_sc_hd__clkbuf_4
X_09876_ _03442_ _05514_ _03374_ vssd1 vssd1 vccd1 vccd1 _05515_ sky130_fd_sc_hd__a21oi_1
Xfanout967 net970 vssd1 vssd1 vccd1 vccd1 net967 sky130_fd_sc_hd__clkbuf_4
XFILLER_161_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1110 _01247_ vssd1 vssd1 vccd1 vccd1 net3667 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout978 net985 vssd1 vssd1 vccd1 vccd1 net978 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1006_X net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1121 top.CPU.registers.data\[224\] vssd1 vssd1 vccd1 vccd1 net3678 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout989 net994 vssd1 vssd1 vccd1 vccd1 net989 sky130_fd_sc_hd__clkbuf_4
Xhold1132 top.CPU.registers.data\[899\] vssd1 vssd1 vccd1 vccd1 net3689 sky130_fd_sc_hd__dlygate4sd3_1
X_08827_ _04465_ vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__inv_2
XANTENNA__09730__A2 net1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1143 top.mmio.mem_data_i\[0\] vssd1 vssd1 vccd1 vccd1 net3700 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1154 top.CPU.registers.data\[745\] vssd1 vssd1 vccd1 vccd1 net3711 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout466_X net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout845_A net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1165 top.CPU.registers.data\[1017\] vssd1 vssd1 vccd1 vccd1 net3722 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1176 top.CPU.registers.data\[672\] vssd1 vssd1 vccd1 vccd1 net3733 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_173_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1187 top.CPU.registers.data\[344\] vssd1 vssd1 vccd1 vccd1 net3744 sky130_fd_sc_hd__dlygate4sd3_1
X_08758_ _04394_ _04395_ vssd1 vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_68_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1198 top.mmio.mem_data_i\[28\] vssd1 vssd1 vccd1 vccd1 net3755 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10628__A1 _05672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11825__B1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07709_ top.CPU.registers.data\[383\] net1307 net1030 top.CPU.registers.data\[351\]
+ net681 vssd1 vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__o221a_1
X_08689_ _04294_ _04326_ vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout633_X net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09494__A1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1375_X net1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10720_ net552 _06333_ vssd1 vssd1 vccd1 vccd1 _06335_ sky130_fd_sc_hd__or2_1
XFILLER_159_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14736__906 clknet_leaf_199_clk vssd1 vssd1 vccd1 vccd1 net2375 sky130_fd_sc_hd__inv_2
XFILLER_110_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10651_ top.CPU.fetch.current_ra\[10\] net1042 net881 top.CPU.handler.toreg\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06269_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout800_X net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10582_ _06202_ vssd1 vssd1 vccd1 vccd1 _06203_ sky130_fd_sc_hd__inv_2
X_13370_ top.mmio.mem_data_i\[17\] _07089_ net555 top.I2C.data_out\[17\] vssd1 vssd1
+ vccd1 vccd1 _02896_ sky130_fd_sc_hd__a22o_1
XFILLER_155_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08733__S net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12321_ net2578 _03984_ net1187 vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__mux2_1
XANTENNA__12255__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15040_ clknet_leaf_91_clk _01285_ net1269 vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_181_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12002__B1 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12252_ net2954 net132 net432 vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__mux2_1
XANTENNA__10283__B net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11356__A2 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11203_ net3599 net297 _06658_ net482 vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__a22o_1
XFILLER_135_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12183_ top.CPU.registers.data\[59\] net170 vssd1 vssd1 vccd1 vccd1 _06858_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_147_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_61_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11134_ net471 _06624_ vssd1 vssd1 vccd1 vccd1 _06626_ sky130_fd_sc_hd__nor2_1
XFILLER_150_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12305__A1 _05054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08509__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_196_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09706__C1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11065_ net3363 net366 _06589_ net323 vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__a22o_1
X_15942_ net2276 _02152_ net1072 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[742\]
+ sky130_fd_sc_hd__dfrtp_1
X_10016_ net417 net374 vssd1 vssd1 vccd1 vccd1 _05655_ sky130_fd_sc_hd__nand2_1
XANTENNA__09182__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_76_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10867__A1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15873_ net2207 _02083_ net1231 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[673\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07732__A1 top.CPU.alu.immediate\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12003__B net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08908__S net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11816__B1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11967_ _06516_ net347 net231 net3186 vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__a22o_1
XANTENNA__08288__A2 net1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13706_ top.SPI.timem\[5\] top.SPI.timem\[6\] _03056_ vssd1 vssd1 vccd1 vccd1 _03058_
+ sky130_fd_sc_hd__and3_1
XFILLER_72_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10918_ net478 net456 _06504_ net220 net3090 vssd1 vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__a32o_1
X_14182__352 clknet_leaf_125_clk vssd1 vssd1 vccd1 vccd1 net1821 sky130_fd_sc_hd__inv_2
X_11898_ _03174_ net570 _06751_ vssd1 vssd1 vccd1 vccd1 _06769_ sky130_fd_sc_hd__or3_1
X_14479__649 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 net2118 sky130_fd_sc_hd__inv_2
X_16425_ clknet_leaf_55_clk _00007_ net1141 vssd1 vssd1 vccd1 vccd1 top.I2C.I2C_state\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_134_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13637_ net3264 _07189_ net664 vssd1 vssd1 vccd1 vccd1 _02571_ sky130_fd_sc_hd__mux2_1
X_10849_ net382 _06414_ vssd1 vssd1 vccd1 vccd1 _06457_ sky130_fd_sc_hd__nand2_1
XFILLER_13_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08445__C1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_14_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16356_ clknet_leaf_28_clk _02565_ net1149 vssd1 vssd1 vccd1 vccd1 top.CPU.fetch.current_ra\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13568_ net1350 _06309_ vssd1 vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__nand2_1
X_14223__393 clknet_leaf_178_clk vssd1 vssd1 vccd1 vccd1 net1862 sky130_fd_sc_hd__inv_2
XANTENNA__07799__A1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14879__1049 clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 net2518 sky130_fd_sc_hd__inv_2
XANTENNA__14942__Q top.CPU.alu.program_counter\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12792__A1 top.CPU.alu.program_counter\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15307_ net1641 _01517_ net1058 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[107\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_118_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12519_ _06977_ _06981_ _06982_ vssd1 vssd1 vccd1 vccd1 _07028_ sky130_fd_sc_hd__or3_1
X_16287_ clknet_leaf_62_clk _02497_ net1161 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.toreg\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13499_ top.CPU.data_out\[8\] net588 _02968_ _02969_ vssd1 vssd1 vccd1 vccd1 _02506_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08460__A2 net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_149_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15238_ net1572 _01448_ net1081 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_160_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11347__A2 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_29_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08748__B1 top.CPU.control_unit.instruction\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10555__A0 _04225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15169_ net1506 _01379_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r1_prev\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08843__S0 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout208 net210 vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__clkbuf_4
Xfanout219 _06525_ vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__clkbuf_8
XFILLER_140_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07991_ top.CPU.registers.data\[856\] net1289 net1009 top.CPU.registers.data\[888\]
+ net932 vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__a221o_1
XANTENNA__10921__B net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_7_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_7_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07971__A1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09730_ top.CPU.registers.data\[603\] net1331 net859 top.CPU.registers.data\[635\]
+ net777 vssd1 vssd1 vccd1 vccd1 _05369_ sky130_fd_sc_hd__a221o_1
XFILLER_101_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10413__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09661_ _04060_ _05299_ _03650_ vssd1 vssd1 vccd1 vccd1 _05300_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_2_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08612_ net1284 _04249_ _04250_ vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__or3_1
X_09592_ top.CPU.control_unit.instruction\[7\] _03152_ _05228_ _05230_ vssd1 vssd1
+ vccd1 vccd1 _05231_ sky130_fd_sc_hd__a22o_1
XANTENNA__11807__B1 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08543_ net935 _04179_ _04181_ net953 vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__o211a_1
XFILLER_70_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout161_A _06760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout259_A net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08474_ net678 _04106_ _04107_ _04112_ vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__a31o_1
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1070_A net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout426_A _06756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1168_A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11586__A2 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08451__A2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout214_X net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1335_A net1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09026_ _04634_ _04663_ vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__nor2_1
XANTENNA__11199__B _06270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout795_A net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11338__A2 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1443_A top.SPI.busy vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09892__B _04698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold240 top.CPU.registers.data\[400\] vssd1 vssd1 vccd1 vccd1 net2797 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10546__B1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08203__A2 net1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold251 top.CPU.registers.data\[913\] vssd1 vssd1 vccd1 vccd1 net2808 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 top.CPU.registers.data\[553\] vssd1 vssd1 vccd1 vccd1 net2819 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 top.SPI.parameters\[25\] vssd1 vssd1 vccd1 vccd1 net2830 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09384__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold284 top.CPU.fetch.current_ra\[26\] vssd1 vssd1 vccd1 vccd1 net2841 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_120_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold295 top.CPU.registers.data\[292\] vssd1 vssd1 vccd1 vccd1 net2852 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout583_X net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout962_A net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout720 net722 vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout731 net734 vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__clkbuf_4
X_09928_ _05564_ _05566_ _05536_ vssd1 vssd1 vccd1 vccd1 _05567_ sky130_fd_sc_hd__a21oi_1
Xfanout742 net746 vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__clkbuf_4
Xfanout753 net760 vssd1 vssd1 vccd1 vccd1 net753 sky130_fd_sc_hd__buf_2
XFILLER_172_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout764 net772 vssd1 vssd1 vccd1 vccd1 net764 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_142_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09164__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout775 net777 vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__clkbuf_4
Xfanout786 net794 vssd1 vssd1 vccd1 vccd1 net786 sky130_fd_sc_hd__buf_2
XANTENNA__09703__A2 net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09859_ _05482_ _05497_ vssd1 vssd1 vccd1 vccd1 _05498_ sky130_fd_sc_hd__or2_4
Xfanout797 net799 vssd1 vssd1 vccd1 vccd1 net797 sky130_fd_sc_hd__clkbuf_4
XFILLER_100_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout848_X net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13634__S net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12870_ top.CPU.alu.program_counter\[23\] _03823_ vssd1 vssd1 vccd1 vccd1 _07317_
+ sky130_fd_sc_hd__or2_1
XFILLER_27_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13799__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11821_ net144 net3674 net156 vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__mux2_1
X_14166__336 clknet_leaf_180_clk vssd1 vssd1 vccd1 vccd1 net1805 sky130_fd_sc_hd__inv_2
XANTENNA__11662__B net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11274__B2 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11752_ _06591_ net199 net192 net3052 vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__a22o_1
XFILLER_26_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10703_ _05632_ _05753_ vssd1 vssd1 vccd1 vccd1 _06318_ sky130_fd_sc_hd__nand2_1
XFILLER_14_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14207__377 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 net1846 sky130_fd_sc_hd__inv_2
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11683_ net463 _06504_ net234 net164 net3217 vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__a32o_1
XFILLER_81_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16210_ net2544 _02420_ net1081 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[1010\]
+ sky130_fd_sc_hd__dfrtp_1
X_13422_ top.I2C.data_out\[31\] net556 _02933_ _07088_ vssd1 vssd1 vccd1 vccd1 _02934_
+ sky130_fd_sc_hd__a22o_1
XFILLER_41_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07868__A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10634_ top.CPU.fetch.current_ra\[11\] net1040 net633 top.CPU.handler.toreg\[11\]
+ _06252_ vssd1 vssd1 vccd1 vccd1 _06253_ sky130_fd_sc_hd__a221o_4
XANTENNA__08427__C1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12223__B1 _03185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16141_ net2475 _02351_ net1076 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[941\]
+ sky130_fd_sc_hd__dfrtp_1
X_13353_ net889 _02883_ vssd1 vssd1 vccd1 vccd1 _02884_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_118_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07587__B net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10565_ _04325_ net507 _06183_ _06186_ vssd1 vssd1 vccd1 vccd1 _06187_ sky130_fd_sc_hd__a211o_1
XFILLER_10_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12304_ net2596 _04986_ net1198 vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__mux2_1
XFILLER_155_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16072_ net2406 _02282_ net1098 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[872\]
+ sky130_fd_sc_hd__dfrtp_1
X_13284_ _03127_ net3467 net895 vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__a21o_1
X_10496_ _05741_ _06120_ _06119_ vssd1 vssd1 vccd1 vccd1 _06121_ sky130_fd_sc_hd__a21oi_1
XFILLER_6_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15023_ clknet_leaf_83_clk _01268_ net1261 vssd1 vssd1 vccd1 vccd1 top.SPI.parameters\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_136_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12235_ top.CPU.registers.data\[33\] net655 _03185_ vssd1 vssd1 vccd1 vccd1 _06884_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__12940__C top.CPU.alu.program_counter\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12166_ top.CPU.registers.data\[69\] net645 net360 vssd1 vssd1 vccd1 vccd1 _06851_
+ sky130_fd_sc_hd__o21a_1
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10741__B _06354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07953__A1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11117_ net3864 net302 _06616_ net313 vssd1 vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__a22o_1
X_13896__66 clknet_leaf_125_clk vssd1 vssd1 vccd1 vccd1 net1535 sky130_fd_sc_hd__inv_2
XANTENNA__09155__A0 _04792_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12097_ _06631_ _06770_ _06816_ net176 net3769 vssd1 vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__a32o_1
XFILLER_77_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11048_ net325 net133 net538 net368 net2970 vssd1 vssd1 vccd1 vccd1 _02329_ sky130_fd_sc_hd__a32o_1
X_15925_ net2259 _02135_ net1210 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[725\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12949__A top.CPU.alu.program_counter\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput8 DAT_I[15] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11501__A2 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08902__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15856_ net2190 _02066_ net1154 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[656\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12668__B top.CPU.alu.program_counter\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15787_ net2121 _01997_ net1058 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[587\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_91_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12999_ _07426_ vssd1 vssd1 vccd1 vccd1 _07427_ sky130_fd_sc_hd__inv_2
XANTENNA__11291__C net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11265__B2 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08666__C1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08130__A1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11804__A3 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13006__A2 _07429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16408_ clknet_leaf_56_clk net3658 net1145 vssd1 vssd1 vccd1 vccd1 top.I2C.I2C_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_08190_ top.CPU.registers.data\[247\] net1381 net987 top.CPU.registers.data\[215\]
+ net911 vssd1 vssd1 vccd1 vccd1 _03829_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_41_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08373__S net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08969__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16339_ clknet_leaf_69_clk _02548_ net1167 vssd1 vssd1 vccd1 vccd1 top.CPU.addressnew\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10776__B1 _06383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1027 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_778 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12517__A1 _04155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_144_Left_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10932__A net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10528__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08197__A1 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11740__A2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07974_ net1033 _03610_ _03612_ vssd1 vssd1 vccd1 vccd1 _03613_ sky130_fd_sc_hd__a21oi_4
XFILLER_102_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09713_ net960 _05351_ _05348_ net614 vssd1 vssd1 vccd1 vccd1 _05352_ sky130_fd_sc_hd__a211o_1
XANTENNA__12859__A top.CPU.alu.program_counter\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13454__S net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09644_ _04533_ _04534_ vssd1 vssd1 vccd1 vccd1 _05283_ sky130_fd_sc_hd__or2_2
XFILLER_67_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_153_Left_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09575_ top.CPU.registers.data\[160\] top.CPU.registers.data\[128\] net973 vssd1
+ vssd1 vccd1 vccd1 _05214_ sky130_fd_sc_hd__mux2_1
XFILLER_55_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout164_X net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout543_A net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08526_ top.CPU.registers.data\[976\] net1290 net1011 top.CPU.registers.data\[1008\]
+ net907 vssd1 vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__a221o_1
XANTENNA__12453__B1 _03241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08121__A1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout710_A net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08457_ top.CPU.registers.data\[401\] net1296 net1016 top.CPU.registers.data\[433\]
+ net913 vssd1 vssd1 vccd1 vccd1 _04096_ sky130_fd_sc_hd__a221o_1
XANTENNA__08672__A2 net1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout429_X net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout808_A net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11008__B2 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12205__B1 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07880__B1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08388_ net619 _04022_ _04026_ net604 vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__a211o_1
XFILLER_149_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11559__A2 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09621__A1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09082__C1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_162_Left_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1338_X net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14551__721 clknet_leaf_76_clk vssd1 vssd1 vccd1 vccd1 net2190 sky130_fd_sc_hd__inv_2
X_10350_ net412 _05752_ vssd1 vssd1 vccd1 vccd1 _05981_ sky130_fd_sc_hd__nor2_1
XANTENNA__12508__A1 _04222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout798_X net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13629__S net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12508__B2 _04324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09009_ top.CPU.registers.data\[329\] net1369 net964 top.CPU.registers.data\[361\]
+ net1280 vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__o221a_1
X_10281_ net402 _05913_ vssd1 vssd1 vccd1 vccd1 _05914_ sky130_fd_sc_hd__nand2_1
XFILLER_117_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12020_ net133 net3436 net151 vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_76_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11192__A0 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout965_X net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16302__Q top.CPU.data_out\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11731__A2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout550 _03316_ vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__clkbuf_4
Xfanout561 _06933_ vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__buf_2
XFILLER_116_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout572 net575 vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__clkbuf_4
Xfanout583 _02994_ vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__clkbuf_4
XFILLER_47_913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09688__A1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_171_Left_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15710_ net2044 _01920_ net1238 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[510\]
+ sky130_fd_sc_hd__dfrtp_1
X_12922_ top.CPU.alu.program_counter\[27\] _07364_ net1361 vssd1 vssd1 vccd1 vccd1
+ _01190_ sky130_fd_sc_hd__mux2_1
XANTENNA__11495__A1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14878__1048 clknet_leaf_152_clk vssd1 vssd1 vccd1 vccd1 net2517 sky130_fd_sc_hd__inv_2
XFILLER_76_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08458__S net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15641_ net1975 _01851_ net1246 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[441\]
+ sky130_fd_sc_hd__dfrtp_1
X_12853_ top.CPU.alu.program_counter\[21\] _03756_ vssd1 vssd1 vccd1 vccd1 _07302_
+ sky130_fd_sc_hd__xor2_1
X_11804_ _06483_ _06648_ net241 net157 net3008 vssd1 vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__a32o_1
XANTENNA__11247__A1 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15572_ net1906 _01782_ net1073 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[372\]
+ sky130_fd_sc_hd__dfrtp_1
X_12784_ top.CPU.alu.program_counter\[14\] _07228_ vssd1 vssd1 vccd1 vccd1 _07240_
+ sky130_fd_sc_hd__and2_1
X_11735_ _06581_ net209 net195 net2907 vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_155_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11612__S net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08046__X _03685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11666_ net468 _06476_ net240 net166 net2915 vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_172_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_14_0_clk_X clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13405_ top.CPU.control_unit.instruction\[26\] _02921_ net670 vssd1 vssd1 vccd1 vccd1
+ _02460_ sky130_fd_sc_hd__mux2_1
X_10617_ _04603_ _06235_ _05533_ vssd1 vssd1 vccd1 vccd1 _06236_ sky130_fd_sc_hd__a21o_1
XFILLER_128_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09073__C1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11597_ net137 net3153 net214 vssd1 vssd1 vccd1 vccd1 _01952_ sky130_fd_sc_hd__mux2_1
XFILLER_127_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_133_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16124_ net2458 _02334_ net1234 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[924\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10222__A2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13336_ top.mmio.mem_data_i\[8\] _07089_ net554 top.I2C.data_out\[8\] vssd1 vssd1
+ vccd1 vccd1 _02871_ sky130_fd_sc_hd__a22o_1
X_10548_ _06160_ _06168_ _06169_ _06170_ vssd1 vssd1 vccd1 vccd1 _06171_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_133_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14294__464 clknet_leaf_180_clk vssd1 vssd1 vccd1 vccd1 net1933 sky130_fd_sc_hd__inv_2
XFILLER_109_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16055_ net2389 _02265_ net1182 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[855\]
+ sky130_fd_sc_hd__dfrtp_1
X_13267_ net3931 _02814_ _02818_ net1053 vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__a22o_1
XFILLER_170_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10479_ top.CPU.fetch.current_ra\[18\] net1044 net882 top.CPU.handler.toreg\[18\]
+ _06104_ vssd1 vssd1 vccd1 vccd1 _06105_ sky130_fd_sc_hd__a221o_2
XANTENNA__08179__A1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15006_ clknet_leaf_94_clk _01251_ net1267 vssd1 vssd1 vccd1 vccd1 top.SPI.parameters\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_130_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12218_ top.CPU.registers.data\[42\] net647 net365 _06687_ net562 vssd1 vssd1 vccd1
+ vccd1 _06876_ sky130_fd_sc_hd__o2111a_1
XFILLER_151_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13198_ top.I2C.data_out\[17\] net892 _02774_ vssd1 vssd1 vccd1 vccd1 _02778_ sky130_fd_sc_hd__mux2_1
XFILLER_111_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07926__A1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11722__A2 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12149_ net3955 net172 _06842_ _06500_ vssd1 vssd1 vccd1 vccd1 _01488_ sky130_fd_sc_hd__a22o_1
XFILLER_97_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09128__B1 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13475__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12679__A net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07780__B net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15908_ net2242 _02118_ net1211 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[708\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11486__A1 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07690_ _03285_ _03298_ _03304_ _03310_ vssd1 vssd1 vccd1 vccd1 _03329_ sky130_fd_sc_hd__and4_1
XFILLER_38_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15839_ net2173 _02049_ net1224 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[639\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_18_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09360_ top.CPU.registers.data\[451\] net1297 net1018 top.CPU.registers.data\[483\]
+ net915 vssd1 vssd1 vccd1 vccd1 _04999_ sky130_fd_sc_hd__a221o_1
XFILLER_52_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08639__C1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08103__A1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10446__C1 _05742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08311_ top.CPU.registers.data\[819\] top.CPU.registers.data\[787\] net826 vssd1
+ vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__mux2_1
XFILLER_162_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09291_ top.CPU.registers.data\[4\] net992 vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__and2_1
XFILLER_61_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10927__A _05694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08242_ net753 _03879_ _03880_ net776 vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__o211a_1
XANTENNA_wire599_X net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07862__B1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14535__705 clknet_leaf_186_clk vssd1 vssd1 vccd1 vccd1 net2174 sky130_fd_sc_hd__inv_2
X_08173_ top.CPU.registers.data\[663\] net1325 net856 top.CPU.registers.data\[695\]
+ net723 vssd1 vssd1 vccd1 vccd1 _03812_ sky130_fd_sc_hd__a221o_1
XFILLER_146_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08406__A2 net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16614__A net1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1033_A net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09367__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout493_A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10381__B net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12493__A2_N _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11713__A2 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1200_A net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09515__X _05154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07957_ top.CPU.registers.data\[664\] net1321 net852 top.CPU.registers.data\[696\]
+ net706 vssd1 vssd1 vccd1 vccd1 _03596_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout281_X net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout660_A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout758_A net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout379_X net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08278__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11477__B2 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07888_ top.CPU.registers.data\[252\] net1394 net832 top.CPU.registers.data\[220\]
+ net778 vssd1 vssd1 vccd1 vccd1 _03527_ sky130_fd_sc_hd__a221o_1
XFILLER_83_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09627_ top.CPU.alu.program_counter\[0\] _05265_ net1034 vssd1 vssd1 vccd1 vccd1
+ _05266_ sky130_fd_sc_hd__mux2_2
XANTENNA_fanout546_X net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout925_A _03353_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09558_ top.CPU.registers.data\[736\] net1377 net973 top.CPU.registers.data\[704\]
+ net902 vssd1 vssd1 vccd1 vccd1 _05197_ sky130_fd_sc_hd__a221o_1
XANTENNA__11229__B2 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09250__X _04889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08509_ top.CPU.registers.data\[784\] net820 net745 _04147_ vssd1 vssd1 vccd1 vccd1
+ _04148_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout713_X net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08645__A2 net1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09489_ top.CPU.registers.data\[161\] top.CPU.registers.data\[129\] net998 vssd1
+ vssd1 vccd1 vccd1 _05128_ sky130_fd_sc_hd__mux2_1
XANTENNA__09842__A1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11520_ net484 _05962_ net354 net250 net2940 vssd1 vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__a32o_1
XFILLER_168_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07853__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11451_ net141 net3447 net263 vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__mux2_1
X_14278__448 clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 net1917 sky130_fd_sc_hd__inv_2
XFILLER_11_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10402_ _06029_ _06030_ _06013_ _06028_ vssd1 vssd1 vccd1 vccd1 _06031_ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_150_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08802__C1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11382_ net473 _06501_ net272 net3246 vssd1 vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__a22o_1
XANTENNA__12771__B top.CPU.alu.program_counter\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09070__A2 net1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13121_ net2776 _02725_ net897 vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__mux2_1
XFILLER_125_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11952__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14022__192 clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 net1661 sky130_fd_sc_hd__inv_2
XFILLER_139_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10333_ _05290_ _05292_ _05297_ _04125_ vssd1 vssd1 vccd1 vccd1 _05964_ sky130_fd_sc_hd__a211oi_2
XFILLER_125_748 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12263__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14319__489 clknet_leaf_179_clk vssd1 vssd1 vccd1 vccd1 net1958 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_111_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09358__B1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13052_ net2896 _07451_ net895 vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__mux2_1
XANTENNA__09138__A net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10264_ net417 net385 net391 vssd1 vssd1 vccd1 vccd1 _05898_ sky130_fd_sc_hd__a21o_1
XFILLER_152_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12003_ net1402 net651 net538 net362 vssd1 vssd1 vccd1 vccd1 _06778_ sky130_fd_sc_hd__and4b_1
XANTENNA__11704__A2 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1301 _03113_ vssd1 vssd1 vccd1 vccd1 net1301 sky130_fd_sc_hd__clkbuf_4
X_10195_ _03576_ net507 net510 _03578_ vssd1 vssd1 vccd1 vccd1 _05831_ sky130_fd_sc_hd__o2bb2a_1
Xfanout1312 net1323 vssd1 vssd1 vccd1 vccd1 net1312 sky130_fd_sc_hd__clkbuf_2
Xfanout1323 _03109_ vssd1 vssd1 vccd1 vccd1 net1323 sky130_fd_sc_hd__buf_4
XFILLER_78_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1334 net1337 vssd1 vssd1 vccd1 vccd1 net1334 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09572__S net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08581__A1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1345 net67 vssd1 vssd1 vccd1 vccd1 net1345 sky130_fd_sc_hd__clkbuf_2
Xfanout1356 top.SPI.state\[2\] vssd1 vssd1 vccd1 vccd1 net1356 sky130_fd_sc_hd__buf_2
X_13866__36 clknet_leaf_149_clk vssd1 vssd1 vccd1 vccd1 net1505 sky130_fd_sc_hd__inv_2
XFILLER_38_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1367 net1368 vssd1 vssd1 vccd1 vccd1 net1367 sky130_fd_sc_hd__buf_2
XANTENNA__13457__A2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1378 net1379 vssd1 vssd1 vccd1 vccd1 net1378 sky130_fd_sc_hd__buf_4
Xfanout380 _05234_ vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__buf_2
XFILLER_94_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout391 net392 vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1389 net1395 vssd1 vssd1 vccd1 vccd1 net1389 sky130_fd_sc_hd__buf_4
XANTENNA__11607__S net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12905_ top.CPU.alu.program_counter\[26\] _05499_ vssd1 vssd1 vccd1 vccd1 _07349_
+ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_194_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_194_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12011__B _06781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12836_ top.CPU.alu.program_counter\[19\] top.CPU.alu.program_counter\[18\] _07270_
+ vssd1 vssd1 vccd1 vccd1 _07287_ sky130_fd_sc_hd__and3_1
X_15624_ net1958 _01834_ net1089 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[424\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08916__S net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_174_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07820__S net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14720__890 clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 net2359 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_174_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15555_ net1889 _01765_ net1207 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[355\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08097__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12767_ top.CPU.alu.program_counter\[13\] _04392_ vssd1 vssd1 vccd1 vccd1 _07224_
+ sky130_fd_sc_hd__and2_1
XANTENNA__09294__C1 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11718_ _06558_ net197 net420 net3035 vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__a22o_1
XANTENNA__07844__B1 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15486_ net1820 _01696_ net1237 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[286\]
+ sky130_fd_sc_hd__dfrtp_1
X_12698_ top.CPU.alu.program_counter\[6\] _07152_ vssd1 vssd1 vccd1 vccd1 _07162_
+ sky130_fd_sc_hd__xor2_1
Xinput11 DAT_I[18] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
XFILLER_128_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09046__C1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11649_ _06233_ net201 net424 net3750 vssd1 vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__a22o_1
Xinput22 DAT_I[28] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__buf_1
Xinput33 DAT_I[9] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09747__S net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12196__A2 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold806 top.CPU.registers.data\[909\] vssd1 vssd1 vccd1 vccd1 net3363 sky130_fd_sc_hd__dlygate4sd3_1
Xhold817 top.CPU.registers.data\[762\] vssd1 vssd1 vccd1 vccd1 net3374 sky130_fd_sc_hd__dlygate4sd3_1
X_16107_ net2441 _02317_ net1064 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[907\]
+ sky130_fd_sc_hd__dfrtp_1
X_13319_ top.CPU.control_unit.instruction\[3\] _02858_ net669 vssd1 vssd1 vccd1 vccd1
+ _02437_ sky130_fd_sc_hd__mux2_1
XANTENNA__11943__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold828 top.CPU.registers.data\[589\] vssd1 vssd1 vccd1 vccd1 net3385 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold839 top.CPU.registers.data\[523\] vssd1 vssd1 vccd1 vccd1 net3396 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13145__A1 top.CPU.data_out\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16038_ net2372 _02248_ net1075 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[838\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_36_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08860_ net688 _04497_ _04498_ vssd1 vssd1 vccd1 vccd1 _04499_ sky130_fd_sc_hd__a21o_1
XFILLER_111_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07811_ top.CPU.registers.data\[573\] top.CPU.registers.data\[541\] net817 vssd1
+ vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__mux2_1
X_08791_ net879 net450 _04429_ vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__o21ai_4
XFILLER_96_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07742_ net755 _03379_ _03380_ vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__o21ai_1
XFILLER_93_860 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12120__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07673_ _03285_ _03311_ _03308_ _03307_ vssd1 vssd1 vccd1 vccd1 _03312_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_185_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_185_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_19_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09412_ net751 _05049_ _05050_ net708 vssd1 vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__o211a_1
X_13880__50 clknet_leaf_166_clk vssd1 vssd1 vccd1 vccd1 net1519 sky130_fd_sc_hd__inv_2
XFILLER_53_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09343_ top.CPU.registers.data\[452\] net1329 net860 top.CPU.registers.data\[484\]
+ net726 vssd1 vssd1 vccd1 vccd1 _04982_ sky130_fd_sc_hd__a221o_1
XFILLER_34_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout241_A net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08627__A2 net1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09824__A1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_158_Right_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09274_ net672 _04896_ _04897_ vssd1 vssd1 vccd1 vccd1 _04913_ sky130_fd_sc_hd__and3_1
XANTENNA__07835__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08127__A net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10249__A2_N net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08225_ top.CPU.registers.data\[182\] top.CPU.registers.data\[150\] net835 vssd1
+ vssd1 vccd1 vccd1 _03864_ sky130_fd_sc_hd__mux2_1
XANTENNA__09037__C1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout127_X net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14006__176 clknet_leaf_182_clk vssd1 vssd1 vccd1 vccd1 net1645 sky130_fd_sc_hd__inv_2
XANTENNA__12187__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08156_ top.CPU.registers.data\[247\] net1391 net824 top.CPU.registers.data\[215\]
+ net773 vssd1 vssd1 vccd1 vccd1 _03795_ sky130_fd_sc_hd__a221o_1
XFILLER_146_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09052__A2 net1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14877__1047 clknet_leaf_134_clk vssd1 vssd1 vccd1 vccd1 net2516 sky130_fd_sc_hd__inv_2
XFILLER_162_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11395__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08260__B1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08087_ top.CPU.registers.data\[597\] net1330 net861 top.CPU.registers.data\[629\]
+ net776 vssd1 vssd1 vccd1 vccd1 _03726_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_56_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1036_X net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_73_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout496_X net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout875_A net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08797__A net1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09392__S net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14663__833 clknet_leaf_184_clk vssd1 vssd1 vccd1 vccd1 net2302 sky130_fd_sc_hd__inv_2
XANTENNA_fanout663_X net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08989_ net783 _04626_ _04627_ net713 vssd1 vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__o211a_1
XFILLER_102_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08315__A1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09512__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12111__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10658__C1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10951_ net520 net138 net545 vssd1 vssd1 vccd1 vccd1 _06526_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_176_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_176_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout928_X net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14704__874 clknet_leaf_196_clk vssd1 vssd1 vccd1 vccd1 net2343 sky130_fd_sc_hd__inv_2
XANTENNA__13642__S net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13670_ net2828 net331 _03048_ top.CPU.addressnew\[3\] vssd1 vssd1 vccd1 vccd1 _02598_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10673__A2 _06288_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10882_ _05693_ _05934_ _06471_ vssd1 vssd1 vccd1 vccd1 _06483_ sky130_fd_sc_hd__and3_1
XANTENNA__10838__Y _06447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12766__B _04392_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08079__A0 _03716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12621_ _07062_ _07081_ vssd1 vssd1 vccd1 vccd1 _00025_ sky130_fd_sc_hd__and2b_1
XANTENNA__13072__A0 top.CPU.data_out\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09276__C1 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12258__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_125_Right_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15340_ net1674 _01550_ net1077 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[140\]
+ sky130_fd_sc_hd__dfrtp_1
X_12552_ top.CPU.done top.CPU.handler.state\[0\] _07059_ vssd1 vssd1 vccd1 vccd1 _00022_
+ sky130_fd_sc_hd__a21o_1
XFILLER_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11503_ net466 _06636_ vssd1 vssd1 vccd1 vccd1 _06730_ sky130_fd_sc_hd__nor2_1
XFILLER_156_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15271_ net1605 _01481_ net1197 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[71\]
+ sky130_fd_sc_hd__dfrtp_1
X_12483_ _03819_ _03854_ vssd1 vssd1 vccd1 vccd1 _06992_ sky130_fd_sc_hd__or2_1
X_11434_ _05808_ net3836 net263 vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__mux2_1
XANTENNA__10189__A1 _03544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08471__S net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11386__B1 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11925__A2 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_100_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_100_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11365_ net490 net474 net520 _06473_ _06715_ vssd1 vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__a41o_1
X_13104_ top.SPI.count\[2\] top.SPI.count\[1\] top.SPI.count\[0\] vssd1 vssd1 vccd1
+ vccd1 _02717_ sky130_fd_sc_hd__nand3_1
X_10316_ net397 _05839_ vssd1 vssd1 vccd1 vccd1 _05948_ sky130_fd_sc_hd__nand2_1
X_11296_ net476 _06479_ net428 vssd1 vssd1 vccd1 vccd1 _06706_ sky130_fd_sc_hd__and3_1
XANTENNA__12006__B _06575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13035_ top.SPI.parameters\[19\] top.SPI.paroutput\[11\] net1356 vssd1 vssd1 vccd1
+ vccd1 _07443_ sky130_fd_sc_hd__mux2_1
XANTENNA__08003__B1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10247_ _05300_ _05367_ _05503_ _05507_ vssd1 vssd1 vccd1 vccd1 _05881_ sky130_fd_sc_hd__o211ai_1
XANTENNA__12721__S net1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09200__C1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1120 net1122 vssd1 vssd1 vccd1 vccd1 net1120 sky130_fd_sc_hd__clkbuf_4
Xfanout1131 net1136 vssd1 vssd1 vccd1 vccd1 net1131 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09751__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1142 net1143 vssd1 vssd1 vccd1 vccd1 net1142 sky130_fd_sc_hd__clkbuf_2
XFILLER_121_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1153 net1170 vssd1 vssd1 vccd1 vccd1 net1153 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_128_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10178_ net382 _05703_ vssd1 vssd1 vccd1 vccd1 _05814_ sky130_fd_sc_hd__or2_1
XANTENNA__08500__A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1164 net1170 vssd1 vssd1 vccd1 vccd1 net1164 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_128_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1175 net1179 vssd1 vssd1 vccd1 vccd1 net1175 sky130_fd_sc_hd__clkbuf_4
XFILLER_120_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1186 net1187 vssd1 vssd1 vccd1 vccd1 net1186 sky130_fd_sc_hd__buf_2
XANTENNA__08994__X _04633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1197 net1200 vssd1 vssd1 vccd1 vccd1 net1197 sky130_fd_sc_hd__clkbuf_4
X_14986_ clknet_leaf_84_clk _01231_ net1264 vssd1 vssd1 vccd1 vccd1 top.SPI.paroutput\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_167_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_167_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11310__B1 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_141_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12676__B top.CPU.alu.program_counter\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12819_ _07270_ _07271_ vssd1 vssd1 vccd1 vccd1 _07272_ sky130_fd_sc_hd__nor2_1
X_15607_ net1941 _01817_ net1181 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[407\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09267__C1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13799_ net2959 net338 net329 top.CPU.data_out\[1\] vssd1 vssd1 vccd1 vccd1 _02679_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13602__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15538_ net1872 _01748_ net1100 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[338\]
+ sky130_fd_sc_hd__dfrtp_1
X_15469_ net1803 _01679_ net1059 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[269\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08490__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12692__A top.CPU.alu.program_counter\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08010_ _03613_ _03647_ vssd1 vssd1 vccd1 vccd1 _03649_ sky130_fd_sc_hd__nand2_2
XANTENNA__12169__A2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09034__A2 net1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11377__B1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold603 top.CPU.registers.data\[709\] vssd1 vssd1 vccd1 vccd1 net3160 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11916__A2 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold614 top.CPU.registers.data\[910\] vssd1 vssd1 vccd1 vccd1 net3171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold625 top.CPU.registers.data\[565\] vssd1 vssd1 vccd1 vccd1 net3182 sky130_fd_sc_hd__dlygate4sd3_1
Xhold636 top.CPU.registers.data\[390\] vssd1 vssd1 vccd1 vccd1 net3193 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07596__A2 net1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold647 top.CPU.registers.data\[694\] vssd1 vssd1 vccd1 vccd1 net3204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 top.SPI.parameters\[20\] vssd1 vssd1 vccd1 vccd1 net3215 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09961_ _05399_ _05431_ _05436_ _05528_ vssd1 vssd1 vccd1 vccd1 _05600_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_90_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold669 top.CPU.registers.data\[531\] vssd1 vssd1 vccd1 vccd1 net3226 sky130_fd_sc_hd__dlygate4sd3_1
X_14350__520 clknet_leaf_121_clk vssd1 vssd1 vccd1 vccd1 net1989 sky130_fd_sc_hd__inv_2
XFILLER_143_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11129__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08912_ top.CPU.registers.data_out_r1_prev\[10\] net871 net691 _04543_ _04550_ vssd1
+ vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__o2111a_1
X_14647__817 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 net2286 sky130_fd_sc_hd__inv_2
XFILLER_131_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09892_ _04729_ _04698_ vssd1 vssd1 vccd1 vccd1 _05531_ sky130_fd_sc_hd__and2b_1
XANTENNA__10940__A _03167_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09742__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08843_ _04478_ _04479_ _04480_ _04481_ net672 net900 vssd1 vssd1 vccd1 vccd1 _04482_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09506__A net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1303 top.CPU.registers.data\[1021\] vssd1 vssd1 vccd1 vccd1 net3860 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10352__A1 _05793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1314 top.CPU.registers.data\[58\] vssd1 vssd1 vccd1 vccd1 net3871 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1325 top.I2C.output_state\[11\] vssd1 vssd1 vccd1 vccd1 net3882 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout289_A net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1336 top.CPU.registers.data\[794\] vssd1 vssd1 vccd1 vccd1 net3893 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10004__X _05643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1347 top.SPI.command\[6\] vssd1 vssd1 vccd1 vccd1 net3904 sky130_fd_sc_hd__dlygate4sd3_1
X_08774_ top.CPU.registers.data\[236\] net1388 net807 top.CPU.registers.data\[204\]
+ net767 vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__a221o_1
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1358 top.CPU.registers.data\[736\] vssd1 vssd1 vccd1 vccd1 net3915 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1369 top.I2C.data_out\[0\] vssd1 vssd1 vccd1 vccd1 net3926 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07725_ net923 _03362_ _03363_ net622 vssd1 vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__o211a_1
X_13837__7 clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 net1476 sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_158_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_158_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11301__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout456_A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_2_0_clk_X clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07656_ _03249_ _03259_ vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__nand2_1
XANTENNA__10655__A2 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08409__X _04048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09241__A net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10387__A _03756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09258__C1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07587_ top.CPU.registers.data\[287\] net865 vssd1 vssd1 vccd1 vccd1 _03226_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout244_X net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09326_ net726 _04960_ _04961_ _04964_ vssd1 vssd1 vccd1 vccd1 _04965_ sky130_fd_sc_hd__a31o_1
XANTENNA__07808__B1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09273__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09257_ top.CPU.registers.data\[325\] net1286 net1004 top.CPU.registers.data\[357\]
+ net926 vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout411_X net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08481__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1153_X net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08208_ top.CPU.registers.data\[311\] net1014 net937 vssd1 vssd1 vccd1 vccd1 _03847_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__08291__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08144__X _03783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09188_ _04823_ _04826_ net641 vssd1 vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout992_A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11368__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11907__A2 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08139_ top.CPU.registers.data\[245\] net1382 net993 top.CPU.registers.data\[213\]
+ net917 vssd1 vssd1 vccd1 vccd1 _03778_ sky130_fd_sc_hd__a221o_1
XANTENNA__09430__C1 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1320_X net1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08784__A1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11150_ net479 net456 _06634_ net301 net3424 vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__a32o_1
XFILLER_49_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout780_X net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10591__A1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14093__263 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 net1732 sky130_fd_sc_hd__inv_2
X_10101_ net391 net309 _05737_ vssd1 vssd1 vccd1 vccd1 _05739_ sky130_fd_sc_hd__and3_1
XANTENNA__13637__S net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07992__C1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11081_ net440 _06428_ net535 vssd1 vssd1 vccd1 vccd1 _06595_ sky130_fd_sc_hd__and3_1
XFILLER_150_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08536__A1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10032_ _03311_ _03322_ _03319_ vssd1 vssd1 vccd1 vccd1 _05671_ sky130_fd_sc_hd__a21oi_4
XANTENNA__08958__C net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09733__B1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_145_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11540__B1 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07744__C1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10894__A2 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input17_A DAT_I[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_149_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_149_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11983_ _06542_ net347 net182 net2839 vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__a22o_1
XANTENNA__12777__A top.CPU.alu.program_counter\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13372__S net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13722_ _07109_ _03060_ vssd1 vssd1 vccd1 vccd1 _03069_ sky130_fd_sc_hd__nand2_1
X_16510_ clknet_leaf_58_clk _02672_ net1144 vssd1 vssd1 vccd1 vccd1 top.mmio.mem_data_i\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_123_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10934_ net147 net437 vssd1 vssd1 vccd1 vccd1 _06514_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_86_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08466__S net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10568__Y _06190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12496__B _05190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16441_ clknet_leaf_80_clk net3048 net1241 vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__dfrtp_1
X_13653_ net3022 _07338_ net666 vssd1 vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__mux2_1
XANTENNA__16258__RESET_B net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10297__A _05367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10865_ net577 net502 vssd1 vssd1 vccd1 vccd1 _06472_ sky130_fd_sc_hd__or2_2
XFILLER_13_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12604_ top.SPI.timem\[21\] top.SPI.timem\[23\] top.SPI.timem\[22\] top.SPI.timem\[20\]
+ vssd1 vssd1 vccd1 vccd1 _07104_ sky130_fd_sc_hd__or4b_1
XFILLER_31_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16372_ clknet_leaf_76_clk _02581_ net1154 vssd1 vssd1 vccd1 vccd1 top.CPU.fetch.current_ra\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13584_ top.CPU.alu.program_counter\[14\] _06188_ net1352 vssd1 vssd1 vccd1 vccd1
+ _03017_ sky130_fd_sc_hd__mux2_1
X_10796_ _05754_ _05869_ _06405_ _06406_ vssd1 vssd1 vccd1 vccd1 _06407_ sky130_fd_sc_hd__o211a_1
XFILLER_158_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14791__961 clknet_leaf_184_clk vssd1 vssd1 vccd1 vccd1 net2430 sky130_fd_sc_hd__inv_2
X_15323_ net1657 _01533_ net1215 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[123\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12535_ _04991_ _05367_ _05541_ _05703_ vssd1 vssd1 vccd1 vccd1 _07044_ sky130_fd_sc_hd__and4_1
XFILLER_157_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15254_ net1588 _01464_ net1231 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_149_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12466_ _03610_ _03645_ _05330_ _05361_ vssd1 vssd1 vccd1 vccd1 _06975_ sky130_fd_sc_hd__a22oi_1
XANTENNA__11359__B1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_169_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_169_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11417_ _06552_ net277 net268 net2760 vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__a22o_1
X_14334__504 clknet_leaf_154_clk vssd1 vssd1 vccd1 vccd1 net1973 sky130_fd_sc_hd__inv_2
X_13998__168 clknet_leaf_166_clk vssd1 vssd1 vccd1 vccd1 net1637 sky130_fd_sc_hd__inv_2
XANTENNA__08224__B1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15185_ net1522 _01395_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r1_prev\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_12397_ top.I2C.inter_received top.I2C.I2C_state\[0\] net2624 vssd1 vssd1 vccd1 vccd1
+ _00030_ sky130_fd_sc_hd__a21o_1
XANTENNA__09421__C1 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11348_ net3487 net286 net279 _06193_ vssd1 vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__a22o_1
XFILLER_153_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07983__C1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11279_ net528 _06429_ net543 vssd1 vssd1 vccd1 vccd1 _06697_ sky130_fd_sc_hd__and3_1
XANTENNA__09724__A0 _05361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13018_ net2695 _07434_ net894 vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__mux2_1
XANTENNA__11531__B1 _06734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14969_ clknet_leaf_94_clk _01214_ net1260 vssd1 vssd1 vccd1 vccd1 top.SPI.paroutput\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12687__A top.CPU.alu.program_counter\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14876__1046 clknet_leaf_137_clk vssd1 vssd1 vccd1 vccd1 net2515 sky130_fd_sc_hd__inv_2
XANTENNA__12626__A3 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07510_ net1409 net1408 vssd1 vssd1 vccd1 vccd1 _03149_ sky130_fd_sc_hd__nand2b_1
XANTENNA__11591__A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10637__A2 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08490_ top.CPU.registers.data\[80\] net1321 net852 top.CPU.registers.data\[112\]
+ net770 vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__a221o_1
XANTENNA__08160__C1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10919__B net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13850__20 clknet_leaf_163_clk vssd1 vssd1 vccd1 vccd1 net1489 sky130_fd_sc_hd__inv_2
XFILLER_50_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09255__A2 net1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11598__A0 _05808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09111_ top.CPU.registers.data\[743\] net1393 net825 top.CPU.registers.data\[711\]
+ net724 vssd1 vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__a221o_1
XFILLER_149_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08463__B1 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13942__112 clknet_leaf_177_clk vssd1 vssd1 vccd1 vccd1 net1581 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_44_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09042_ _04677_ _04680_ net640 vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__a21o_1
XANTENNA__10654__B net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10146__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold400 top.CPU.registers.data\[619\] vssd1 vssd1 vccd1 vccd1 net2957 sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 top.I2C.output_state\[8\] vssd1 vssd1 vccd1 vccd1 net2968 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09412__C1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold422 top.CPU.registers.data\[471\] vssd1 vssd1 vccd1 vccd1 net2979 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout204_A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14077__247 clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 net1716 sky130_fd_sc_hd__inv_2
XANTENNA__11365__A3 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold433 top.CPU.registers.data\[406\] vssd1 vssd1 vccd1 vccd1 net2990 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold444 top.CPU.registers.data\[556\] vssd1 vssd1 vccd1 vccd1 net3001 sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 top.CPU.registers.data\[11\] vssd1 vssd1 vccd1 vccd1 net3012 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold466 top.CPU.registers.data\[965\] vssd1 vssd1 vccd1 vccd1 net3023 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11770__B1 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold477 top.CPU.registers.data\[868\] vssd1 vssd1 vccd1 vccd1 net3034 sky130_fd_sc_hd__dlygate4sd3_1
X_09944_ _04159_ _04190_ vssd1 vssd1 vccd1 vccd1 _05583_ sky130_fd_sc_hd__or2_1
Xfanout902 net903 vssd1 vssd1 vccd1 vccd1 net902 sky130_fd_sc_hd__clkbuf_4
Xhold488 top.CPU.registers.data\[789\] vssd1 vssd1 vccd1 vccd1 net3045 sky130_fd_sc_hd__dlygate4sd3_1
Xhold499 top.CPU.registers.data\[448\] vssd1 vssd1 vccd1 vccd1 net3056 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout913 net914 vssd1 vssd1 vccd1 vccd1 net913 sky130_fd_sc_hd__clkbuf_4
XFILLER_89_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1113_A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout924 net925 vssd1 vssd1 vccd1 vccd1 net924 sky130_fd_sc_hd__clkbuf_4
X_14118__288 clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 net1757 sky130_fd_sc_hd__inv_2
Xfanout935 net949 vssd1 vssd1 vccd1 vccd1 net935 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09715__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13511__B2 _02975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout946 net948 vssd1 vssd1 vccd1 vccd1 net946 sky130_fd_sc_hd__buf_2
XFILLER_38_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09875_ _03579_ _05509_ _05510_ _03511_ _03445_ vssd1 vssd1 vccd1 vccd1 _05514_ sky130_fd_sc_hd__a311o_1
XANTENNA_input9_A DAT_I[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout957 net962 vssd1 vssd1 vccd1 vccd1 net957 sky130_fd_sc_hd__buf_2
Xhold1100 top.I2C.I2C_state\[23\] vssd1 vssd1 vccd1 vccd1 net3657 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout968 net970 vssd1 vssd1 vccd1 vccd1 net968 sky130_fd_sc_hd__buf_2
XFILLER_38_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout194_X net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout573_A net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1111 top.CPU.registers.data\[1006\] vssd1 vssd1 vccd1 vccd1 net3668 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout979 net980 vssd1 vssd1 vccd1 vccd1 net979 sky130_fd_sc_hd__clkbuf_4
XFILLER_161_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08826_ _04431_ _04464_ vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_5_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1122 top.CPU.registers.data\[213\] vssd1 vssd1 vccd1 vccd1 net3679 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1133 net85 vssd1 vssd1 vccd1 vccd1 net3690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1144 top.CPU.registers.data\[140\] vssd1 vssd1 vccd1 vccd1 net3701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1155 top.CPU.registers.data\[964\] vssd1 vssd1 vccd1 vccd1 net3712 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07741__A2 net1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1166 top.CPU.registers.data\[1008\] vssd1 vssd1 vccd1 vccd1 net3723 sky130_fd_sc_hd__dlygate4sd3_1
X_08757_ _04394_ _04395_ vssd1 vssd1 vccd1 vccd1 _04396_ sky130_fd_sc_hd__and2b_1
Xhold1177 top.CPU.registers.data\[186\] vssd1 vssd1 vccd1 vccd1 net3734 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1188 top.CPU.registers.data\[71\] vssd1 vssd1 vccd1 vccd1 net3745 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout740_A net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout361_X net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1199 top.CPU.registers.data\[876\] vssd1 vssd1 vccd1 vccd1 net3756 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout838_A net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout459_X net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07708_ top.CPU.registers.data\[319\] top.CPU.registers.data\[287\] net999 vssd1
+ vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__mux2_1
X_08688_ _04294_ _04326_ vssd1 vssd1 vccd1 vccd1 _04327_ sky130_fd_sc_hd__nand2_1
XFILLER_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07639_ top.CPU.control_unit.instruction\[30\] _03258_ _03260_ vssd1 vssd1 vccd1
+ vccd1 _03278_ sky130_fd_sc_hd__and3_1
XFILLER_41_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14775__945 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 net2414 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_101_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout626_X net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1368_X net1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08129__S0 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10650_ _06239_ _06257_ _06267_ vssd1 vssd1 vccd1 vccd1 _06268_ sky130_fd_sc_hd__a21o_1
XFILLER_110_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09309_ net680 _04926_ _04927_ net613 vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__a31o_1
XFILLER_166_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07697__Y _03336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12250__A1 _06033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10581_ _06141_ _06201_ vssd1 vssd1 vccd1 vccd1 _06202_ sky130_fd_sc_hd__or2_1
XANTENNA__08454__B1 _04092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14816__986 clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 net2455 sky130_fd_sc_hd__inv_2
XFILLER_166_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13221__A _06948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12320_ net2591 _03716_ net1113 vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__mux2_1
XFILLER_10_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout995_X net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_39_Left_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08206__B1 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12251_ net3247 _06056_ net432 vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__mux2_1
XFILLER_163_971 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11202_ _06313_ _06644_ vssd1 vssd1 vccd1 vccd1 _06658_ sky130_fd_sc_hd__nor2_1
XFILLER_135_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12182_ net567 _06666_ net240 net171 net2900 vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__a32o_1
XFILLER_79_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08852__S1 net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_857 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11133_ _06624_ vssd1 vssd1 vccd1 vccd1 _06625_ sky130_fd_sc_hd__inv_2
XANTENNA__10580__A net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12271__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09706__B1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09146__A net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07980__A2 net1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15941_ net2275 _02151_ net1086 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[741\]
+ sky130_fd_sc_hd__dfrtp_1
X_11064_ _06212_ net534 vssd1 vssd1 vccd1 vccd1 _06589_ sky130_fd_sc_hd__and2_1
XFILLER_48_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07717__C1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11513__B1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10015_ _03243_ net379 vssd1 vssd1 vccd1 vccd1 _05654_ sky130_fd_sc_hd__nor2_1
XFILLER_23_1028 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15872_ net2206 _02082_ net1090 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[672\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10867__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12003__C net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_48_Left_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16439__RESET_B net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11615__S net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11816__A1 _06500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11966_ _06515_ net348 net231 net3462 vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__a22o_1
XFILLER_32_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13705_ net3400 _03056_ vssd1 vssd1 vccd1 vccd1 _02624_ sky130_fd_sc_hd__xor2_1
X_10917_ net142 net435 vssd1 vssd1 vccd1 vccd1 _06504_ sky130_fd_sc_hd__and2_1
X_11897_ net131 net3376 net188 vssd1 vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__mux2_1
XANTENNA__13569__A1 top.CPU.alu.program_counter\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16424_ clknet_leaf_54_clk _00006_ net1135 vssd1 vssd1 vccd1 vccd1 top.I2C.I2C_state\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_13636_ net3868 _07175_ net664 vssd1 vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__mux2_1
X_10848_ net382 _05701_ _06452_ vssd1 vssd1 vccd1 vccd1 _06456_ sky130_fd_sc_hd__or3_1
X_13567_ top.CPU.addressnew\[7\] _03006_ net581 vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__mux2_1
X_16355_ clknet_leaf_75_clk _02564_ net1154 vssd1 vssd1 vccd1 vccd1 top.CPU.fetch.current_ra\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12241__A1 _05808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10779_ net601 _06389_ _06390_ vssd1 vssd1 vccd1 vccd1 _06391_ sky130_fd_sc_hd__a21o_2
XANTENNA__13131__A _06887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_57_Left_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12792__A2 _04325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15306_ net1640 _01516_ net1085 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[106\]
+ sky130_fd_sc_hd__dfrtp_1
X_12518_ _06976_ _06985_ _06986_ _06978_ vssd1 vssd1 vccd1 vccd1 _07027_ sky130_fd_sc_hd__or4b_1
X_16286_ clknet_leaf_33_clk _02496_ net1120 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.toreg\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_13498_ _03369_ _02967_ net587 vssd1 vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__o21ai_4
XTAP_TAPCELL_ROW_136_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12449_ net3919 _06891_ _06904_ top.I2C.output_state\[0\] vssd1 vssd1 vccd1 vccd1
+ _00047_ sky130_fd_sc_hd__a22o_1
X_15237_ net1571 _01447_ net1065 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08748__A1 net1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15168_ net1505 _01378_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r1_prev\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10555__A1 _04294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08843__S1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11752__B1 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15099_ net1481 _01312_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r2_prev\[11\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout209 net210 vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__clkbuf_4
X_07990_ top.CPU.registers.data_out_r2_prev\[24\] net685 net618 _03621_ _03628_ vssd1
+ vssd1 vccd1 vccd1 _03629_ sky130_fd_sc_hd__o2111a_1
XFILLER_87_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09173__A1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_66_Left_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09660_ _05290_ _05292_ _05298_ _04125_ vssd1 vssd1 vccd1 vccd1 _05299_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_2_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10858__A2 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09490__S net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08611_ top.CPU.registers.data\[591\] net1375 net974 top.CPU.registers.data\[623\]
+ net903 vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__o221a_1
XFILLER_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09591_ _03151_ net1045 _03159_ _05229_ _03177_ vssd1 vssd1 vccd1 vccd1 _05230_ sky130_fd_sc_hd__a41o_1
X_14462__632 clknet_leaf_153_clk vssd1 vssd1 vccd1 vccd1 net2101 sky130_fd_sc_hd__inv_2
X_08542_ net909 _04180_ vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__or2_1
X_14759__929 clknet_leaf_183_clk vssd1 vssd1 vccd1 vccd1 net2398 sky130_fd_sc_hd__inv_2
XANTENNA__08133__C1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13009__B1 _07431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08473_ net958 _04109_ _04111_ net614 vssd1 vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_46_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16617__A net1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout154_A net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10491__B1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14503__673 clknet_leaf_183_clk vssd1 vssd1 vccd1 vccd1 net2142 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_63_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09228__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_75_Left_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_754 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11035__A2 _05769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08436__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout321_A net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1063_A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09025_ _04634_ _04663_ vssd1 vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__nand2_1
XANTENNA__11991__B1 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12880__A top.CPU.alu.program_counter\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11199__C net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout207_X net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1328_A net1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08739__A1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold230 top.CPU.registers.data\[169\] vssd1 vssd1 vccd1 vccd1 net2787 sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 top.CPU.registers.data\[554\] vssd1 vssd1 vccd1 vccd1 net2798 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10671__Y _06288_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout690_A net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold252 top.CPU.registers.data\[161\] vssd1 vssd1 vccd1 vccd1 net2809 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10546__B2 _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11743__B1 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold263 top.CPU.registers.data\[815\] vssd1 vssd1 vccd1 vccd1 net2820 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout788_A net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold274 _01267_ vssd1 vssd1 vccd1 vccd1 net2831 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07693__B _03262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold285 top.CPU.registers.data\[559\] vssd1 vssd1 vccd1 vccd1 net2842 sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 top.mmio.mem_data_i\[23\] vssd1 vssd1 vccd1 vccd1 net2853 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout710 net711 vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__clkbuf_4
XFILLER_172_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout721 net722 vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__buf_2
XFILLER_132_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout732 net734 vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07962__A2 net1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09927_ _04603_ _05283_ _05565_ vssd1 vssd1 vccd1 vccd1 _05566_ sky130_fd_sc_hd__and3_1
XANTENNA__12299__A1 _04633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout743 net746 vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout576_X net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout955_A net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout754 net759 vssd1 vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_142_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout765 net766 vssd1 vssd1 vccd1 vccd1 net765 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_142_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout776 net777 vssd1 vssd1 vccd1 vccd1 net776 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout787 net788 vssd1 vssd1 vccd1 vccd1 net787 sky130_fd_sc_hd__clkbuf_4
X_09858_ net628 _05488_ _05496_ vssd1 vssd1 vccd1 vccd1 _05497_ sky130_fd_sc_hd__and3_1
Xfanout798 net799 vssd1 vssd1 vccd1 vccd1 net798 sky130_fd_sc_hd__clkbuf_4
XFILLER_58_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07714__A2 _03154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08911__A1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08372__C1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08809_ net1283 _04446_ _04447_ vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__or3_1
XFILLER_100_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10399__X _06028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09789_ net627 _05424_ _05427_ _05422_ vssd1 vssd1 vccd1 vccd1 _05428_ sky130_fd_sc_hd__a31o_4
XANTENNA_fanout743_X net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11435__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11820_ net1401 _06657_ net233 net156 net2874 vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__a32o_1
XANTENNA__13799__B2 top.CPU.data_out\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09467__A2 net1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11751_ _06590_ net498 net192 net2863 vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout910_X net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11274__A2 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_80_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_121_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13650__S net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10702_ _05664_ _05979_ _06316_ vssd1 vssd1 vccd1 vccd1 _06317_ sky130_fd_sc_hd__o21a_1
XANTENNA__10482__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11682_ net459 _06503_ net234 net164 net3279 vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__a32o_1
X_13421_ top.mmio.mem_data_i\[31\] net593 net1345 vssd1 vssd1 vccd1 vccd1 _02933_
+ sky130_fd_sc_hd__a21o_1
X_10633_ net600 _06251_ vssd1 vssd1 vccd1 vccd1 _06252_ sky130_fd_sc_hd__nor2_1
XANTENNA__08427__B1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12266__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10575__A net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08316__Y _03955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08978__A1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16140_ net2474 _02350_ net1079 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[940\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_167_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13352_ top.I2C.data_out\[12\] net554 _02882_ net597 vssd1 vssd1 vccd1 vccd1 _02883_
+ sky130_fd_sc_hd__a22o_1
X_10564_ _05642_ _05722_ _06182_ _06185_ vssd1 vssd1 vccd1 vccd1 _06186_ sky130_fd_sc_hd__a211o_1
XFILLER_139_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12303_ net2586 _04889_ net1063 vssd1 vssd1 vccd1 vccd1 _01380_ sky130_fd_sc_hd__mux2_1
XANTENNA__11982__B1 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16071_ net2405 _02281_ net1197 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[871\]
+ sky130_fd_sc_hd__dfrtp_1
X_13283_ net3795 net3467 top.SPI.register\[1\] vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__mux2_1
XANTENNA__07650__A1 top.CPU.control_unit.instruction\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10495_ _05922_ _06113_ net405 vssd1 vssd1 vccd1 vccd1 _06120_ sky130_fd_sc_hd__mux2_1
XFILLER_5_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15022_ clknet_leaf_84_clk net2831 net1264 vssd1 vssd1 vccd1 vccd1 top.SPI.parameters\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09575__S net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14875__1045 clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 net2514 sky130_fd_sc_hd__inv_2
XANTENNA__12526__A2 _05265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12234_ _06697_ _06770_ _06883_ net168 net3172 vssd1 vssd1 vccd1 vccd1 _01444_ sky130_fd_sc_hd__a32o_1
XFILLER_6_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11734__B1 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12165_ net3763 net173 _06850_ vssd1 vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__a21o_1
XFILLER_123_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11116_ net573 net526 net439 _06057_ vssd1 vssd1 vccd1 vccd1 _06616_ sky130_fd_sc_hd__and4_1
XANTENNA__13487__A0 top.CPU.data_out\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12096_ top.CPU.registers.data\[104\] net645 vssd1 vssd1 vccd1 vccd1 _06816_ sky130_fd_sc_hd__or2_1
XANTENNA__09155__A1 _04793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_10_0_clk_X clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15924_ net2258 _02134_ net1112 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[724\]
+ sky130_fd_sc_hd__dfrtp_1
X_11047_ net3508 net367 _06582_ net324 vssd1 vssd1 vccd1 vccd1 _02330_ sky130_fd_sc_hd__a22o_1
X_14446__616 clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 net2085 sky130_fd_sc_hd__inv_2
Xinput9 DAT_I[16] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15855_ net2189 _02065_ net1104 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[655\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_92_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15786_ net2120 _01996_ net1085 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[586\]
+ sky130_fd_sc_hd__dfrtp_1
X_12998_ net1354 net1358 vssd1 vssd1 vccd1 vccd1 _07426_ sky130_fd_sc_hd__nand2_2
XFILLER_91_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11265__A2 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08666__B1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11949_ _06493_ net345 net230 net3560 vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_71_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_20_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16407_ clknet_leaf_56_clk net3213 net1145 vssd1 vssd1 vccd1 vccd1 top.I2C.I2C_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_138_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13619_ top.CPU.alu.program_counter\[28\] _05845_ net1351 vssd1 vssd1 vccd1 vccd1
+ _03038_ sky130_fd_sc_hd__mux2_1
XANTENNA__07778__B net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09615__C1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11080__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16338_ clknet_leaf_68_clk _02547_ net1165 vssd1 vssd1 vccd1 vccd1 top.CPU.addressnew\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10776__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11973__B1 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16269_ clknet_leaf_46_clk _02479_ net1137 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.toreg\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_69_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12517__A2 _04188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10932__B _06373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11725__B1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09394__A1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07944__A2 net1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07973_ top.CPU.alu.program_counter\[24\] net1033 vssd1 vssd1 vccd1 vccd1 _03612_
+ sky130_fd_sc_hd__nor2_1
XFILLER_101_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09712_ _05349_ _05350_ net946 vssd1 vssd1 vccd1 vccd1 _05351_ sky130_fd_sc_hd__mux2_1
XFILLER_19_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12150__B1 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08354__C1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09697__A2 net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12859__B _03916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14189__359 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 net1828 sky130_fd_sc_hd__inv_2
X_09643_ _04535_ _04601_ _04533_ vssd1 vssd1 vccd1 vccd1 _05282_ sky130_fd_sc_hd__a21o_1
XFILLER_55_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout271_A _06714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09574_ top.CPU.registers.data\[224\] top.CPU.registers.data\[192\] net973 vssd1
+ vssd1 vccd1 vccd1 _05213_ sky130_fd_sc_hd__mux2_1
XFILLER_43_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_180_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08106__C1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08525_ top.CPU.registers.data\[848\] net1290 net1011 top.CPU.registers.data\[880\]
+ net933 vssd1 vssd1 vccd1 vccd1 _04164_ sky130_fd_sc_hd__a221o_1
XANTENNA__12875__A top.CPU.alu.program_counter\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1180_A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout536_A net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09854__C1 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12453__B2 _03369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_62_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_60_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13470__S net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout157_X net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08456_ top.CPU.registers.data\[305\] top.CPU.registers.data\[273\] net988 vssd1
+ vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11008__A2 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12205__A1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10395__A net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13402__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09606__C1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_195_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08387_ net908 _04025_ _04024_ net626 vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout324_X net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout703_A _03212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09082__B1 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_75_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11964__B1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14590__760 clknet_leaf_153_clk vssd1 vssd1 vccd1 vccd1 net2229 sky130_fd_sc_hd__inv_2
XANTENNA_fanout1233_X net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12508__A2 _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09008_ top.CPU.registers.data\[457\] net1369 net964 top.CPU.registers.data\[489\]
+ net1364 vssd1 vssd1 vccd1 vccd1 _04647_ sky130_fd_sc_hd__o221a_1
X_10280_ _05785_ _05898_ _05912_ net395 vssd1 vssd1 vccd1 vccd1 _05913_ sky130_fd_sc_hd__o22a_1
XFILLER_105_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11716__B1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout693_X net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08188__A2 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1400_X net1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14133__303 clknet_leaf_173_clk vssd1 vssd1 vccd1 vccd1 net1772 sky130_fd_sc_hd__inv_2
XFILLER_120_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13469__B1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout860_X net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_133_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout540 net541 vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout958_X net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13645__S net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout551 _03172_ vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__buf_4
XANTENNA__09137__A1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout562 net564 vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__clkbuf_8
Xfanout573 net575 vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__buf_2
Xfanout584 net586 vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_13_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12921_ _07363_ _07360_ net129 vssd1 vssd1 vccd1 vccd1 _07364_ sky130_fd_sc_hd__mux2_1
XANTENNA__11495__A2 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_51 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_148_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15640_ net1974 _01850_ net1151 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[440\]
+ sky130_fd_sc_hd__dfrtp_1
X_12852_ top.CPU.alu.program_counter\[20\] _07301_ net1359 vssd1 vssd1 vccd1 vccd1
+ _01183_ sky130_fd_sc_hd__mux2_1
XFILLER_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11803_ _06649_ net241 net157 net3406 vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__a22o_1
X_12783_ _07237_ _07238_ vssd1 vssd1 vccd1 vccd1 _07239_ sky130_fd_sc_hd__nor2_1
X_15571_ net1905 _01781_ net1178 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[371\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11247__A2 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12785__A top.CPU.alu.program_counter\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_28_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09845__C1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_53_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__10455__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08112__A2 net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11734_ _06580_ net209 net194 net3719 vssd1 vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__a22o_1
XANTENNA__08743__S0 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11665_ net460 _06475_ net235 net164 net3031 vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__a32o_1
Xclkbuf_4_6_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_6_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_30_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13404_ _02830_ _02920_ vssd1 vssd1 vccd1 vccd1 _02921_ sky130_fd_sc_hd__nor2_1
X_10616_ _05564_ _05565_ _05532_ vssd1 vssd1 vccd1 vccd1 _06235_ sky130_fd_sc_hd__a21o_1
X_11596_ net3375 net215 net208 _06702_ vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__a22o_1
XFILLER_128_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09612__A2 net1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11955__B1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13335_ top.CPU.control_unit.instruction\[7\] _02870_ net667 vssd1 vssd1 vccd1 vccd1
+ _02441_ sky130_fd_sc_hd__mux2_1
X_16123_ net2457 _02333_ net1218 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[923\]
+ sky130_fd_sc_hd__dfrtp_1
X_10547_ _05641_ _05642_ _06167_ net413 _06166_ vssd1 vssd1 vccd1 vccd1 _06170_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_133_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10592__X _06213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13266_ net891 top.I2C.data_out\[3\] _02782_ vssd1 vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__mux2_1
XFILLER_109_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16054_ net2388 _02264_ net1221 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[854\]
+ sky130_fd_sc_hd__dfrtp_1
X_10478_ _06087_ _06102_ net600 vssd1 vssd1 vccd1 vccd1 _06104_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11707__B1 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09376__A1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15005_ clknet_leaf_94_clk _01250_ net1260 vssd1 vssd1 vccd1 vccd1 top.SPI.parameters\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_12217_ net360 _06745_ _06875_ net168 net3024 vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__a32o_1
X_13197_ top.I2C.output_state\[28\] top.I2C.which_data_address\[2\] _02775_ _02776_
+ vssd1 vssd1 vccd1 vccd1 _02777_ sky130_fd_sc_hd__and4_1
XFILLER_111_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12148_ top.CPU.registers.data\[78\] net648 _06749_ vssd1 vssd1 vccd1 vccd1 _06842_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__16454__RESET_B net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11864__A net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12079_ net563 net361 _06618_ _06808_ _06807_ vssd1 vssd1 vccd1 vccd1 _01524_ sky130_fd_sc_hd__a41o_1
XFILLER_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12132__B1 _06749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09679__A2 net1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14948__Q top.CPU.alu.program_counter\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15907_ net2241 _02117_ net1183 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[707\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11486__A2 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_139_Right_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08887__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15838_ net2172 _02048_ net1202 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[638\]
+ sky130_fd_sc_hd__dfrtp_1
X_15769_ net2103 _01979_ net1244 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[569\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_44_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_clk sky130_fd_sc_hd__clkbuf_8
X_08310_ net749 _03947_ _03948_ net695 vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_23_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11789__A3 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09290_ top.CPU.registers.data\[452\] net1299 net1020 top.CPU.registers.data\[484\]
+ net918 vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__a221o_1
XANTENNA__08384__S net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10997__B2 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09851__A2 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08241_ top.CPU.registers.data\[918\] net1330 net861 top.CPU.registers.data\[950\]
+ net728 vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__a221o_1
XFILLER_166_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14574__744 clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 net2213 sky130_fd_sc_hd__inv_2
XANTENNA__12199__B1 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11104__A net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13797__Y _03096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08172_ top.CPU.registers.data\[567\] top.CPU.registers.data\[535\] net824 vssd1
+ vssd1 vccd1 vccd1 _03811_ sky130_fd_sc_hd__mux2_1
XANTENNA__11410__A2 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10943__A _05693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14615__785 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 net2254 sky130_fd_sc_hd__inv_2
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__buf_2
XFILLER_161_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08413__A _04020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_974 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10381__C _06010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1026_A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08575__C1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07917__A2 net1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout486_A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07956_ net706 _03591_ _03592_ _03593_ _03594_ vssd1 vssd1 vccd1 vccd1 _03595_ sky130_fd_sc_hd__o32a_1
XANTENNA__08559__S net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07887_ top.CPU.registers.data\[188\] top.CPU.registers.data\[156\] net833 vssd1
+ vssd1 vccd1 vccd1 _03526_ sky130_fd_sc_hd__mux2_1
XANTENNA__11477__A2 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout653_A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout274_X net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_106_Right_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09626_ net640 _05263_ _05264_ _05250_ vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__o211a_2
XFILLER_102_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13623__A0 top.CPU.alu.program_counter\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14874__1044 clknet_leaf_162_clk vssd1 vssd1 vccd1 vccd1 net2513 sky130_fd_sc_hd__inv_2
X_09557_ top.CPU.registers.data\[64\] net1286 vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__and2_1
XANTENNA__11229__A2 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout441_X net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout820_A net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12809__S net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout918_A net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout539_X net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_35_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_8
X_08508_ net1048 _03164_ net1039 net1390 top.CPU.registers.data\[816\] vssd1 vssd1
+ vccd1 vccd1 _04147_ sky130_fd_sc_hd__o311a_1
X_09488_ _05124_ _05125_ vssd1 vssd1 vccd1 vccd1 _05127_ sky130_fd_sc_hd__nand2_2
XANTENNA__12503__A_N _04828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10988__B2 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08439_ net695 _04076_ _04077_ vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout706_X net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11450_ net3655 net265 _06724_ net487 vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__a22o_1
XANTENNA__09055__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11937__B1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10401_ _03789_ _05971_ net444 vssd1 vssd1 vccd1 vccd1 _06030_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_78_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11381_ net481 net471 _06496_ net271 net3190 vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__a32o_1
XANTENNA__11401__A2 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13120_ top.SPI.command\[6\] net1410 top.SPI.paroutput\[30\] net1358 vssd1 vssd1
+ vccd1 vccd1 _02725_ sky130_fd_sc_hd__a22o_1
XFILLER_109_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_12_Left_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10332_ net3471 net225 net313 _05963_ vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__a22o_1
XANTENNA__09419__A net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13051_ top.SPI.parameters\[27\] top.SPI.paroutput\[19\] net1358 vssd1 vssd1 vccd1
+ vccd1 _07451_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10263_ net403 _05894_ _05896_ _05643_ vssd1 vssd1 vccd1 vccd1 _05897_ sky130_fd_sc_hd__a211o_1
XFILLER_3_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08042__B net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12002_ _06573_ net342 net180 net2774 vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__a22o_1
XANTENNA__08566__C1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07908__A2 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1302 net1304 vssd1 vssd1 vccd1 vccd1 net1302 sky130_fd_sc_hd__clkbuf_4
X_10194_ net411 _05829_ vssd1 vssd1 vccd1 vccd1 _05830_ sky130_fd_sc_hd__and2_1
Xfanout1313 net1315 vssd1 vssd1 vccd1 vccd1 net1313 sky130_fd_sc_hd__clkbuf_4
XFILLER_87_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1324 net1327 vssd1 vssd1 vccd1 vccd1 net1324 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10912__B2 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1335 net1336 vssd1 vssd1 vccd1 vccd1 net1335 sky130_fd_sc_hd__clkbuf_4
Xfanout1346 net1347 vssd1 vssd1 vccd1 vccd1 net1346 sky130_fd_sc_hd__clkbuf_4
Xfanout1357 top.SPI.state\[2\] vssd1 vssd1 vccd1 vccd1 net1357 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08469__S net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout370 net371 vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__clkbuf_4
Xfanout1368 top.CPU.control_unit.instruction\[21\] vssd1 vssd1 vccd1 vccd1 net1368
+ sky130_fd_sc_hd__buf_4
Xfanout1379 net1380 vssd1 vssd1 vccd1 vccd1 net1379 sky130_fd_sc_hd__buf_4
Xfanout381 net382 vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__buf_2
XFILLER_93_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout392 net393 vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_21_Left_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12904_ top.CPU.alu.program_counter\[26\] _05499_ vssd1 vssd1 vccd1 vccd1 _07348_
+ sky130_fd_sc_hd__and2_1
XANTENNA__07541__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15623_ net1957 _01833_ net1201 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[423\]
+ sky130_fd_sc_hd__dfrtp_1
X_12835_ _07284_ _07285_ vssd1 vssd1 vccd1 vccd1 _07286_ sky130_fd_sc_hd__xnor2_1
XFILLER_36_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_26_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_174_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10428__B1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11623__S net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13404__A _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14261__431 clknet_leaf_173_clk vssd1 vssd1 vccd1 vccd1 net1900 sky130_fd_sc_hd__inv_2
X_15554_ net1888 _01764_ net1173 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[354\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12766_ top.CPU.alu.program_counter\[13\] _04392_ vssd1 vssd1 vccd1 vccd1 _07223_
+ sky130_fd_sc_hd__nor2_1
X_14558__728 clknet_leaf_152_clk vssd1 vssd1 vccd1 vccd1 net2197 sky130_fd_sc_hd__inv_2
XANTENNA__09833__A2 net1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11717_ _06556_ net199 net420 net2675 vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__a22o_1
X_12697_ net125 _07160_ vssd1 vssd1 vccd1 vccd1 _07161_ sky130_fd_sc_hd__nand2_1
X_15485_ net1819 _01695_ net1117 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[285\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11640__A2 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11648_ _06214_ net196 net424 net3675 vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__a22o_1
XANTENNA__09046__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14302__472 clknet_leaf_153_clk vssd1 vssd1 vccd1 vccd1 net1941 sky130_fd_sc_hd__inv_2
Xinput12 DAT_I[19] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput23 DAT_I[29] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__buf_1
XANTENNA__11928__B1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput34 en vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_2
XFILLER_128_554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11579_ _06690_ _06726_ net246 net3407 vssd1 vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__a2bb2o_1
Xhold807 top.CPU.registers.data\[648\] vssd1 vssd1 vccd1 vccd1 net3364 sky130_fd_sc_hd__dlygate4sd3_1
X_16106_ net2440 _02316_ net1084 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[906\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_143_524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13318_ _02830_ _02857_ vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__nor2_1
Xhold818 top.CPU.registers.data\[543\] vssd1 vssd1 vccd1 vccd1 net3375 sky130_fd_sc_hd__dlygate4sd3_1
Xhold829 top.CPU.registers.data\[701\] vssd1 vssd1 vccd1 vccd1 net3386 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16037_ net2371 _02247_ net1086 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[837\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_170_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13249_ net891 top.I2C.data_out\[11\] _02782_ vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__mux2_1
XFILLER_42_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08557__C1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09763__S net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08021__A1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11594__A net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07810_ top.CPU.registers.data\[765\] net1389 net816 top.CPU.registers.data\[733\]
+ net705 vssd1 vssd1 vccd1 vccd1 _03449_ sky130_fd_sc_hd__a221o_1
X_08790_ top.CPU.alu.program_counter\[12\] net878 vssd1 vssd1 vccd1 vccd1 _04429_
+ sky130_fd_sc_hd__nand2_1
XFILLER_69_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08309__C1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09064__A net1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07741_ top.CPU.registers.data\[670\] net1333 net864 top.CPU.registers.data\[702\]
+ net730 vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__a221o_1
XANTENNA__12202__B net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08324__A2 net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07672_ _03297_ _03304_ _03310_ vssd1 vssd1 vccd1 vccd1 _03311_ sky130_fd_sc_hd__and3_2
XFILLER_93_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10003__A net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09411_ top.CPU.registers.data\[899\] net1328 net859 top.CPU.registers.data\[931\]
+ net727 vssd1 vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__a221o_1
XFILLER_16_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13605__A0 top.CPU.alu.program_counter\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09809__C1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10938__A net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_17_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__13314__A _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09342_ top.CPU.registers.data\[324\] net1329 net860 top.CPU.registers.data\[356\]
+ net752 vssd1 vssd1 vccd1 vccd1 _04981_ sky130_fd_sc_hd__a221o_1
XANTENNA__08088__A1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09003__S net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09273_ top.CPU.registers.data_out_r2_prev\[5\] net686 _04910_ _04911_ net617 vssd1
+ vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__o221a_1
XANTENNA__11631__A2 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout234_A net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08224_ top.CPU.registers.data\[86\] net1337 net866 top.CPU.registers.data\[118\]
+ net779 vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__a221o_1
XANTENNA__08842__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11919__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08155_ top.CPU.registers.data\[183\] top.CPU.registers.data\[151\] net824 vssd1
+ vssd1 vccd1 vccd1 _03794_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout401_A net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1143_A net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08796__C1 net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08086_ top.CPU.registers.data\[565\] top.CPU.registers.data\[533\] net830 vssd1
+ vssd1 vccd1 vccd1 _03725_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1310_A net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12344__B1 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1408_A top.CPU.control_unit.instruction\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1029_X net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09673__S net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout770_A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11698__A2 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout489_X net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout868_A net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09760__A1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08289__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08988_ top.CPU.registers.data\[841\] net1309 net840 top.CPU.registers.data\[873\]
+ net761 vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__a221o_1
X_07939_ _03544_ _03577_ vssd1 vssd1 vccd1 vccd1 _03578_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout656_X net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10658__B1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11009__A _06333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09512__A1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10950_ net1403 net323 net542 vssd1 vssd1 vccd1 vccd1 _06525_ sky130_fd_sc_hd__nand3_1
XFILLER_28_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15940__RESET_B net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14245__415 clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 net1884 sky130_fd_sc_hd__inv_2
X_09609_ net788 _05242_ _05243_ net741 vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout823_X net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10881_ _05934_ _06471_ vssd1 vssd1 vccd1 vccd1 _06482_ sky130_fd_sc_hd__and2_1
XANTENNA__11870__A2 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11443__S net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12620_ _03127_ net1358 _07101_ _07116_ vssd1 vssd1 vccd1 vccd1 _00071_ sky130_fd_sc_hd__a22o_1
XANTENNA__08079__A1 _03685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09815__A2 net1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15083__SET_B net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12551_ top.CPU.done top.CPU.handler.state\[2\] _07054_ vssd1 vssd1 vccd1 vccd1 _07059_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_14_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11502_ _06635_ net260 net256 net3603 vssd1 vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__a22o_1
XFILLER_40_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12482_ _03610_ _03645_ vssd1 vssd1 vccd1 vccd1 _06991_ sky130_fd_sc_hd__nor2_1
X_15270_ net1604 _01480_ net1074 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[70\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10854__Y _06462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11433_ _06577_ net283 net265 net3106 vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__a22o_1
XFILLER_153_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11017__C_N net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11364_ top.CPU.registers.data\[735\] net273 vssd1 vssd1 vccd1 vccd1 _06715_ sky130_fd_sc_hd__and2_1
XFILLER_125_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13103_ top.SPI.count\[1\] top.SPI.count\[0\] _02713_ vssd1 vssd1 vccd1 vccd1 _02716_
+ sky130_fd_sc_hd__and3_1
X_10315_ _03646_ net507 vssd1 vssd1 vccd1 vccd1 _05947_ sky130_fd_sc_hd__nand2_1
XFILLER_125_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13926__96 clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 net1565 sky130_fd_sc_hd__inv_2
XFILLER_152_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11295_ net3459 net291 net359 net135 vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__a22o_1
XANTENNA__08539__C1 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13034_ net3088 _07442_ net894 vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_167_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10246_ net3735 net226 net317 _05880_ vssd1 vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__a22o_1
XANTENNA__08003__A1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11689__A2 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1110 net1111 vssd1 vssd1 vccd1 vccd1 net1110 sky130_fd_sc_hd__buf_2
XFILLER_121_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1121 net1122 vssd1 vssd1 vccd1 vccd1 net1121 sky130_fd_sc_hd__buf_2
XFILLER_26_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11618__S net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1132 net1133 vssd1 vssd1 vccd1 vccd1 net1132 sky130_fd_sc_hd__clkbuf_4
XFILLER_152_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10177_ _05509_ net447 _05812_ vssd1 vssd1 vccd1 vccd1 _05813_ sky130_fd_sc_hd__and3_1
XFILLER_113_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1143 net1146 vssd1 vssd1 vccd1 vccd1 net1143 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_128_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1154 net1157 vssd1 vssd1 vccd1 vccd1 net1154 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10361__A2 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07762__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1165 net1169 vssd1 vssd1 vccd1 vccd1 net1165 sky130_fd_sc_hd__clkbuf_4
XFILLER_120_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1176 net1179 vssd1 vssd1 vccd1 vccd1 net1176 sky130_fd_sc_hd__clkbuf_2
X_14985_ clknet_leaf_93_clk _01230_ net1267 vssd1 vssd1 vccd1 vccd1 top.SPI.paroutput\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1187 net1188 vssd1 vssd1 vccd1 vccd1 net1187 sky130_fd_sc_hd__buf_2
XANTENNA__12022__B net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1198 net1200 vssd1 vssd1 vccd1 vccd1 net1198 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08306__A2 net1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11310__B2 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11861__A2 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12676__C top.CPU.alu.program_counter\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15606_ net1940 _01816_ net1227 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[406\]
+ sky130_fd_sc_hd__dfrtp_1
X_12818_ top.CPU.alu.program_counter\[17\] _07260_ vssd1 vssd1 vccd1 vccd1 _07271_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__13063__A1 top.CPU.data_out\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13798_ net2745 net335 net328 top.CPU.data_out\[0\] vssd1 vssd1 vccd1 vccd1 _02678_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09806__A2 net1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15537_ net1871 _01747_ net1105 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[337\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07817__A1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12749_ top.CPU.alu.program_counter\[11\] _07191_ vssd1 vssd1 vccd1 vccd1 _07208_
+ sky130_fd_sc_hd__and2_1
XANTENNA__11613__A2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14029__199 clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 net1668 sky130_fd_sc_hd__inv_2
XFILLER_72_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10821__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15468_ net1802 _01678_ net1071 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[268\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12692__B _04856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11589__A net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13366__A2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15399_ net1733 _01609_ net1200 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[199\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_144_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08778__C1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold604 top.CPU.fetch.current_ra\[7\] vssd1 vssd1 vccd1 vccd1 net3161 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08242__A1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold615 top.CPU.registers.data\[34\] vssd1 vssd1 vccd1 vccd1 net3172 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold626 top.CPU.registers.data\[274\] vssd1 vssd1 vccd1 vccd1 net3183 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13118__A2 net1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold637 top.SPI.parameters\[15\] vssd1 vssd1 vccd1 vccd1 net3194 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold648 top.CPU.registers.data\[211\] vssd1 vssd1 vccd1 vccd1 net3205 sky130_fd_sc_hd__dlygate4sd3_1
X_09960_ _05503_ _05598_ _05528_ vssd1 vssd1 vccd1 vccd1 _05599_ sky130_fd_sc_hd__a21oi_1
X_14873__1043 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 net2512 sky130_fd_sc_hd__inv_2
Xhold659 top.CPU.registers.data\[532\] vssd1 vssd1 vccd1 vccd1 net3216 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_6_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__11129__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08911_ net741 _04545_ _04546_ _04549_ net636 vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__a311o_1
X_14686__856 clknet_leaf_154_clk vssd1 vssd1 vccd1 vccd1 net2325 sky130_fd_sc_hd__inv_2
X_09891_ _04260_ _04330_ vssd1 vssd1 vccd1 vccd1 _05530_ sky130_fd_sc_hd__and2_1
XFILLER_69_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10940__B _06447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10888__B1 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08545__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08842_ top.CPU.registers.data\[875\] top.CPU.registers.data\[843\] net964 vssd1
+ vssd1 vccd1 vccd1 _04481_ sky130_fd_sc_hd__mux2_1
Xhold1304 top.CPU.registers.data\[116\] vssd1 vssd1 vccd1 vccd1 net3861 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_98_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1315 top.CPU.registers.data\[36\] vssd1 vssd1 vccd1 vccd1 net3872 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1326 top.CPU.registers.data\[120\] vssd1 vssd1 vccd1 vccd1 net3883 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1337 top.CPU.handler.toreg\[5\] vssd1 vssd1 vccd1 vccd1 net3894 sky130_fd_sc_hd__dlygate4sd3_1
X_08773_ top.CPU.registers.data\[172\] top.CPU.registers.data\[140\] net808 vssd1
+ vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__mux2_1
XANTENNA__13826__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14727__897 clknet_leaf_183_clk vssd1 vssd1 vccd1 vccd1 net2366 sky130_fd_sc_hd__inv_2
Xhold1348 top.CPU.registers.data\[121\] vssd1 vssd1 vccd1 vccd1 net3905 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1359 top.CPU.registers.data\[94\] vssd1 vssd1 vccd1 vccd1 net3916 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout184_A net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07724_ net681 _03341_ net947 _03338_ vssd1 vssd1 vccd1 vccd1 _03363_ sky130_fd_sc_hd__a211o_1
XFILLER_66_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08702__C1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09522__A net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07655_ net1038 _03293_ vssd1 vssd1 vccd1 vccd1 _03294_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11852__A2 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout351_A net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1093_A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12586__C _07089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07586_ top.CPU.control_unit.instruction\[19\] _03200_ vssd1 vssd1 vccd1 vccd1 _03225_
+ sky130_fd_sc_hd__or2_1
XANTENNA__09258__B1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10387__B net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09325_ net752 _04962_ _04963_ net637 vssd1 vssd1 vccd1 vccd1 _04964_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_66_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout237_X net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1358_A top.SPI.state\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09256_ top.CPU.registers.data\[421\] top.CPU.registers.data\[389\] top.CPU.registers.data\[293\]
+ top.CPU.registers.data\[261\] net966 net901 vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_32_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08481__A1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08572__S net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08207_ top.CPU.registers.data\[407\] net987 _03845_ vssd1 vssd1 vccd1 vccd1 _03846_
+ sky130_fd_sc_hd__a21o_1
XFILLER_138_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09187_ net704 _04824_ _04825_ vssd1 vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout404_X net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1146_X net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08769__C1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08138_ top.CPU.registers.data\[85\] net1300 net1021 top.CPU.registers.data\[117\]
+ net940 vssd1 vssd1 vccd1 vccd1 _03777_ sky130_fd_sc_hd__a221o_1
X_14630__800 clknet_leaf_123_clk vssd1 vssd1 vccd1 vccd1 net2269 sky130_fd_sc_hd__inv_2
XANTENNA__08233__A1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout985_A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08069_ top.CPU.registers.data\[436\] net1008 net905 vssd1 vssd1 vccd1 vccd1 _03708_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_108_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1313_X net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10100_ net308 _05737_ vssd1 vssd1 vccd1 vccd1 _05738_ sky130_fd_sc_hd__and2_1
XANTENNA__10591__A2 _06210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07992__B1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07916__S net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11080_ net148 net3689 net368 vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__mux2_1
XFILLER_108_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout773_X net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10031_ net509 vssd1 vssd1 vccd1 vccd1 _05670_ sky130_fd_sc_hd__inv_2
XANTENNA__13219__A top.I2C.output_state\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11540__A1 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07744__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout940_X net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13653__S net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11982_ _06540_ net346 net181 net2805 vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__a22o_1
XANTENNA__12777__B _04325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13721_ top.SPI.timem\[11\] top.SPI.timem\[10\] _03064_ vssd1 vssd1 vccd1 vccd1 _03068_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_123_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10933_ net479 net456 _06513_ net220 net3023 vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_86_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12269__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11843__A2 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11173__S net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16440_ clknet_leaf_80_clk _02603_ net1241 vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__dfrtp_1
X_13652_ net3101 _07334_ net666 vssd1 vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__mux2_1
XANTENNA__09249__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10864_ net576 net502 vssd1 vssd1 vccd1 vccd1 _06471_ sky130_fd_sc_hd__nor2_2
XFILLER_71_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12603_ _07102_ top.SPI.nextwrx vssd1 vssd1 vccd1 vccd1 _07103_ sky130_fd_sc_hd__and2_1
X_16371_ clknet_leaf_71_clk _02580_ net1169 vssd1 vssd1 vccd1 vccd1 top.CPU.fetch.current_ra\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_13583_ net3974 _03016_ net580 vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__mux2_1
X_10795_ _05056_ net508 net504 _05058_ net443 vssd1 vssd1 vccd1 vccd1 _06406_ sky130_fd_sc_hd__o221a_1
XFILLER_13_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10865__X _06472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09578__S net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10803__B1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15322_ net1656 _01532_ net1243 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[122\]
+ sky130_fd_sc_hd__dfrtp_1
X_12534_ _03650_ _05127_ _06402_ _07042_ vssd1 vssd1 vccd1 vccd1 _07043_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_30_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15253_ net1587 _01463_ net1228 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16227__RESET_B net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12465_ _06969_ _06970_ _06973_ vssd1 vssd1 vccd1 vccd1 _06974_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_169_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11416_ _06551_ net275 net267 net3043 vssd1 vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_169_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12396_ _06917_ net560 vssd1 vssd1 vccd1 vccd1 _07456_ sky130_fd_sc_hd__nand2_1
XANTENNA__09421__B1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15184_ net1521 _01394_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r1_prev\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_14373__543 clknet_leaf_112_clk vssd1 vssd1 vccd1 vccd1 net2012 sky130_fd_sc_hd__inv_2
X_11347_ net3911 net287 net276 _06175_ vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__a22o_1
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07983__B1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07826__S net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09607__A net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11278_ net2928 net295 _06696_ net317 vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__a22o_1
X_14414__584 clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 net2053 sky130_fd_sc_hd__inv_2
XFILLER_3_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09724__A1 _05362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09185__C1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08527__A2 net1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10229_ net395 _05660_ vssd1 vssd1 vccd1 vccd1 _05864_ sky130_fd_sc_hd__nor2_1
X_13017_ top.SPI.parameters\[10\] top.SPI.paroutput\[2\] net1355 vssd1 vssd1 vccd1
+ vccd1 _07434_ sky130_fd_sc_hd__mux2_1
XFILLER_67_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11531__B2 _06500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1 top.CPU.handler.next_counter_on vssd1 vssd1 vccd1 vccd1 net2558 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14968_ clknet_leaf_97_clk net3065 net1253 vssd1 vssd1 vccd1 vccd1 top.SPI.paroutput\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12087__A2 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10098__A1 _03315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11591__B net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11295__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11834__A2 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10919__C net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09110_ top.CPU.registers.data\[583\] net1327 net858 top.CPU.registers.data\[615\]
+ net749 vssd1 vssd1 vccd1 vccd1 _04749_ sky130_fd_sc_hd__a221o_1
XFILLER_148_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13981__151 clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 net1620 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_44_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09041_ net703 _04678_ _04679_ vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__or3_1
XANTENNA__13339__A2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10654__C net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11112__A net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold401 top.CPU.registers.data\[464\] vssd1 vssd1 vccd1 vccd1 net2958 sky130_fd_sc_hd__dlygate4sd3_1
Xhold412 _06897_ vssd1 vssd1 vccd1 vccd1 net2969 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold423 top.CPU.registers.data\[348\] vssd1 vssd1 vccd1 vccd1 net2980 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold434 top.CPU.registers.data\[816\] vssd1 vssd1 vccd1 vccd1 net2991 sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 top.CPU.registers.data\[176\] vssd1 vssd1 vccd1 vccd1 net3002 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10951__A net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold456 top.CPU.registers.data\[449\] vssd1 vssd1 vccd1 vccd1 net3013 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11770__A1 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold467 top.CPU.registers.data\[43\] vssd1 vssd1 vccd1 vccd1 net3024 sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 top.CPU.registers.data\[425\] vssd1 vssd1 vccd1 vccd1 net3035 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09943_ _03684_ _03718_ vssd1 vssd1 vccd1 vccd1 _05582_ sky130_fd_sc_hd__nor2_1
Xhold489 top.CPU.registers.data\[939\] vssd1 vssd1 vccd1 vccd1 net3046 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout903 net910 vssd1 vssd1 vccd1 vccd1 net903 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout914 net925 vssd1 vssd1 vccd1 vccd1 net914 sky130_fd_sc_hd__buf_2
XANTENNA__09176__C1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout925 _03353_ vssd1 vssd1 vccd1 vccd1 net925 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout399_A net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout936 net938 vssd1 vssd1 vccd1 vccd1 net936 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09715__A1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09874_ _05512_ vssd1 vssd1 vccd1 vccd1 _05513_ sky130_fd_sc_hd__inv_2
Xfanout947 net948 vssd1 vssd1 vccd1 vccd1 net947 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10325__A2 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07726__B1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout958 net961 vssd1 vssd1 vccd1 vccd1 net958 sky130_fd_sc_hd__buf_4
Xhold1101 _00032_ vssd1 vssd1 vccd1 vccd1 net3658 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11522__B2 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout969 net970 vssd1 vssd1 vccd1 vccd1 net969 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1106_A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1112 top.CPU.registers.data\[752\] vssd1 vssd1 vccd1 vccd1 net3669 sky130_fd_sc_hd__dlygate4sd3_1
X_08825_ _04460_ _04463_ net452 vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__mux2_1
Xhold1123 top.CPU.registers.data\[1003\] vssd1 vssd1 vccd1 vccd1 net3680 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1134 _02703_ vssd1 vssd1 vccd1 vccd1 net3691 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_86_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout566_A net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout187_X net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1145 top.CPU.registers.data\[142\] vssd1 vssd1 vccd1 vccd1 net3702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1156 top.CPU.registers.data\[744\] vssd1 vssd1 vccd1 vccd1 net3713 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1167 top.CPU.registers.data\[486\] vssd1 vssd1 vccd1 vccd1 net3724 sky130_fd_sc_hd__dlygate4sd3_1
X_08756_ _04363_ _04393_ vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__nand2_1
Xhold1178 top.CPU.registers.data\[1019\] vssd1 vssd1 vccd1 vccd1 net3735 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11970__D_N net1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1189 top.CPU.registers.data\[88\] vssd1 vssd1 vccd1 vccd1 net3746 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07707_ top.CPU.registers.data\[895\] top.CPU.registers.data\[863\] net999 vssd1
+ vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__mux2_1
XANTENNA__11825__A2 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08687_ _04324_ _04325_ net453 vssd1 vssd1 vccd1 vccd1 _04326_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout733_A net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout354_X net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07638_ top.CPU.control_unit.instruction\[4\] _03177_ _03274_ _03275_ _03276_ vssd1
+ vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13578__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10548__D _06170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08129__S1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10685__X _06301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout900_A net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout521_X net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07569_ net1048 _03164_ net1039 top.CPU.control_unit.instruction\[17\] vssd1 vssd1
+ vccd1 vccd1 _03208_ sky130_fd_sc_hd__o31a_1
XFILLER_55_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1263_X net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout619_X net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09100__C1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13502__A _04593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09308_ net680 _04928_ _04929_ _04946_ vssd1 vssd1 vccd1 vccd1 _04947_ sky130_fd_sc_hd__a31o_1
X_10580_ net402 _05674_ vssd1 vssd1 vccd1 vccd1 _06201_ sky130_fd_sc_hd__nor2_1
XANTENNA__08454__A1 _03198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14060__230 clknet_leaf_195_clk vssd1 vssd1 vccd1 vccd1 net1699 sky130_fd_sc_hd__inv_2
XFILLER_166_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14357__527 clknet_leaf_173_clk vssd1 vssd1 vccd1 vccd1 net1996 sky130_fd_sc_hd__inv_2
X_09239_ top.CPU.registers.data\[581\] net1313 net844 top.CPU.registers.data\[613\]
+ net737 vssd1 vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__a221o_1
XFILLER_166_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12250_ net2865 _06033_ net433 vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout890_X net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12002__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11210__A0 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11201_ net144 net3572 net297 vssd1 vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout988_X net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14101__271 clknet_leaf_173_clk vssd1 vssd1 vccd1 vccd1 net1740 sky130_fd_sc_hd__inv_2
XANTENNA__09954__A1 _03822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13648__S net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12181_ _06740_ net237 net169 net3566 vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__a22o_1
XFILLER_163_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10861__A net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10564__A2 _05722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07965__B1 net1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11132_ net551 net515 _06232_ vssd1 vssd1 vccd1 vccd1 _06624_ sky130_fd_sc_hd__or3_1
XFILLER_79_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold990 top.CPU.registers.data\[655\] vssd1 vssd1 vccd1 vccd1 net3547 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_164_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11168__S net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08509__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15940_ net2274 _02150_ net1212 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[740\]
+ sky130_fd_sc_hd__dfrtp_1
X_11063_ net3171 net367 _06588_ net314 vssd1 vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__a22o_1
XFILLER_135_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12710__A0 top.CPU.alu.program_counter\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11513__A1 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10014_ net384 net374 _03407_ vssd1 vssd1 vccd1 vccd1 _05653_ sky130_fd_sc_hd__or3b_1
XANTENNA__09861__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08914__C1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09182__A2 net1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_160_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15871_ net2205 _02081_ net1199 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[671\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10867__A3 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12003__D net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11965_ _06514_ net348 net231 net3541 vssd1 vssd1 vccd1 vccd1 _01606_ sky130_fd_sc_hd__a22o_1
XFILLER_44_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11816__A2 _06648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08142__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13704_ _03056_ _03057_ vssd1 vssd1 vccd1 vccd1 _02623_ sky130_fd_sc_hd__nor2_1
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10916_ net483 net459 _06503_ net220 net3131 vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__a32o_1
X_14872__1042 clknet_leaf_160_clk vssd1 vssd1 vccd1 vccd1 net2511 sky130_fd_sc_hd__inv_2
XFILLER_71_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11896_ _06711_ net241 net191 net2738 vssd1 vssd1 vccd1 vccd1 _01667_ sky130_fd_sc_hd__a22o_1
X_16423_ clknet_leaf_56_clk _00005_ net1142 vssd1 vssd1 vccd1 vccd1 top.I2C.I2C_state\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13965__135 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 net1604 sky130_fd_sc_hd__inv_2
X_13635_ net3161 _07166_ net664 vssd1 vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__mux2_1
XANTENNA__16408__RESET_B net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10847_ _05268_ net504 _05754_ _05937_ _06454_ vssd1 vssd1 vccd1 vccd1 _06455_ sky130_fd_sc_hd__o221a_1
XFILLER_158_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13412__A net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16354_ clknet_leaf_75_clk _02563_ net1158 vssd1 vssd1 vccd1 vccd1 top.CPU.fetch.current_ra\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08445__A1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13566_ top.CPU.alu.program_counter\[7\] _06331_ net1349 vssd1 vssd1 vccd1 vccd1
+ _03006_ sky130_fd_sc_hd__mux2_1
X_10778_ top.CPU.fetch.current_ra\[4\] net1040 net633 top.CPU.handler.toreg\[4\] vssd1
+ vssd1 vccd1 vccd1 _06390_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_4_Left_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09101__S net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15305_ net1639 _01515_ net1055 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[105\]
+ sky130_fd_sc_hd__dfrtp_1
X_12517_ _04155_ _04188_ _06979_ _06984_ _06992_ vssd1 vssd1 vccd1 vccd1 _07026_ sky130_fd_sc_hd__o2111ai_1
X_16285_ clknet_leaf_58_clk _02495_ net1145 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.toreg\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_117_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13497_ _04726_ _02966_ vssd1 vssd1 vccd1 vccd1 _02968_ sky130_fd_sc_hd__nor2_1
XFILLER_9_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15236_ net1570 _01446_ net1212 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[36\]
+ sky130_fd_sc_hd__dfrtp_1
X_12448_ net1054 _06960_ vssd1 vssd1 vccd1 vccd1 _00048_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_136_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11201__A0 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15167_ net1504 _01377_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r1_prev\[2\]
+ sky130_fd_sc_hd__dfxtp_2
X_12379_ _03127_ top.SPI.state\[5\] vssd1 vssd1 vccd1 vccd1 _06917_ sky130_fd_sc_hd__or2_1
XFILLER_125_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15098_ net1480 _01311_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r2_prev\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_141_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16231__Q top.CPU.control_unit.instruction\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12477__A1_N net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11504__B2 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12698__A top.CPU.alu.program_counter\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13910__80 clknet_leaf_178_clk vssd1 vssd1 vccd1 vccd1 net1549 sky130_fd_sc_hd__inv_2
XANTENNA__08895__B _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11806__S net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13146__X _02738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08610_ top.CPU.registers.data\[719\] net1375 net976 top.CPU.registers.data\[751\]
+ net929 vssd1 vssd1 vccd1 vccd1 _04249_ sky130_fd_sc_hd__o221a_1
X_09590_ _03144_ _03157_ net1363 vssd1 vssd1 vccd1 vccd1 _05229_ sky130_fd_sc_hd__a21o_1
XFILLER_67_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14798__968 clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 net2437 sky130_fd_sc_hd__inv_2
X_08541_ top.CPU.registers.data\[688\] top.CPU.registers.data\[656\] net984 vssd1
+ vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__mux2_1
XFILLER_70_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08133__B1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08472_ net919 _04110_ vssd1 vssd1 vccd1 vccd1 _04111_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_46_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08684__A1 _03342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14925__RESET_B net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14044__214 clknet_leaf_140_clk vssd1 vssd1 vccd1 vccd1 net1683 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_63_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07892__C1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout147_A _06391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12232__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10243__A1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout314_A net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09024_ net452 _04658_ _04661_ vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout1056_A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09397__C1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold220 top.CPU.registers.data\[969\] vssd1 vssd1 vccd1 vccd1 net2777 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10681__A net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold231 top.CPU.registers.data\[396\] vssd1 vssd1 vccd1 vccd1 net2788 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold242 top.I2C.data_out\[31\] vssd1 vssd1 vccd1 vccd1 net2799 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold253 net87 vssd1 vssd1 vccd1 vccd1 net2810 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11743__A1 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_1004 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold264 top.CPU.registers.data\[942\] vssd1 vssd1 vccd1 vccd1 net2821 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold275 top.CPU.registers.data\[162\] vssd1 vssd1 vccd1 vccd1 net2832 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout683_A net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold286 top.CPU.registers.data\[312\] vssd1 vssd1 vccd1 vccd1 net2843 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout700 net701 vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__clkbuf_4
Xhold297 top.CPU.fetch.current_ra\[29\] vssd1 vssd1 vccd1 vccd1 net2854 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09149__C1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout711 net712 vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__clkbuf_4
X_09926_ _04732_ _05279_ vssd1 vssd1 vccd1 vccd1 _05565_ sky130_fd_sc_hd__and2_1
Xfanout722 net736 vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__buf_2
XFILLER_131_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13496__A1 net1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout733 net734 vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__clkbuf_2
Xfanout744 net746 vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1109_X net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout755 net759 vssd1 vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__buf_2
XANTENNA__09164__A2 net1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14742__912 clknet_leaf_181_clk vssd1 vssd1 vccd1 vccd1 net2381 sky130_fd_sc_hd__inv_2
Xfanout766 net772 vssd1 vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__clkbuf_4
Xfanout777 net782 vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__buf_2
X_09857_ net960 _05490_ _05492_ _05495_ vssd1 vssd1 vccd1 vccd1 _05496_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout850_A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout788 net794 vssd1 vssd1 vccd1 vccd1 net788 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout471_X net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout569_X net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout799 net804 vssd1 vssd1 vccd1 vccd1 net799 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08372__B1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout948_A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08808_ top.CPU.registers.data\[844\] net1372 net977 top.CPU.registers.data\[876\]
+ net1282 vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__o221a_1
XANTENNA__13248__B2 _02803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09788_ net613 _05425_ _05426_ vssd1 vssd1 vccd1 vccd1 _05427_ sky130_fd_sc_hd__or3_1
XFILLER_39_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13799__A2 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08739_ net624 _04370_ _04376_ _04377_ vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1380_X net1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13949__119 clknet_leaf_130_clk vssd1 vssd1 vccd1 vccd1 net1588 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_83_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout736_X net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11017__A net1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11750_ net145 net535 net498 net192 net2657 vssd1 vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__a32o_1
XFILLER_157_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10701_ _05757_ _05978_ _05671_ vssd1 vssd1 vccd1 vccd1 _06316_ sky130_fd_sc_hd__a21o_1
XFILLER_92_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07883__C1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11681_ _06502_ net196 net164 net3684 vssd1 vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout903_X net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11451__S net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13420_ top.CPU.control_unit.instruction\[30\] _02932_ net670 vssd1 vssd1 vccd1 vccd1
+ _02464_ sky130_fd_sc_hd__mux2_1
XFILLER_139_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10632_ _06237_ _06240_ _06250_ vssd1 vssd1 vccd1 vccd1 _06251_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_157_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13420__A1 _02932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12223__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10563_ net550 _04330_ _06184_ vssd1 vssd1 vccd1 vccd1 _06185_ sky130_fd_sc_hd__o21ai_1
X_13351_ top.mmio.mem_data_i\[12\] net592 net1344 vssd1 vssd1 vccd1 vccd1 _02882_
+ sky130_fd_sc_hd__a21o_1
XFILLER_155_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12302_ net2587 _04828_ net1082 vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__mux2_1
X_16070_ net2404 _02280_ net1072 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[870\]
+ sky130_fd_sc_hd__dfrtp_1
X_13282_ top.CPU.handler.readout _02826_ _02827_ _02828_ vssd1 vssd1 vccd1 vccd1 _01374_
+ sky130_fd_sc_hd__a31o_1
X_10494_ _05733_ _05919_ _05924_ _05753_ _06118_ vssd1 vssd1 vccd1 vccd1 _06119_ sky130_fd_sc_hd__a221o_1
XANTENNA__08760__S net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12790__B _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10862__Y _06469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15021_ clknet_leaf_83_clk net2883 net1261 vssd1 vssd1 vccd1 vccd1 top.SPI.parameters\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_108_663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12233_ top.CPU.registers.data\[34\] net647 vssd1 vssd1 vccd1 vccd1 _06883_ sky130_fd_sc_hd__or2_1
XANTENNA__07938__A0 _03575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09157__A _04765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12164_ top.CPU.registers.data\[70\] net649 _06355_ net361 net355 vssd1 vssd1 vccd1
+ vccd1 _06850_ sky130_fd_sc_hd__o2111a_1
XANTENNA__08060__C1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11115_ net490 net467 _06615_ net303 net2931 vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__a32o_1
XFILLER_151_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12095_ net562 _06629_ net234 net176 net3036 vssd1 vssd1 vccd1 vccd1 _01515_ sky130_fd_sc_hd__a32o_1
XANTENNA__13487__A1 _05154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15923_ net2257 _02133_ net1184 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[723\]
+ sky130_fd_sc_hd__dfrtp_1
X_11046_ _05960_ _06575_ vssd1 vssd1 vccd1 vccd1 _06582_ sky130_fd_sc_hd__nor2_1
XANTENNA__13279__C_N net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08589__S1 net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11498__B1 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14485__655 clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 net2124 sky130_fd_sc_hd__inv_2
XFILLER_162_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08363__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08902__A2 net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15854_ net2188 _02064_ net1193 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[654\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10170__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15785_ net2119 _01995_ net1055 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[585\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12997_ top.SPI.csx _07425_ _07424_ vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__mux2_1
XFILLER_80_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14526__696 clknet_leaf_151_clk vssd1 vssd1 vccd1 vccd1 net2165 sky130_fd_sc_hd__inv_2
XFILLER_33_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11948_ _06492_ net347 net231 net3205 vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_28_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11670__B1 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11879_ net141 net3183 net189 vssd1 vssd1 vccd1 vccd1 _01684_ sky130_fd_sc_hd__mux2_1
X_16406_ clknet_leaf_55_clk net3839 net1143 vssd1 vssd1 vccd1 vccd1 top.I2C.I2C_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_138_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13618_ net2913 _03037_ net581 vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_138_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09615__B1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13411__B2 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16337_ clknet_leaf_66_clk _02546_ net1165 vssd1 vssd1 vccd1 vccd1 top.CPU.addressnew\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08969__A2 net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11422__B1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13549_ top.CPU.alu.program_counter\[0\] _06462_ net1350 vssd1 vssd1 vccd1 vccd1
+ _02996_ sky130_fd_sc_hd__mux2_1
XFILLER_158_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16268_ clknet_leaf_45_clk _02478_ net1138 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.toreg\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_127_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15219_ net1553 _01429_ net1175 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_145_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16199_ net2533 _02409_ net1198 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[999\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12922__A0 top.CPU.alu.program_counter\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07929__B1 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10528__A2 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10932__C net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08051__C1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07972_ _03610_ vssd1 vssd1 vccd1 vccd1 _03611_ sky130_fd_sc_hd__inv_2
X_13887__57 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 net1526 sky130_fd_sc_hd__inv_2
X_09711_ top.CPU.registers.data\[697\] top.CPU.registers.data\[665\] net1001 vssd1
+ vssd1 vccd1 vccd1 _05350_ sky130_fd_sc_hd__mux2_1
XANTENNA__11489__B1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08354__B1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09642_ _04603_ _05280_ vssd1 vssd1 vccd1 vccd1 _05281_ sky130_fd_sc_hd__nor2_1
XFILLER_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09573_ net676 _05211_ _05210_ net902 vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__o211a_1
XFILLER_24_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout264_A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12989__B1 _07418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09303__C1 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08524_ top.CPU.registers.data\[912\] net1291 net1010 top.CPU.registers.data\[944\]
+ net907 vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__a221o_1
XANTENNA__08845__S net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08455_ net880 _04090_ _04092_ vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__o21a_1
XANTENNA__11661__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07865__C1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10676__A net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout431_A net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1173_A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout529_A net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08386_ top.CPU.registers.data\[434\] top.CPU.registers.data\[402\] net982 vssd1
+ vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__mux2_1
XANTENNA__08409__A1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13402__A1 net1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12205__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07880__A2 net1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11413__B1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout317_X net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15965__RESET_B net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08290__C1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09007_ top.CPU.registers.data\[425\] top.CPU.registers.data\[393\] top.CPU.registers.data\[297\]
+ top.CPU.registers.data\[265\] net965 net1280 vssd1 vssd1 vccd1 vccd1 _04646_ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout1226_X net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14172__342 clknet_leaf_139_clk vssd1 vssd1 vccd1 vccd1 net1811 sky130_fd_sc_hd__inv_2
XANTENNA_fanout686_X net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14871__1041 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 net2510 sky130_fd_sc_hd__inv_2
XFILLER_160_783 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13469__A1 net1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14469__639 clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 net2108 sky130_fd_sc_hd__inv_2
XFILLER_116_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout530 net532 vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__clkbuf_4
Xfanout541 _06524_ vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__buf_4
X_09909_ _05195_ _05547_ vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__nand2_1
Xfanout552 _03172_ vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__clkbuf_4
Xfanout563 net564 vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__buf_4
Xfanout574 net575 vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__buf_4
XANTENNA_fanout853_X net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout585 net586 vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__buf_1
XANTENNA__09542__C1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14213__383 clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 net1852 sky130_fd_sc_hd__inv_2
X_12920_ _07361_ _07362_ vssd1 vssd1 vccd1 vccd1 _07363_ sky130_fd_sc_hd__nor2_1
XANTENNA__13227__A _02782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout596 net598 vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__buf_2
XANTENNA__07699__A2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12851_ _07300_ _07297_ net126 vssd1 vssd1 vccd1 vccd1 _07301_ sky130_fd_sc_hd__mux2_1
XFILLER_92_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11970__A net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11802_ net136 net3495 net157 vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__mux2_1
XFILLER_14_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15570_ net1904 _01780_ net1101 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[370\]
+ sky130_fd_sc_hd__dfrtp_1
X_12782_ _07234_ _07236_ vssd1 vssd1 vccd1 vccd1 _07238_ sky130_fd_sc_hd__and2_1
XANTENNA__11247__A3 _06678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09440__A net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11652__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11733_ net135 net539 net500 net194 net2754 vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__a32o_1
XANTENNA__08743__S1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11664_ net468 _06474_ net240 net167 net3080 vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_172_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13403_ top.I2C.data_out\[26\] net555 _02919_ vssd1 vssd1 vccd1 vccd1 _02920_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_172_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10615_ _05281_ net370 vssd1 vssd1 vccd1 vccd1 _06234_ sky130_fd_sc_hd__nor2_1
XANTENNA__11404__B1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09073__A1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11595_ net457 net233 vssd1 vssd1 vccd1 vccd1 _06754_ sky130_fd_sc_hd__nand2_1
X_16122_ net2456 _02332_ net1251 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[922\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_155_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13334_ net888 _02869_ vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__and2_1
XFILLER_6_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10546_ net550 _04260_ net507 _04256_ vssd1 vssd1 vccd1 vccd1 _06169_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08820__A1 _03342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16053_ net2387 _02263_ net1211 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[853\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_143_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13265_ net3927 _02814_ _02817_ net1053 vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_94_Left_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10477_ _06087_ _06102_ vssd1 vssd1 vccd1 vccd1 _06103_ sky130_fd_sc_hd__and2_1
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15004_ clknet_leaf_97_clk _01249_ net1254 vssd1 vssd1 vccd1 vccd1 top.SPI.parameters\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12216_ top.CPU.registers.data\[43\] net645 vssd1 vssd1 vccd1 vccd1 _06875_ sky130_fd_sc_hd__or2_1
XFILLER_155_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13196_ net36 top.I2C.initiate_read_bit vssd1 vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__nand2b_2
XFILLER_155_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09781__C1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12740__S net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12147_ _06497_ _06749_ _06841_ net172 net3768 vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__a32o_1
XFILLER_110_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09128__A2 net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11864__B _03180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12078_ top.CPU.registers.data\[114\] net649 vssd1 vssd1 vccd1 vccd1 _06808_ sky130_fd_sc_hd__or2_1
XFILLER_110_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09533__C1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11029_ net513 net438 net130 net543 vssd1 vssd1 vccd1 vccd1 _06573_ sky130_fd_sc_hd__and4_1
X_15906_ net2240 _02116_ net1173 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[706\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08887__A1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11891__A0 _06354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15837_ net2171 _02047_ net1114 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[637\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_92_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15125__Q top.CPU.done vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08639__A1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08665__S net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15768_ net2102 _01978_ net1102 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[568\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10446__A1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09350__A net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11643__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07847__C1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15699_ net2033 _01909_ net1178 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[499\]
+ sky130_fd_sc_hd__dfrtp_1
X_08240_ top.CPU.registers.data\[822\] top.CPU.registers.data\[790\] net829 vssd1
+ vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__mux2_1
XANTENNA__10997__A2 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12199__A1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08171_ net695 _03805_ _03806_ _03809_ vssd1 vssd1 vccd1 vccd1 _03810_ sky130_fd_sc_hd__a31o_1
XFILLER_174_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09496__S net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08272__C1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10943__B _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput100 net100 vssd1 vssd1 vccd1 vccd1 SEL_O[0] sky130_fd_sc_hd__buf_2
XFILLER_173_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14156__326 clknet_leaf_194_clk vssd1 vssd1 vccd1 vccd1 net1795 sky130_fd_sc_hd__inv_2
Xoutput111 net111 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_58_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11120__A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09367__A2 net1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08024__C1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10382__B1 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1019_A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13318__Y _02858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07955_ net744 _03589_ _03590_ net694 vssd1 vssd1 vccd1 vccd1 _03594_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_71_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout479_A net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09524__C1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07886_ net801 _03524_ _03518_ net642 vssd1 vssd1 vccd1 vccd1 _03525_ sky130_fd_sc_hd__a211o_1
XFILLER_95_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10685__A1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09625_ top.CPU.registers.data_out_r1_prev\[0\] net877 vssd1 vssd1 vccd1 vccd1 _05264_
+ sky130_fd_sc_hd__or2_1
XANTENNA__11882__A0 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout267_X net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout646_A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1290_A net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1388_A net1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09556_ net381 _05192_ vssd1 vssd1 vccd1 vccd1 _05195_ sky130_fd_sc_hd__xnor2_2
XANTENNA__13623__A1 _05767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08507_ top.CPU.registers.data\[656\] net1322 net853 top.CPU.registers.data\[688\]
+ net721 vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__a221o_1
XANTENNA__11634__B1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09487_ _05125_ vssd1 vssd1 vccd1 vccd1 _05126_ sky130_fd_sc_hd__inv_2
XFILLER_24_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout813_A _03204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout434_X net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10988__A2 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08438_ top.CPU.registers.data\[753\] net1393 net825 top.CPU.registers.data\[721\]
+ net725 vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__a221o_1
XANTENNA__07853__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13387__A0 net1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09055__A1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout601_X net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08369_ top.CPU.registers.data\[434\] top.CPU.registers.data\[402\] net818 vssd1
+ vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__mux2_1
X_10400_ _03789_ _05971_ vssd1 vssd1 vccd1 vccd1 _06029_ sky130_fd_sc_hd__nor2_1
XANTENNA__13510__A _04323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08263__C1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11380_ _06495_ net279 net272 net3267 vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_150_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08604__A net1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10331_ net573 net515 _05962_ vssd1 vssd1 vccd1 vccd1 _05963_ sky130_fd_sc_hd__and3_1
XFILLER_127_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13050_ net3115 _07450_ net895 vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__mux2_1
X_10262_ net399 _05895_ vssd1 vssd1 vccd1 vccd1 _05896_ sky130_fd_sc_hd__nor2_1
XANTENNA__09358__A2 net1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout970_X net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13656__S net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08566__B1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12001_ _06571_ net351 net183 net2809 vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__a22o_1
XFILLER_133_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10193_ _05758_ _05828_ vssd1 vssd1 vccd1 vccd1 _05829_ sky130_fd_sc_hd__nor2_1
XANTENNA__10373__B1 _05754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1303 net1304 vssd1 vssd1 vccd1 vccd1 net1303 sky130_fd_sc_hd__clkbuf_4
Xfanout1314 net1315 vssd1 vssd1 vccd1 vccd1 net1314 sky130_fd_sc_hd__clkbuf_4
Xfanout1325 net1327 vssd1 vssd1 vccd1 vccd1 net1325 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10912__A2 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09435__A net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1336 net1337 vssd1 vssd1 vccd1 vccd1 net1336 sky130_fd_sc_hd__clkbuf_4
Xfanout1347 net67 vssd1 vssd1 vccd1 vccd1 net1347 sky130_fd_sc_hd__clkbuf_2
Xfanout1358 top.SPI.state\[2\] vssd1 vssd1 vccd1 vccd1 net1358 sky130_fd_sc_hd__clkbuf_4
Xfanout360 net365 vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__buf_4
XFILLER_94_829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout371 _05518_ vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__buf_2
Xfanout1369 net1370 vssd1 vssd1 vccd1 vccd1 net1369 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout382 net383 vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__clkbuf_2
XFILLER_47_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout393 _05090_ vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10125__B1 _05762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12903_ _07345_ _07346_ vssd1 vssd1 vccd1 vccd1 _07347_ sky130_fd_sc_hd__nor2_1
XANTENNA__09722__X _05361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07541__A1 top.CPU.control_unit.instruction\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_28_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15622_ net1956 _01832_ net1080 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[422\]
+ sky130_fd_sc_hd__dfrtp_1
X_12834_ _07275_ _07280_ vssd1 vssd1 vccd1 vccd1 _07285_ sky130_fd_sc_hd__nor2_1
XANTENNA__08485__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11625__A0 _06428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15553_ net1887 _01763_ net1225 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[353\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07829__C1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12765_ top.CPU.alu.program_counter\[12\] _07222_ net1361 vssd1 vssd1 vccd1 vccd1
+ _01175_ sky130_fd_sc_hd__mux2_1
XANTENNA__08097__A2 net1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09294__B2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14597__767 clknet_leaf_110_clk vssd1 vssd1 vccd1 vccd1 net2236 sky130_fd_sc_hd__inv_2
X_11716_ _06554_ net196 net420 net3321 vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__a22o_1
X_15484_ net1818 _01694_ net1234 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[284\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07844__A2 net1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12696_ _07158_ _07159_ vssd1 vssd1 vccd1 vccd1 _07160_ sky130_fd_sc_hd__xnor2_1
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11647_ _06193_ net200 net425 net3358 vssd1 vssd1 vccd1 vccd1 _01904_ sky130_fd_sc_hd__a22o_1
Xinput13 DAT_I[1] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput24 DAT_I[2] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
Xinput35 gpio_in[0] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08254__C1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11578_ net2819 net246 _06746_ net478 vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__a22o_1
XFILLER_128_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16105_ net2439 _02315_ net1060 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[905\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_171_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13317_ top.I2C.data_out\[3\] net553 _02856_ vssd1 vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__a21oi_1
Xhold808 top.CPU.registers.data\[706\] vssd1 vssd1 vccd1 vccd1 net3365 sky130_fd_sc_hd__dlygate4sd3_1
X_10529_ _04469_ _05284_ vssd1 vssd1 vccd1 vccd1 _06152_ sky130_fd_sc_hd__or2_1
Xhold819 top.CPU.registers.data\[256\] vssd1 vssd1 vccd1 vccd1 net3376 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_172_Right_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16036_ net2370 _02246_ net1185 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[836\]
+ sky130_fd_sc_hd__dfrtp_1
X_13248_ net3803 _02805_ _02808_ _02803_ vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__a22o_1
XFILLER_170_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08557__B1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13179_ top.I2C.I2C_state\[23\] top.I2C.I2C_state\[2\] _06911_ top.I2C.which_data_address\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__o22a_1
XANTENNA__10364__B1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13857__27 clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 net1496 sky130_fd_sc_hd__inv_2
XANTENNA__08309__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_194_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07740_ top.CPU.registers.data\[574\] top.CPU.registers.data\[542\] net833 vssd1
+ vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__mux2_1
XFILLER_42_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_74_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07671_ _03291_ _03309_ vssd1 vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__nor2_4
XANTENNA__10003__B _05616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10778__X _06390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14541__711 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 net2180 sky130_fd_sc_hd__inv_2
XFILLER_93_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09410_ top.CPU.registers.data\[803\] top.CPU.registers.data\[771\] net828 vssd1
+ vssd1 vccd1 vccd1 _05049_ sky130_fd_sc_hd__mux2_1
XANTENNA__13605__A1 _06008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10938__B _06428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11616__A0 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09341_ top.CPU.registers.data\[228\] net1391 net829 top.CPU.registers.data\[196\]
+ net726 vssd1 vssd1 vccd1 vccd1 _04980_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_89_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14870__1040 clknet_leaf_181_clk vssd1 vssd1 vccd1 vccd1 net2509 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09272_ net928 _04902_ _04904_ net605 vssd1 vssd1 vccd1 vccd1 _04911_ sky130_fd_sc_hd__a31o_1
XFILLER_20_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07835__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13369__A0 top.CPU.control_unit.instruction\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_21_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_132_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08223_ top.CPU.registers.data\[54\] top.CPU.registers.data\[22\] net836 vssd1 vssd1
+ vccd1 vccd1 _03862_ sky130_fd_sc_hd__mux2_1
XANTENNA__09037__A1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout227_A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08154_ top.CPU.registers.data\[87\] net1325 net856 top.CPU.registers.data\[119\]
+ net773 vssd1 vssd1 vccd1 vccd1 _03793_ sky130_fd_sc_hd__a221o_1
XANTENNA__12041__B1 _06781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_12_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11395__A2 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10165__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08085_ top.CPU.alu.program_counter\[21\] net1034 vssd1 vssd1 vccd1 vccd1 _03724_
+ sky130_fd_sc_hd__nor2_1
XFILLER_146_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08260__A2 net1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1136_A net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_147_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout596_A net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13476__S net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09745__C1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_27_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10355__B1 _05742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1303_A net1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09760__A2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08987_ top.CPU.registers.data\[809\] top.CPU.registers.data\[777\] net805 vssd1
+ vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout763_A net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_5_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_5_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_57_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07938_ _03575_ _03576_ net453 vssd1 vssd1 vccd1 vccd1 _03577_ sky130_fd_sc_hd__mux2_1
XFILLER_169_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11855__B1 net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11009__B net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout551_X net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout930_A net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07869_ _03492_ _03507_ vssd1 vssd1 vccd1 vccd1 _03508_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_108_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1293_X net1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14284__454 clknet_leaf_195_clk vssd1 vssd1 vccd1 vccd1 net1923 sky130_fd_sc_hd__inv_2
XANTENNA__08720__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout649_X net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09608_ net787 _05236_ _05237_ net715 vssd1 vssd1 vccd1 vccd1 _05247_ sky130_fd_sc_hd__o211a_1
X_13871__41 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 net1510 sky130_fd_sc_hd__inv_2
X_10880_ net495 net469 _06481_ net223 net2939 vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__a32o_1
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11607__A0 _06056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09539_ net802 _05177_ _05176_ net756 vssd1 vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__o211a_1
XANTENNA__09276__A1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout816_X net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_159_Left_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11025__A _06447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12550_ top.CPU.handler.state\[5\] _07053_ _07054_ _07058_ vssd1 vssd1 vccd1 vccd1
+ _00021_ sky130_fd_sc_hd__a31o_1
X_14325__495 clknet_leaf_173_clk vssd1 vssd1 vccd1 vccd1 net1964 sky130_fd_sc_hd__inv_2
XFILLER_106_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11501_ net480 net472 _06634_ net254 net2947 vssd1 vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__a32o_1
X_12481_ _06977_ _06989_ _06976_ vssd1 vssd1 vccd1 vccd1 _06990_ sky130_fd_sc_hd__o21ba_1
XANTENNA__10864__A net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12032__A0 _06149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08236__C1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11432_ net3479 net265 _06718_ net487 vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__a22o_1
XFILLER_22_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_886 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11386__A2 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08787__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10075__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11363_ net457 _06468_ _06603_ vssd1 vssd1 vccd1 vccd1 _06714_ sky130_fd_sc_hd__or3_4
XANTENNA_hold975_A top.CPU.data_out\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10594__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13102_ _02713_ _02714_ _02715_ _02712_ net4011 vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__a32o_1
XFILLER_4_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10314_ _05821_ _05837_ net387 vssd1 vssd1 vccd1 vccd1 _05946_ sky130_fd_sc_hd__mux2_1
X_11294_ net3499 net289 net359 _05847_ vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__a22o_1
XANTENNA__12335__A1 _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_168_Left_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13239__X _02803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13033_ top.SPI.parameters\[18\] top.SPI.paroutput\[10\] net1355 vssd1 vssd1 vccd1
+ vccd1 _07442_ sky130_fd_sc_hd__mux2_1
XANTENNA__11695__A net1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_167_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10245_ net1406 net577 net517 net135 vssd1 vssd1 vccd1 vccd1 _05880_ sky130_fd_sc_hd__and4_1
XANTENNA__09200__A1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1100 net1109 vssd1 vssd1 vccd1 vccd1 net1100 sky130_fd_sc_hd__buf_2
Xfanout1111 net1277 vssd1 vssd1 vccd1 vccd1 net1111 sky130_fd_sc_hd__buf_2
X_10176_ _03581_ _05506_ _05508_ vssd1 vssd1 vccd1 vccd1 _05812_ sky130_fd_sc_hd__nand3_1
XFILLER_152_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1122 net1127 vssd1 vssd1 vccd1 vccd1 net1122 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09751__A2 net1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1133 net1136 vssd1 vssd1 vccd1 vccd1 net1133 sky130_fd_sc_hd__clkbuf_4
XFILLER_26_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1144 net1145 vssd1 vssd1 vccd1 vccd1 net1144 sky130_fd_sc_hd__clkbuf_4
XFILLER_94_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07762__A1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1155 net1157 vssd1 vssd1 vccd1 vccd1 net1155 sky130_fd_sc_hd__clkbuf_2
Xfanout1166 net1169 vssd1 vssd1 vccd1 vccd1 net1166 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10104__A net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14984_ clknet_leaf_98_clk _01229_ net1256 vssd1 vssd1 vccd1 vccd1 top.SPI.paroutput\[23\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1177 net1179 vssd1 vssd1 vccd1 vccd1 net1177 sky130_fd_sc_hd__clkbuf_4
Xfanout1188 net1205 vssd1 vssd1 vccd1 vccd1 net1188 sky130_fd_sc_hd__clkbuf_2
Xfanout190 net191 vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__buf_6
Xfanout1199 net1200 vssd1 vssd1 vccd1 vccd1 net1199 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11846__B1 net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09503__A2 net1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11310__A2 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13415__A net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload5_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15605_ net1939 _01815_ net1216 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[405\]
+ sky130_fd_sc_hd__dfrtp_1
X_12817_ top.CPU.alu.program_counter\[17\] _07260_ vssd1 vssd1 vccd1 vccd1 _07270_
+ sky130_fd_sc_hd__and2_1
XFILLER_50_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13797_ top.CPU.handler.readout _07054_ _03045_ vssd1 vssd1 vccd1 vccd1 _03096_ sky130_fd_sc_hd__a21boi_4
X_15536_ net1870 _01746_ net1108 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[336\]
+ sky130_fd_sc_hd__dfrtp_1
X_12748_ _07205_ _07206_ vssd1 vssd1 vccd1 vccd1 _07207_ sky130_fd_sc_hd__xor2_1
XANTENNA__08475__C1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11074__B2 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11613__A3 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15467_ net1801 _01677_ net1058 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[267\]
+ sky130_fd_sc_hd__dfrtp_1
X_12679_ net125 _07144_ vssd1 vssd1 vccd1 vccd1 _07145_ sky130_fd_sc_hd__or2_1
XANTENNA__08490__A2 net1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15398_ net1732 _01608_ net1072 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[198\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11377__A2 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08778__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_834 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwire591 _02964_ vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__buf_2
Xhold605 top.CPU.registers.data\[625\] vssd1 vssd1 vccd1 vccd1 net3162 sky130_fd_sc_hd__dlygate4sd3_1
Xhold616 top.CPU.handler.toreg\[31\] vssd1 vssd1 vccd1 vccd1 net3173 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10585__B1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold627 top.CPU.registers.data\[126\] vssd1 vssd1 vccd1 vccd1 net3184 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09627__X _05266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold638 top.CPU.registers.data\[453\] vssd1 vssd1 vccd1 vccd1 net3195 sky130_fd_sc_hd__dlygate4sd3_1
Xhold649 top.I2C.I2C_state\[21\] vssd1 vssd1 vccd1 vccd1 net3206 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12326__A1 _04324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11129__A2 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08910_ net787 _04547_ _04548_ net715 vssd1 vssd1 vccd1 vccd1 _04549_ sky130_fd_sc_hd__o211a_1
X_16019_ net2353 _02229_ net1197 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[819\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11809__S net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09890_ _03647_ _03613_ vssd1 vssd1 vccd1 vccd1 _05529_ sky130_fd_sc_hd__and2b_1
XANTENNA__08250__Y _03889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08841_ top.CPU.registers.data\[811\] top.CPU.registers.data\[779\] net964 vssd1
+ vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__mux2_1
XANTENNA__10888__A1 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09742__A2 net1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_51_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1305 top.SPI.timem\[21\] vssd1 vssd1 vccd1 vccd1 net3862 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1316 top.CPU.registers.data\[623\] vssd1 vssd1 vccd1 vccd1 net3873 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1327 top.SPI.timem\[11\] vssd1 vssd1 vccd1 vccd1 net3884 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08772_ net704 _04401_ _04404_ _04407_ _04410_ vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__o32a_1
Xhold1338 top.CPU.fetch.current_ra\[20\] vssd1 vssd1 vccd1 vccd1 net3895 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1349 top.CPU.handler.toreg\[27\] vssd1 vssd1 vccd1 vccd1 net3906 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14268__438 clknet_leaf_136_clk vssd1 vssd1 vccd1 vccd1 net1907 sky130_fd_sc_hd__inv_2
X_07723_ top.CPU.registers.data\[767\] top.CPU.registers.data\[735\] top.CPU.registers.data\[703\]
+ top.CPU.registers.data\[671\] net992 net957 vssd1 vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__mux4_1
XANTENNA__11837__B1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10949__A net1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11301__A2 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout177_A _06795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07654_ _03259_ _03108_ _03103_ vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__and3b_1
X_14012__182 clknet_leaf_136_clk vssd1 vssd1 vccd1 vccd1 net1651 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14309__479 clknet_leaf_110_clk vssd1 vssd1 vccd1 vccd1 net1948 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07585_ _03211_ net699 _03216_ _03223_ vssd1 vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__a31oi_2
XFILLER_22_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout344_A net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1086_A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09324_ top.CPU.registers.data\[420\] net1392 net829 top.CPU.registers.data\[388\]
+ net696 vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_66_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11065__B2 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07808__A2 net1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_915 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09255_ top.CPU.registers.data\[901\] net1286 net1004 top.CPU.registers.data\[933\]
+ net900 vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__a221o_1
XFILLER_22_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout132_X net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout609_A _03349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08206_ top.CPU.registers.data\[439\] net1014 net912 vssd1 vssd1 vccd1 vccd1 _03845_
+ sky130_fd_sc_hd__a21o_1
XFILLER_119_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12014__B1 net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09186_ net790 _04818_ _04819_ vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__and3_1
XANTENNA__08769__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11368__A2 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08137_ net620 _03773_ _03774_ _03775_ vssd1 vssd1 vccd1 vccd1 _03776_ sky130_fd_sc_hd__a31o_1
XFILLER_134_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09430__A1 net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08068_ top.CPU.registers.data\[404\] net979 vssd1 vssd1 vccd1 vccd1 _03707_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout880_A _03198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12317__A1 _03854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09718__C1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout978_A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14710__880 clknet_leaf_181_clk vssd1 vssd1 vccd1 vccd1 net2349 sky130_fd_sc_hd__inv_2
XANTENNA_fanout1306_X net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10030_ _03311_ _03323_ _03326_ vssd1 vssd1 vccd1 vccd1 _05669_ sky130_fd_sc_hd__a21oi_2
XANTENNA__09733__A2 net1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout766_X net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_162_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13506__Y _02973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11828__B1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11981_ _06538_ net348 net182 net2707 vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__a22o_1
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout933_X net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10859__A _03170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13720_ _03066_ _03067_ vssd1 vssd1 vccd1 vccd1 _02629_ sky130_fd_sc_hd__nor2_1
XANTENNA__10211__X _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10932_ net439 _06373_ net435 vssd1 vssd1 vccd1 vccd1 _06513_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_123_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16319__Q top.CPU.data_out\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13651_ net4022 _07324_ net663 vssd1 vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__mux2_1
X_10863_ top.CPU.registers.data\[991\] net223 vssd1 vssd1 vccd1 vccd1 _06470_ sky130_fd_sc_hd__and2_1
XFILLER_140_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12602_ net1354 top.SPI.state\[3\] vssd1 vssd1 vccd1 vccd1 top.SPI.nextwrx sky130_fd_sc_hd__and2_1
X_16370_ clknet_leaf_70_clk _02579_ net1169 vssd1 vssd1 vccd1 vccd1 top.CPU.fetch.current_ra\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13582_ top.CPU.alu.program_counter\[13\] _06210_ net1352 vssd1 vssd1 vccd1 vccd1
+ _03016_ sky130_fd_sc_hd__mux2_1
XANTENNA__11056__B2 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08457__C1 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10794_ net548 _06402_ vssd1 vssd1 vccd1 vccd1 _06405_ sky130_fd_sc_hd__or2_1
X_15321_ net1655 _01531_ net1203 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[121\]
+ sky130_fd_sc_hd__dfrtp_1
X_12533_ _05548_ _05601_ vssd1 vssd1 vccd1 vccd1 _07042_ sky130_fd_sc_hd__nor2_1
XFILLER_9_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15252_ net1586 _01462_ net1082 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[52\]
+ sky130_fd_sc_hd__dfrtp_1
X_12464_ _05330_ _05361_ _05466_ _05498_ _06971_ vssd1 vssd1 vccd1 vccd1 _06973_ sky130_fd_sc_hd__o221a_1
XFILLER_138_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11359__A2 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11415_ _06550_ net278 net268 net2897 vssd1 vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_169_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15183_ net1520 _01393_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r1_prev\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_12395_ top.SPI.register\[2\] net599 vssd1 vssd1 vccd1 vccd1 _06933_ sky130_fd_sc_hd__nand2_1
XANTENNA__10567__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08224__A2 net1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11346_ net3669 net286 net278 _06151_ vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__a22o_1
XFILLER_99_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12308__A1 _05265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11277_ net517 _06567_ vssd1 vssd1 vccd1 vccd1 _06696_ sky130_fd_sc_hd__nor2_2
XFILLER_4_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13016_ net2762 _07433_ net895 vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__mux2_1
X_10228_ _03315_ _05435_ _05862_ net410 _05857_ vssd1 vssd1 vccd1 vccd1 _05863_ sky130_fd_sc_hd__a221o_1
XFILLER_121_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11531__A2 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08932__B1 net1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2 top.mmio.s1 vssd1 vssd1 vccd1 vccd1 net2559 sky130_fd_sc_hd__dlygate4sd3_1
X_10159_ _03477_ net507 net505 _05510_ vssd1 vssd1 vccd1 vccd1 _05796_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__13808__B2 top.CPU.data_out\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11872__B net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14967_ clknet_leaf_96_clk net3051 net1254 vssd1 vssd1 vccd1 vccd1 top.SPI.paroutput\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12087__A3 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08696__C1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08160__A1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16229__Q top.CPU.control_unit.instruction\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09769__S net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08448__C1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11047__B2 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08999__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15519_ net1853 _01729_ net1223 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[319\]
+ sky130_fd_sc_hd__dfrtp_1
X_16499_ clknet_leaf_41_clk _02661_ net1115 vssd1 vssd1 vccd1 vccd1 top.mmio.mem_data_i\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08463__A2 net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14653__823 clknet_leaf_133_clk vssd1 vssd1 vccd1 vccd1 net2292 sky130_fd_sc_hd__inv_2
X_09040_ net785 _04672_ _04673_ vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__and3_1
XFILLER_129_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11112__B net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09412__A1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold402 net79 vssd1 vssd1 vccd1 vccd1 net2959 sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 top.CPU.registers.data\[919\] vssd1 vssd1 vccd1 vccd1 net2970 sky130_fd_sc_hd__dlygate4sd3_1
Xhold424 top.CPU.registers.data\[781\] vssd1 vssd1 vccd1 vccd1 net2981 sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 net40 vssd1 vssd1 vccd1 vccd1 net2992 sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 top.CPU.registers.data\[388\] vssd1 vssd1 vccd1 vccd1 net3003 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10951__B net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07974__A1 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold457 net90 vssd1 vssd1 vccd1 vccd1 net3014 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold468 top.CPU.registers.data\[391\] vssd1 vssd1 vccd1 vccd1 net3025 sky130_fd_sc_hd__dlygate4sd3_1
X_09942_ _03755_ _03785_ vssd1 vssd1 vccd1 vccd1 _05581_ sky130_fd_sc_hd__and2_1
XFILLER_89_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10443__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold479 top.CPU.registers.data\[105\] vssd1 vssd1 vccd1 vccd1 net3036 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout904 net909 vssd1 vssd1 vccd1 vccd1 net904 sky130_fd_sc_hd__clkbuf_4
Xfanout915 net925 vssd1 vssd1 vccd1 vccd1 net915 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09176__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout926 net949 vssd1 vssd1 vccd1 vccd1 net926 sky130_fd_sc_hd__clkbuf_4
X_09873_ _03511_ _05510_ vssd1 vssd1 vccd1 vccd1 _05512_ sky130_fd_sc_hd__and2b_1
XFILLER_112_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout937 net938 vssd1 vssd1 vccd1 vccd1 net937 sky130_fd_sc_hd__clkbuf_2
Xfanout948 net949 vssd1 vssd1 vccd1 vccd1 net948 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07726__A1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout294_A _06662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11522__A2 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout959 net961 vssd1 vssd1 vccd1 vccd1 net959 sky130_fd_sc_hd__clkbuf_4
X_08824_ _04462_ vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__inv_2
Xhold1102 top.CPU.registers.data\[987\] vssd1 vssd1 vccd1 vccd1 net3659 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_86_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1113 top.CPU.registers.data\[867\] vssd1 vssd1 vccd1 vccd1 net3670 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1124 top.CPU.registers.data\[974\] vssd1 vssd1 vccd1 vccd1 net3681 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1001_A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1135 net72 vssd1 vssd1 vccd1 vccd1 net3692 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07752__S net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1146 top.CPU.registers.data\[637\] vssd1 vssd1 vccd1 vccd1 net3703 sky130_fd_sc_hd__dlygate4sd3_1
X_08755_ _04363_ _04393_ vssd1 vssd1 vccd1 vccd1 _04394_ sky130_fd_sc_hd__nor2_1
Xhold1157 top.CPU.registers.data\[963\] vssd1 vssd1 vccd1 vccd1 net3714 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09479__A1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout461_A net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1168 top.CPU.registers.data\[929\] vssd1 vssd1 vccd1 vccd1 net3725 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1179 top.CPU.handler.toreg\[7\] vssd1 vssd1 vccd1 vccd1 net3736 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout559_A net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07706_ top.CPU.registers.data\[799\] net1030 net959 _03344_ vssd1 vssd1 vccd1 vccd1
+ _03345_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_68_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08686_ top.CPU.control_unit.instruction\[14\] _03160_ _03985_ vssd1 vssd1 vccd1
+ vccd1 _04325_ sky130_fd_sc_hd__o21a_2
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07637_ _03108_ _03177_ _03259_ _03263_ vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__and4_1
X_13841__11 clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 net1480 sky130_fd_sc_hd__inv_2
XANTENNA__12894__A top.CPU.alu.program_counter\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1370_A net1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout726_A net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout347_X net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12235__B1 _03185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11038__B2 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07568_ top.CPU.registers.data\[703\] top.CPU.registers.data\[671\] net829 vssd1
+ vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__mux2_1
XANTENNA__09100__B1 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09307_ net940 _04924_ _04945_ net957 vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_81_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13502__B _02967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07499_ top.SPI.percount\[3\] vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__inv_2
XANTENNA__08454__A2 _04090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout514_X net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14396__566 clknet_leaf_137_clk vssd1 vssd1 vccd1 vccd1 net2035 sky130_fd_sc_hd__inv_2
X_09238_ top.CPU.registers.data\[837\] net1310 net841 top.CPU.registers.data\[869\]
+ net737 vssd1 vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__a221o_1
XFILLER_139_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12118__B net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08206__A2 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09169_ net790 _04806_ _04807_ net692 vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__o211a_1
XFILLER_163_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10549__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11200_ net1401 net480 _06657_ net297 net2901 vssd1 vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__a32o_1
XFILLER_134_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08611__C1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12180_ net567 _06664_ net240 net170 net2664 vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout883_X net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08612__A net1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07965__A1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11131_ net482 net456 _06623_ net301 net3739 vssd1 vssd1 vccd1 vccd1 _02287_ sky130_fd_sc_hd__a32o_1
Xhold980 top.CPU.registers.data\[883\] vssd1 vssd1 vccd1 vccd1 net3537 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_164_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold991 top.CPU.registers.data\[862\] vssd1 vssd1 vccd1 vccd1 net3548 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09706__A2 net1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11062_ _06190_ _06575_ vssd1 vssd1 vccd1 vccd1 _06588_ sky130_fd_sc_hd__nor2_1
XFILLER_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07717__A1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08914__B1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11513__A2 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10013_ net384 _05651_ vssd1 vssd1 vccd1 vccd1 _05652_ sky130_fd_sc_hd__nand2_1
XFILLER_49_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15870_ net2204 _02080_ net1239 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[670\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_160_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input22_A DAT_I[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_73 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11964_ _06513_ net342 net229 net3300 vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__a22o_1
XANTENNA__08678__C1 net1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11816__A3 net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08142__A1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13703_ net3844 _03054_ vssd1 vssd1 vccd1 vccd1 _03057_ sky130_fd_sc_hd__nor2_1
X_10915_ net660 _06230_ net435 vssd1 vssd1 vccd1 vccd1 _06503_ sky130_fd_sc_hd__and3_1
XFILLER_72_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11895_ _06428_ net3263 net188 vssd1 vssd1 vccd1 vccd1 _01668_ sky130_fd_sc_hd__mux2_1
X_14340__510 clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 net1979 sky130_fd_sc_hd__inv_2
X_16422_ clknet_leaf_55_clk _00004_ net1143 vssd1 vssd1 vccd1 vccd1 top.I2C.I2C_state\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13634_ net3262 _07162_ net664 vssd1 vssd1 vccd1 vccd1 _02568_ sky130_fd_sc_hd__mux2_1
X_10846_ net508 _06453_ _06452_ vssd1 vssd1 vccd1 vccd1 _06454_ sky130_fd_sc_hd__a21o_1
XANTENNA__08493__S net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14637__807 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 net2276 sky130_fd_sc_hd__inv_2
XFILLER_158_723 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16353_ clknet_leaf_72_clk _02562_ net1153 vssd1 vssd1 vccd1 vccd1 top.CPU.fetch.current_ra\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13565_ top.CPU.addressnew\[6\] _03005_ net580 vssd1 vssd1 vccd1 vccd1 _02536_ sky130_fd_sc_hd__mux2_1
X_10777_ _06384_ _06386_ _06388_ vssd1 vssd1 vccd1 vccd1 _06389_ sky130_fd_sc_hd__or3_2
XFILLER_9_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15304_ net1638 _01514_ net1087 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[104\]
+ sky130_fd_sc_hd__dfrtp_1
X_12516_ _07016_ _07021_ _07022_ _07024_ vssd1 vssd1 vccd1 vccd1 _07025_ sky130_fd_sc_hd__a31oi_1
XFILLER_8_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16284_ clknet_leaf_62_clk _02494_ net1161 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.toreg\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16448__RESET_B net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13496_ net1400 net874 _03248_ _02965_ vssd1 vssd1 vccd1 vccd1 _02967_ sky130_fd_sc_hd__a31o_2
XANTENNA__12028__B net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15235_ net1569 _01445_ net1210 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[35\]
+ sky130_fd_sc_hd__dfrtp_1
X_12447_ net1339 top.I2C.output_state\[1\] top.I2C.output_state\[16\] vssd1 vssd1
+ vccd1 vccd1 _06960_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_136_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07837__S net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15166_ net1503 _01376_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r1_prev\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_12378_ _03125_ _06915_ _06916_ vssd1 vssd1 vccd1 vccd1 _00040_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08602__C1 net1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07956__A1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11752__A2 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11329_ _03174_ net570 _06603_ vssd1 vssd1 vccd1 vccd1 _06712_ sky130_fd_sc_hd__or3_4
X_15097_ net1479 _01310_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r2_prev\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11504__A2 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08381__A1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09005__S0 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15999_ net2333 _02209_ net1223 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[799\]
+ sky130_fd_sc_hd__dfrtp_1
X_08540_ top.CPU.registers.data\[560\] top.CPU.registers.data\[528\] net984 vssd1
+ vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__mux2_1
XANTENNA__11268__B2 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11807__A3 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08471_ top.CPU.registers.data\[689\] top.CPU.registers.data\[657\] net995 vssd1
+ vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__mux2_1
XANTENNA__13009__A2 _07429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12217__B1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07892__B1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14083__253 clknet_leaf_114_clk vssd1 vssd1 vccd1 vccd1 net1722 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_63_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10946__B net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10779__B1 _06390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_114_Left_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11440__A1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14124__294 clknet_leaf_188_clk vssd1 vssd1 vccd1 vccd1 net1763 sky130_fd_sc_hd__inv_2
XFILLER_164_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09023_ net452 _04658_ vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__or2_1
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11991__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10962__A _05906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1049_A _03093_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold210 top.CPU.registers.data\[479\] vssd1 vssd1 vccd1 vccd1 net2767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 top.SPI.parameters\[31\] vssd1 vssd1 vccd1 vccd1 net2778 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold232 top.CPU.registers.data\[549\] vssd1 vssd1 vccd1 vccd1 net2789 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08432__A net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold243 top.CPU.addressnew\[29\] vssd1 vssd1 vccd1 vccd1 net2800 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11743__A2 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold254 _02705_ vssd1 vssd1 vccd1 vccd1 net2811 sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 top.CPU.registers.data\[173\] vssd1 vssd1 vccd1 vccd1 net2822 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold276 top.CPU.registers.data\[823\] vssd1 vssd1 vccd1 vccd1 net2833 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold287 top.CPU.registers.data\[30\] vssd1 vssd1 vccd1 vccd1 net2844 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout701 _03213_ vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__buf_4
XFILLER_172_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09925_ _05541_ _05561_ _05563_ vssd1 vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__a21o_2
Xhold298 top.CPU.registers.data\[606\] vssd1 vssd1 vccd1 vccd1 net2855 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout712 _03212_ vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__clkbuf_4
Xfanout723 net724 vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__clkbuf_4
XFILLER_113_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13496__A2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout734 net735 vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13484__S net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_123_Left_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout297_X net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout745 net746 vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__buf_2
XANTENNA_fanout676_A _03336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14781__951 clknet_leaf_134_clk vssd1 vssd1 vccd1 vccd1 net2420 sky130_fd_sc_hd__inv_2
XFILLER_59_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout756 net759 vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_142_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout767 net768 vssd1 vssd1 vccd1 vccd1 net767 sky130_fd_sc_hd__clkbuf_4
X_09856_ net682 _05493_ _05494_ net609 vssd1 vssd1 vccd1 vccd1 _05495_ sky130_fd_sc_hd__a31o_1
XANTENNA__08578__S net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1004_X net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout778 net781 vssd1 vssd1 vccd1 vccd1 net778 sky130_fd_sc_hd__clkbuf_4
Xfanout789 net790 vssd1 vssd1 vccd1 vccd1 net789 sky130_fd_sc_hd__clkbuf_4
XFILLER_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08807_ top.CPU.registers.data\[972\] net1372 net977 top.CPU.registers.data\[1004\]
+ net1364 vssd1 vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__o221a_1
XFILLER_65_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09787_ net680 _05406_ _05407_ vssd1 vssd1 vccd1 vccd1 _05426_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout843_A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout464_X net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07580__C1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08738_ net950 _04373_ net624 vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10202__A net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14822__992 clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 net2461 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_120_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13988__158 clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 net1627 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_83_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11017__B _03170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08669_ net963 _04304_ net625 vssd1 vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__a21o_1
XFILLER_14_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1373_X net1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout729_X net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10700_ _05541_ _05561_ vssd1 vssd1 vccd1 vccd1 _06315_ sky130_fd_sc_hd__or2_1
XFILLER_14_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11680_ net516 _06500_ net200 net165 net3044 vssd1 vssd1 vccd1 vccd1 _01872_ sky130_fd_sc_hd__a32o_1
XANTENNA__07883__B1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10482__A2 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10631_ _05642_ _05872_ _06246_ _06247_ _06249_ vssd1 vssd1 vccd1 vccd1 _06250_ sky130_fd_sc_hd__a221o_2
XTAP_TAPCELL_ROW_157_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09085__C1 top.CPU.control_unit.instruction\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09624__A1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08427__A2 net1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11033__A net1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13350_ top.CPU.control_unit.instruction\[11\] _02881_ net667 vssd1 vssd1 vccd1 vccd1
+ _02445_ sky130_fd_sc_hd__mux2_1
X_10562_ _04328_ net510 _05679_ _04327_ vssd1 vssd1 vccd1 vccd1 _06184_ sky130_fd_sc_hd__o22a_1
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_118_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12301_ net3761 _04764_ net1202 vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__mux2_1
XANTENNA__13659__S net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11982__A2 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13281_ net4007 _02827_ vssd1 vssd1 vccd1 vccd1 _02828_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_153_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10493_ _04123_ net506 _06117_ vssd1 vssd1 vccd1 vccd1 _06118_ sky130_fd_sc_hd__a21o_1
XANTENNA__10872__A net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07650__A3 _03154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15020_ clknet_leaf_98_clk _01265_ net1256 vssd1 vssd1 vccd1 vccd1 top.SPI.parameters\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_12232_ net3842 net653 _06882_ vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__o21a_1
XFILLER_108_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08342__A net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07938__A1 _03576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11734__A2 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11179__S net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12163_ net362 _06737_ _06849_ net174 net3745 vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_9_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11114_ net574 net529 _06035_ vssd1 vssd1 vccd1 vccd1 _06615_ sky130_fd_sc_hd__and3_1
XFILLER_111_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12094_ net3942 net647 _06815_ vssd1 vssd1 vccd1 vccd1 _01516_ sky130_fd_sc_hd__o21a_1
XFILLER_110_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11045_ net3749 net369 _06581_ net319 vssd1 vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__a22o_1
XANTENNA__11498__A1 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15922_ net2256 _02132_ net1101 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[722\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08899__C1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13932__102 clknet_leaf_193_clk vssd1 vssd1 vccd1 vccd1 net1571 sky130_fd_sc_hd__inv_2
XFILLER_49_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15853_ net2187 _02063_ net1077 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[653\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07571__C1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11208__A net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12996_ top.SPI.state\[4\] _07112_ _06917_ vssd1 vssd1 vccd1 vccd1 _07425_ sky130_fd_sc_hd__a21o_1
X_15784_ net2118 _01994_ net1098 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[584\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_80_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14067__237 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 net1706 sky130_fd_sc_hd__inv_2
X_11947_ _06491_ net344 net230 net3509 vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__a22o_1
XANTENNA__08666__A2 net1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11670__A1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11878_ _06084_ net3539 net190 vssd1 vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__mux2_1
XANTENNA__08517__A _04155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16405_ clknet_leaf_64_clk _00076_ net1161 vssd1 vssd1 vccd1 vccd1 top.wm.curr_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13617_ top.CPU.alu.program_counter\[27\] _05876_ net1351 vssd1 vssd1 vccd1 vccd1
+ _03037_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_138_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10829_ net511 _05548_ _06437_ _05918_ _05753_ vssd1 vssd1 vccd1 vccd1 _06438_ sky130_fd_sc_hd__a32o_1
X_14108__278 clknet_leaf_138_clk vssd1 vssd1 vccd1 vccd1 net1747 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_138_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16336_ clknet_leaf_66_clk _02545_ net1165 vssd1 vssd1 vccd1 vccd1 top.CPU.addressnew\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13548_ _07056_ _02993_ vssd1 vssd1 vccd1 vccd1 _02995_ sky130_fd_sc_hd__nand2_1
XFILLER_9_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11973__A2 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16267_ clknet_leaf_44_clk _02477_ net1126 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.toreg\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13479_ net1396 net872 _02929_ net419 vssd1 vssd1 vccd1 vccd1 _02961_ sky130_fd_sc_hd__a31o_1
XFILLER_65_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15218_ net1552 _01428_ net1098 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_161_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16198_ net2532 _02408_ net1072 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[998\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16242__Q top.CPU.control_unit.instruction\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11725__A2 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15149_ clknet_leaf_42_clk _01359_ net1118 vssd1 vssd1 vccd1 vccd1 top.I2C.data_out\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10933__B1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14765__935 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 net2404 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_39_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07971_ net641 _03608_ _03609_ vssd1 vssd1 vccd1 vccd1 _03610_ sky130_fd_sc_hd__o21ai_4
XFILLER_45_1030 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11817__S _06762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09710_ top.CPU.registers.data\[569\] top.CPU.registers.data\[537\] net1001 vssd1
+ vssd1 vccd1 vccd1 _05349_ sky130_fd_sc_hd__mux2_1
XANTENNA__11489__A1 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09000__C1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12502__A _04828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09551__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12150__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09641_ _04732_ _04797_ _05276_ _05279_ _05278_ vssd1 vssd1 vccd1 vccd1 _05280_ sky130_fd_sc_hd__o41a_2
X_14806__976 clknet_leaf_181_clk vssd1 vssd1 vccd1 vccd1 net2445 sky130_fd_sc_hd__inv_2
XANTENNA__10161__A1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11118__A net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09572_ top.CPU.registers.data\[32\] top.CPU.registers.data\[0\] net973 vssd1 vssd1
+ vccd1 vccd1 _05211_ sky130_fd_sc_hd__mux2_1
XANTENNA__08106__A1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12989__A1 top.SPI.busy vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08523_ top.CPU.registers.data\[816\] top.CPU.registers.data\[784\] net984 vssd1
+ vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__mux2_1
XFILLER_70_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout257_A _06728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08454_ _03198_ _04090_ _04092_ vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__o21ai_2
XANTENNA__07602__Y _03241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09606__A1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08385_ net934 _04023_ vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout424_A _06756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1166_A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08814__C1 net1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09082__A2 net1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11964__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08290__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout212_X net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1333_A net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09006_ net617 _04644_ _04639_ _03342_ vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__o211a_1
XFILLER_164_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11177__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout793_A net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11716__A2 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_131_Left_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10924__B1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08593__A1 net1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09790__B1 _03408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout960_A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13469__A2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout520 net522 vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__buf_2
XANTENNA_fanout679_X net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout531 net532 vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__clkbuf_2
XFILLER_116_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout542 net544 vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__buf_2
X_09908_ net372 _05266_ vssd1 vssd1 vccd1 vccd1 _05547_ sky130_fd_sc_hd__or2_1
XANTENNA__13508__A _04390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout553 net554 vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__buf_2
XANTENNA__12677__B1 top.CPU.alu.program_counter\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout564 net569 vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08345__A1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout575 _03171_ vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__buf_4
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12141__A2 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout597 net598 vssd1 vssd1 vccd1 vccd1 net597 sky130_fd_sc_hd__clkbuf_2
X_09839_ top.CPU.registers.data\[570\] top.CPU.registers.data\[538\] net1000 vssd1
+ vssd1 vccd1 vccd1 _05478_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout846_X net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11028__A net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12850_ _07298_ _07299_ vssd1 vssd1 vccd1 vccd1 _07300_ sky130_fd_sc_hd__nor2_1
XANTENNA__09280__X _04919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11801_ net1402 _06647_ net240 net157 net2980 vssd1 vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__a32o_1
XANTENNA__11970__B net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _07218_ _07235_ _07234_ _07223_ vssd1 vssd1 vccd1 vccd1 _07237_ sky130_fd_sc_hd__a211oi_2
XPHY_EDGE_ROW_140_Left_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11462__S net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10455__A2 _06081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11732_ _06579_ net499 net193 net3102 vssd1 vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__a22o_1
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11663_ net520 _06473_ net208 net166 net2767 vssd1 vssd1 vccd1 vccd1 _01889_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_153_Right_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13402_ net1346 top.mmio.mem_data_i\[26\] net598 vssd1 vssd1 vccd1 vccd1 _02919_
+ sky130_fd_sc_hd__o21a_1
XFILLER_174_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_172_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10207__A2 _05824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07608__B1 net1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10614_ net3833 net225 net313 _06233_ vssd1 vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_172_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11594_ net472 _06751_ vssd1 vssd1 vccd1 vccd1 _06753_ sky130_fd_sc_hd__nor2_1
X_16121_ net2455 _02331_ net1245 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[921\]
+ sky130_fd_sc_hd__dfrtp_1
X_13333_ top.I2C.data_out\[7\] net553 _02868_ net596 vssd1 vssd1 vccd1 vccd1 _02869_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11955__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10545_ _04258_ net510 net505 _04259_ vssd1 vssd1 vccd1 vccd1 _06168_ sky130_fd_sc_hd__o22ai_1
XFILLER_127_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12293__S net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_130_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_130_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_133_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16052_ net2386 _02262_ net1112 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[852\]
+ sky130_fd_sc_hd__dfrtp_1
X_13264_ top.I2C.data_out\[4\] net891 _02755_ vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__mux2_1
X_14452__622 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 net2091 sky130_fd_sc_hd__inv_2
X_10476_ net512 _06062_ _06101_ _06100_ vssd1 vssd1 vccd1 vccd1 _06102_ sky130_fd_sc_hd__a31oi_2
XANTENNA__11168__A0 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15003_ clknet_leaf_96_clk _01248_ net1247 vssd1 vssd1 vccd1 vccd1 top.SPI.parameters\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_14749__919 clknet_leaf_134_clk vssd1 vssd1 vccd1 vccd1 net2388 sky130_fd_sc_hd__inv_2
XANTENNA__11707__A2 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12215_ net360 _06744_ _06874_ net168 net3235 vssd1 vssd1 vccd1 vccd1 _01454_ sky130_fd_sc_hd__a32o_1
X_13195_ top.I2C.which_data_address\[0\] top.I2C.which_data_address\[1\] vssd1 vssd1
+ vccd1 vccd1 _02775_ sky130_fd_sc_hd__nand2_1
XANTENNA__10107__A _03822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09230__C1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12146_ top.CPU.registers.data\[79\] net648 vssd1 vssd1 vccd1 vccd1 _06841_ sky130_fd_sc_hd__or2_1
XFILLER_2_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12077_ top.CPU.registers.data\[114\] net177 vssd1 vssd1 vccd1 vccd1 _06807_ sky130_fd_sc_hd__and2_1
XANTENNA__12132__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11028_ net438 net130 net543 vssd1 vssd1 vccd1 vccd1 _06572_ sky130_fd_sc_hd__and3_1
XFILLER_38_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15905_ net2239 _02115_ net1230 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[705\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_197_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_197_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11340__B1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15836_ net2170 _02046_ net1195 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[636\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_66_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09190__X _04829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07703__X _03342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12979_ top.I2C.bit_timer_counter\[5\] _07411_ top.I2C.bit_timer_state\[0\] vssd1
+ vssd1 vccd1 vccd1 _07412_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09836__A1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15767_ net2101 _01977_ net1180 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[567\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07847__B1 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15698_ net2032 _01908_ net1101 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[498\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10851__C1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_120_Right_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09777__S net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08170_ net707 _03807_ _03808_ vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__and3_1
XFILLER_146_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16319_ clknet_leaf_95_clk _02528_ net1260 vssd1 vssd1 vccd1 vccd1 top.CPU.data_out\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13600__B _06054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_121_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_121_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput101 net101 vssd1 vssd1 vccd1 vccd1 SEL_O[1] sky130_fd_sc_hd__buf_2
X_14195__365 clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 net1834 sky130_fd_sc_hd__inv_2
XFILLER_133_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12216__B net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput112 net112 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_58_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08575__A1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15345__RESET_B net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07783__C1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07954_ net793 _03582_ _03583_ net721 vssd1 vssd1 vccd1 vccd1 _03593_ sky130_fd_sc_hd__o211a_1
XFILLER_102_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12123__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09524__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_71_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_188_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_188_clk
+ sky130_fd_sc_hd__clkbuf_8
X_07885_ net712 _03522_ _03523_ _03521_ vssd1 vssd1 vccd1 vccd1 _03524_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout374_A net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09624_ net703 _05261_ _05262_ _05259_ _05260_ vssd1 vssd1 vccd1 vccd1 _05263_ sky130_fd_sc_hd__o32a_1
XFILLER_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07613__X _03252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09555_ net381 _05192_ vssd1 vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__or2_1
XFILLER_71_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09288__C1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout162_X net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout541_A _06524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1283_A net1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08506_ top.CPU.registers.data\[560\] top.CPU.registers.data\[528\] net821 vssd1
+ vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__mux2_1
XANTENNA__07838__B1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09486_ net394 _05123_ vssd1 vssd1 vccd1 vccd1 _05125_ sky130_fd_sc_hd__or2_1
XFILLER_24_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08437_ top.CPU.registers.data\[593\] net1326 net857 top.CPU.registers.data\[625\]
+ net750 vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__a221o_1
XFILLER_12_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout806_A net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout427_X net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1169_X net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08368_ top.CPU.registers.data\[242\] net1389 net818 top.CPU.registers.data\[210\]
+ net769 vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__a221o_1
XANTENNA__10693__Y _06309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11398__B1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11937__A2 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14436__606 clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 net2075 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_115_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13510__B _02966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09460__C1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08299_ net796 _03932_ _03933_ net750 vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_78_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_112_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_112_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_150_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1336_X net1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13139__A1 top.CPU.data_out\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11311__A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10330_ _05697_ _05961_ vssd1 vssd1 vccd1 vccd1 _05962_ sky130_fd_sc_hd__and2_2
XFILLER_125_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout796_X net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10261_ _05720_ _05725_ net387 vssd1 vssd1 vccd1 vccd1 _05895_ sky130_fd_sc_hd__mux2_1
XANTENNA__09212__C1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12000_ _06569_ net347 net180 net2832 vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__a22o_1
XFILLER_79_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10192_ net406 _05827_ vssd1 vssd1 vccd1 vccd1 _05828_ sky130_fd_sc_hd__nor2_1
XANTENNA__08620__A _04225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout963_X net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1304 _03113_ vssd1 vssd1 vccd1 vccd1 net1304 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11570__B1 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1315 net1323 vssd1 vssd1 vccd1 vccd1 net1315 sky130_fd_sc_hd__clkbuf_4
Xfanout1326 net1327 vssd1 vssd1 vccd1 vccd1 net1326 sky130_fd_sc_hd__clkbuf_4
Xfanout1337 net1338 vssd1 vssd1 vccd1 vccd1 net1337 sky130_fd_sc_hd__clkbuf_4
Xfanout1348 net1349 vssd1 vssd1 vccd1 vccd1 net1348 sky130_fd_sc_hd__buf_2
XFILLER_121_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout350 net353 vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__buf_4
Xfanout361 net365 vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__buf_4
XFILLER_143_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1359 net1360 vssd1 vssd1 vccd1 vccd1 net1359 sky130_fd_sc_hd__clkbuf_4
Xfanout372 net373 vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__buf_2
XFILLER_4_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10125__A1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout383 _05157_ vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_179_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_179_clk
+ sky130_fd_sc_hd__clkbuf_8
Xfanout394 net398 vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__buf_2
XANTENNA__11322__B1 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12902_ top.CPU.alu.program_counter\[26\] top.CPU.alu.program_counter\[25\] top.CPU.alu.program_counter\[24\]
+ _07322_ vssd1 vssd1 vccd1 vccd1 _07346_ sky130_fd_sc_hd__and4_1
XFILLER_4_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11873__A1 _05960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08766__S net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07541__A2 net1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13075__A0 top.CPU.data_out\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12833_ top.CPU.alu.program_counter\[19\] _03986_ vssd1 vssd1 vccd1 vccd1 _07284_
+ sky130_fd_sc_hd__xor2_1
X_15621_ net1955 _01831_ net1063 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[421\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_62_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09818__A1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11192__S net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ _07221_ _07220_ net128 vssd1 vssd1 vccd1 vccd1 _07222_ sky130_fd_sc_hd__mux2_1
X_15552_ net1886 _01762_ net1096 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[352\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_174_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10833__C1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11715_ _06552_ net201 net421 net2876 vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__a22o_1
X_15483_ net1817 _01693_ net1214 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[283\]
+ sky130_fd_sc_hd__dfrtp_1
X_12695_ _07148_ _07150_ _07147_ vssd1 vssd1 vccd1 vccd1 _07159_ sky130_fd_sc_hd__a21oi_2
XFILLER_147_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09597__S net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11646_ _06175_ net199 net426 net3430 vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__a22o_1
XANTENNA__09046__A2 net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11389__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput14 DAT_I[20] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11928__A2 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput25 DAT_I[30] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14179__349 clknet_leaf_114_clk vssd1 vssd1 vccd1 vccd1 net1818 sky130_fd_sc_hd__inv_2
Xinput36 gpio_in[1] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_1
XFILLER_128_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11577_ net570 _06688_ vssd1 vssd1 vccd1 vccd1 _06746_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_103_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_103_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_156_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13316_ net1343 top.mmio.mem_data_i\[3\] net596 vssd1 vssd1 vccd1 vccd1 _02856_ sky130_fd_sc_hd__o21a_1
XFILLER_7_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16104_ net2438 _02314_ net1087 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[904\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_128_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10528_ net3723 net228 net314 _06151_ vssd1 vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__a22o_1
XFILLER_170_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold809 top.CPU.registers.data\[904\] vssd1 vssd1 vccd1 vccd1 net3366 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13247_ top.I2C.data_out\[12\] net892 _02755_ vssd1 vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__mux2_1
X_16035_ net2369 _02245_ net1182 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[835\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12889__B1 net1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10459_ net574 net518 net440 net132 vssd1 vssd1 vccd1 vccd1 _06086_ sky130_fd_sc_hd__and4_1
X_13178_ _06913_ _02757_ _02759_ _02756_ net3891 vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__a32o_1
XANTENNA__13419__Y _02932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11561__B1 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12129_ net3746 net173 _06832_ vssd1 vssd1 vccd1 vccd1 _01498_ sky130_fd_sc_hd__a21o_1
XANTENNA__10124__X _05762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12052__A net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12105__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11313__B1 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07670_ _03251_ _03301_ _03160_ _03162_ vssd1 vssd1 vccd1 vccd1 _03309_ sky130_fd_sc_hd__o211ai_4
X_14580__750 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 net2219 sky130_fd_sc_hd__inv_2
XANTENNA__08190__C1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13066__A0 top.CPU.data_out\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15819_ net2153 _02029_ net1058 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[619\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_80_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08248__Y _03887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10938__C net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09340_ top.CPU.registers.data\[68\] net1329 net860 top.CPU.registers.data\[100\]
+ net752 vssd1 vssd1 vccd1 vccd1 _04979_ sky130_fd_sc_hd__a221o_1
XFILLER_34_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14621__791 clknet_leaf_133_clk vssd1 vssd1 vccd1 vccd1 net2260 sky130_fd_sc_hd__inv_2
X_09271_ net672 _04900_ _04901_ net900 vssd1 vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_16_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11830__S net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08222_ top.CPU.registers.data\[374\] top.CPU.registers.data\[342\] top.CPU.registers.data\[310\]
+ top.CPU.registers.data\[278\] net835 net780 vssd1 vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__mux4_1
XFILLER_119_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11919__A2 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09300__S net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08153_ top.CPU.registers.data\[55\] top.CPU.registers.data\[23\] net823 vssd1 vssd1
+ vccd1 vccd1 _03792_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout122_A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09442__C1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10052__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08084_ _03722_ vssd1 vssd1 vccd1 vccd1 _03723_ sky130_fd_sc_hd__inv_2
XFILLER_161_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12661__S net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1031_A net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1129_A net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07755__S net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08548__A1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09745__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10355__B2 _05979_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout491_A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07756__C1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout589_A net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10181__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08986_ net635 _04621_ _04624_ vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__or3_1
XFILLER_103_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07937_ top.CPU.control_unit.instruction\[28\] net1046 net899 vssd1 vssd1 vccd1 vccd1
+ _03576_ sky130_fd_sc_hd__o21a_1
XANTENNA__11304__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout756_A net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10658__A2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07868_ net625 _03498_ _03506_ vssd1 vssd1 vccd1 vccd1 _03507_ sky130_fd_sc_hd__and3_1
XFILLER_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08720__A1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09607_ net703 _05244_ _05245_ vssd1 vssd1 vccd1 vccd1 _05246_ sky130_fd_sc_hd__or3_1
XFILLER_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16314__RESET_B net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout544_X net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout923_A net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07799_ net621 _03433_ _03434_ _03437_ vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout1286_X net1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09538_ top.CPU.registers.data\[161\] top.CPU.registers.data\[129\] net835 vssd1
+ vssd1 vccd1 vccd1 _05177_ sky130_fd_sc_hd__mux2_1
XFILLER_12_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11025__B net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12280__A1 _05465_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout711_X net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09469_ net695 _05106_ _05107_ vssd1 vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__and3_1
XANTENNA__09681__C1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout809_X net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11500_ _06633_ net258 net255 net3312 vssd1 vssd1 vccd1 vccd1 _02024_ sky130_fd_sc_hd__a22o_1
XANTENNA__13521__A _03984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12480_ _06979_ _06988_ _06978_ vssd1 vssd1 vccd1 vccd1 _06989_ sky130_fd_sc_hd__a21boi_1
XFILLER_12_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10864__B net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11431_ net565 net138 net539 vssd1 vssd1 vccd1 vccd1 _06718_ sky130_fd_sc_hd__and3_1
XFILLER_22_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08236__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09433__C1 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10043__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11362_ net3915 net285 net276 _06465_ vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__a22o_1
X_13101_ top.SPI.count\[1\] top.SPI.count\[0\] vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__nand2_1
XANTENNA__11791__B1 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07995__C1 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10313_ net403 _05943_ vssd1 vssd1 vccd1 vccd1 _05945_ sky130_fd_sc_hd__nand2_1
XFILLER_138_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11293_ net3391 net290 net357 _05808_ vssd1 vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__a22o_1
XFILLER_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13032_ net2768 _07441_ net895 vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__mux2_1
XFILLER_112_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09446__A _05084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11695__B net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10244_ _03167_ _05878_ vssd1 vssd1 vccd1 vccd1 _05879_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_167_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11543__B1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07747__C1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1101 net1103 vssd1 vssd1 vccd1 vccd1 net1101 sky130_fd_sc_hd__clkbuf_4
Xfanout1112 net1113 vssd1 vssd1 vccd1 vccd1 net1112 sky130_fd_sc_hd__clkbuf_4
X_10175_ net3860 net225 net313 _05811_ vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__a22o_1
XFILLER_121_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1123 net1127 vssd1 vssd1 vccd1 vccd1 net1123 sky130_fd_sc_hd__clkbuf_4
Xfanout1134 net1135 vssd1 vssd1 vccd1 vccd1 net1134 sky130_fd_sc_hd__clkbuf_4
XFILLER_120_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1145 net1146 vssd1 vssd1 vccd1 vccd1 net1145 sky130_fd_sc_hd__clkbuf_4
XFILLER_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_128_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1156 net1157 vssd1 vssd1 vccd1 vccd1 net1156 sky130_fd_sc_hd__clkbuf_4
Xfanout1167 net1168 vssd1 vssd1 vccd1 vccd1 net1167 sky130_fd_sc_hd__clkbuf_4
X_14564__734 clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 net2203 sky130_fd_sc_hd__inv_2
X_14983_ clknet_leaf_96_clk _01228_ net1247 vssd1 vssd1 vccd1 vccd1 top.SPI.paroutput\[22\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout180 _06777_ vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__buf_4
XANTENNA__10104__B _05665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1178 net1179 vssd1 vssd1 vccd1 vccd1 net1178 sky130_fd_sc_hd__clkbuf_2
Xfanout191 _06767_ vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__clkbuf_8
Xfanout1189 net1192 vssd1 vssd1 vccd1 vccd1 net1189 sky130_fd_sc_hd__clkbuf_4
XFILLER_47_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11846__A1 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14605__775 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 net2244 sky130_fd_sc_hd__inv_2
XANTENNA__13599__A1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11216__A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15604_ net1938 _01814_ net1119 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[404\]
+ sky130_fd_sc_hd__dfrtp_1
X_12816_ _07267_ _07268_ vssd1 vssd1 vccd1 vccd1 _07269_ sky130_fd_sc_hd__or2_1
X_13796_ net26 net1050 net885 net3952 vssd1 vssd1 vccd1 vccd1 _02677_ sky130_fd_sc_hd__o22a_1
XANTENNA__09267__A2 net1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15535_ net1869 _01745_ net1096 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[335\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11074__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12747_ _07196_ _07198_ _07194_ vssd1 vssd1 vccd1 vccd1 _07206_ sky130_fd_sc_hd__o21ai_1
XFILLER_97_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09672__C1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10282__B1 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12678_ _07142_ _07143_ vssd1 vssd1 vccd1 vccd1 _07144_ sky130_fd_sc_hd__nor2_1
XANTENNA__10821__A2 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15466_ net1800 _01676_ net1089 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[266\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09019__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11629_ _03173_ net498 vssd1 vssd1 vccd1 vccd1 _06756_ sky130_fd_sc_hd__nand2_4
XANTENNA__12023__A1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09424__C1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15397_ net1731 _01607_ net1083 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[197\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08322__S0 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold606 top.CPU.registers.data\[653\] vssd1 vssd1 vccd1 vccd1 net3163 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11782__B1 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold617 top.CPU.registers.data\[371\] vssd1 vssd1 vccd1 vccd1 net3174 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold628 top.CPU.registers.data\[733\] vssd1 vssd1 vccd1 vccd1 net3185 sky130_fd_sc_hd__dlygate4sd3_1
X_13917__87 clknet_leaf_130_clk vssd1 vssd1 vccd1 vccd1 net1556 sky130_fd_sc_hd__inv_2
XFILLER_171_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold639 top.CPU.registers.data\[433\] vssd1 vssd1 vccd1 vccd1 net3196 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07575__S net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16018_ net2352 _02228_ net1103 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[818\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_143_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11534__B1 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08840_ top.CPU.registers.data\[1003\] top.CPU.registers.data\[971\] net964 vssd1
+ vssd1 vccd1 vccd1 _04479_ sky130_fd_sc_hd__mux2_1
XANTENNA__10888__A2 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12988__Y _07418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1306 top.CPU.registers.data_out_r1_prev\[19\] vssd1 vssd1 vccd1 vccd1 net3863
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1317 top.SPI.timem\[18\] vssd1 vssd1 vccd1 vccd1 net3874 sky130_fd_sc_hd__dlygate4sd3_1
X_08771_ net789 _04408_ _04409_ net692 vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__a31o_1
Xhold1328 top.I2C.data_out\[5\] vssd1 vssd1 vccd1 vccd1 net3885 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1339 top.SPI.timem\[16\] vssd1 vssd1 vccd1 vccd1 net3896 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13826__A2 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07722_ net621 _03356_ _03357_ _03360_ vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__a31oi_2
XFILLER_66_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11837__A1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_7_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08163__C1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10949__B _03170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08702__A1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07604__A net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09091__A _04698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07653_ _03245_ _03262_ _03264_ vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__or3_4
XFILLER_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07910__C1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11126__A net1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07584_ net756 _03218_ _03219_ _03222_ net711 vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__o311a_1
XANTENNA__09258__A2 net1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09323_ top.CPU.registers.data\[164\] net1392 net829 top.CPU.registers.data\[132\]
+ net708 vssd1 vssd1 vccd1 vccd1 _04962_ sky130_fd_sc_hd__a221o_1
XFILLER_22_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12262__A1 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11065__A2 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10965__A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09663__C1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout337_A net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09254_ top.CPU.registers.data\[805\] top.CPU.registers.data\[773\] net966 vssd1
+ vssd1 vccd1 vccd1 _04893_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1079_A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08435__A net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10684__B _06139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08205_ net677 _03839_ _03840_ _03843_ net612 vssd1 vssd1 vccd1 vccd1 _03844_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_32_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12014__A1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10585__A2_N net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09185_ net742 _04817_ _04816_ net768 vssd1 vssd1 vccd1 vccd1 _04824_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout504_A net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout125_X net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08136_ net627 _03771_ _03772_ net612 vssd1 vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__a31o_1
XFILLER_174_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08722__X _04361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11773__B1 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08067_ net674 _03701_ _03702_ _03705_ net610 vssd1 vssd1 vccd1 vccd1 _03706_ sky130_fd_sc_hd__a311oi_1
XFILLER_162_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07992__A2 net1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08170__A net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14251__421 clknet_leaf_149_clk vssd1 vssd1 vccd1 vccd1 net1890 sky130_fd_sc_hd__inv_2
XFILLER_68_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout494_X net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11525__B1 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout873_A net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14548__718 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 net2187 sky130_fd_sc_hd__inv_2
XANTENNA__07744__A2 net1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11540__A3 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout661_X net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08969_ top.CPU.registers.data\[745\] net1386 net805 top.CPU.registers.data\[713\]
+ net761 vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout759_X net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_162_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11980_ _06537_ net351 net182 net3609 vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__a22o_1
XFILLER_84_47 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08154__C1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10859__B _03180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10931_ net483 net459 _06512_ net221 net3328 vssd1 vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__a32o_1
XFILLER_17_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout926_X net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13650_ net3191 _07315_ net663 vssd1 vssd1 vccd1 vccd1 _02584_ sky130_fd_sc_hd__mux2_1
X_10862_ net323 net435 vssd1 vssd1 vccd1 vccd1 _06469_ sky130_fd_sc_hd__nand2_4
XFILLER_71_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12601_ _03139_ top.SPI.count\[3\] _07100_ vssd1 vssd1 vccd1 vccd1 _07102_ sky130_fd_sc_hd__a21o_1
X_13581_ net3970 net579 _03014_ _03015_ vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__a22o_1
XFILLER_140_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11056__A2 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08457__B1 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12253__A1 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12419__X _06945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10793_ _05124_ _05270_ _06402_ net371 vssd1 vssd1 vccd1 vccd1 _06404_ sky130_fd_sc_hd__a31o_1
XANTENNA__08616__Y _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12532_ net547 _03323_ _07040_ vssd1 vssd1 vccd1 vccd1 _07041_ sky130_fd_sc_hd__and3_1
X_15320_ net1654 _01530_ net1103 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[120\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10803__A2 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12463_ _06970_ _06971_ _06969_ vssd1 vssd1 vccd1 vccd1 _06972_ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_193_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15251_ net1585 _01461_ net1176 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[51\]
+ sky130_fd_sc_hd__dfrtp_1
X_11414_ _06548_ net276 net267 net3411 vssd1 vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__a22o_1
X_15182_ net1519 _01392_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r1_prev\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_166_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12394_ net599 vssd1 vssd1 vccd1 vccd1 _06932_ sky130_fd_sc_hd__inv_2
XFILLER_137_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_169_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_73_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09421__A2 net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11764__B1 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13397__S net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11345_ net3704 net287 net281 _06127_ vssd1 vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__a22o_1
XFILLER_152_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13505__A1 top.CPU.data_out\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07983__A2 net1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13505__B2 _02972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10319__A1 _03650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08080__A _03683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11276_ net3015 net295 _06695_ net318 vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__a22o_1
XFILLER_141_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11516__B1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13015_ top.SPI.parameters\[9\] top.SPI.paroutput\[1\] net1357 vssd1 vssd1 vccd1
+ vccd1 _07433_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_18_Left_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09185__A1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10227_ _05667_ _05861_ vssd1 vssd1 vccd1 vccd1 _05862_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_88_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10115__A net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10158_ _05647_ _05658_ net308 vssd1 vssd1 vccd1 vccd1 _05795_ sky130_fd_sc_hd__mux2_1
XFILLER_121_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_131_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold3 top.I2C.I2C_state\[0\] vssd1 vssd1 vccd1 vccd1 net2560 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_12_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11819__A1 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10089_ _03889_ net379 vssd1 vssd1 vccd1 vccd1 _05727_ sky130_fd_sc_hd__or2_1
X_14966_ clknet_leaf_97_clk net3222 net1253 vssd1 vssd1 vccd1 vccd1 top.SPI.paroutput\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_11_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11295__A2 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08696__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_146_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11047__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_26_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13779_ net7 net1051 net886 top.mmio.mem_data_i\[14\] vssd1 vssd1 vccd1 vccd1 _02660_
+ sky130_fd_sc_hd__a22o_1
XFILLER_95_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15518_ net1852 _01728_ net1237 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[318\]
+ sky130_fd_sc_hd__dfrtp_1
X_16498_ clknet_leaf_41_clk _02660_ net1116 vssd1 vssd1 vccd1 vccd1 top.mmio.mem_data_i\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_14692__862 clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 net2331 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_44_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_4_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_4_0_clk sky130_fd_sc_hd__clkbuf_8
X_15449_ net1783 _01659_ net1245 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[249\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_159_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11112__C _06010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11755__B1 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold403 top.CPU.registers.data\[431\] vssd1 vssd1 vccd1 vccd1 net2960 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07959__C1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold414 net77 vssd1 vssd1 vccd1 vccd1 net2971 sky130_fd_sc_hd__dlygate4sd3_1
Xhold425 top.CPU.addressnew\[23\] vssd1 vssd1 vccd1 vccd1 net2982 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14235__405 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 net1874 sky130_fd_sc_hd__inv_2
Xhold436 top.CPU.registers.data\[886\] vssd1 vssd1 vccd1 vccd1 net2993 sky130_fd_sc_hd__dlygate4sd3_1
Xhold447 top.CPU.registers.data\[772\] vssd1 vssd1 vccd1 vccd1 net3004 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10951__C net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07974__A2 _03610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold458 top.CPU.registers.data\[804\] vssd1 vssd1 vccd1 vccd1 net3015 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09941_ _05577_ _05578_ _05579_ vssd1 vssd1 vccd1 vccd1 _05580_ sky130_fd_sc_hd__or3_2
Xhold469 top.CPU.registers.data\[864\] vssd1 vssd1 vccd1 vccd1 net3026 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11770__A3 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11507__B1 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout905 net906 vssd1 vssd1 vccd1 vccd1 net905 sky130_fd_sc_hd__clkbuf_4
Xfanout916 net925 vssd1 vssd1 vccd1 vccd1 net916 sky130_fd_sc_hd__clkbuf_2
Xfanout927 net949 vssd1 vssd1 vccd1 vccd1 net927 sky130_fd_sc_hd__buf_2
X_09872_ _03511_ _03579_ _05510_ vssd1 vssd1 vccd1 vccd1 _05511_ sky130_fd_sc_hd__o21a_1
Xfanout938 net949 vssd1 vssd1 vccd1 vccd1 net938 sky130_fd_sc_hd__clkbuf_4
Xfanout949 _03352_ vssd1 vssd1 vccd1 vccd1 net949 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12180__B1 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08823_ net1400 _03160_ _03985_ vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__o21a_1
Xhold1103 top.SPI.paroutput\[31\] vssd1 vssd1 vccd1 vccd1 net3660 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1114 top.CPU.registers.data\[115\] vssd1 vssd1 vccd1 vccd1 net3671 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout287_A net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1125 top.CPU.registers.data\[952\] vssd1 vssd1 vccd1 vccd1 net3682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1136 top.CPU.registers.data\[994\] vssd1 vssd1 vccd1 vccd1 net3693 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08754_ _04391_ _04392_ net453 vssd1 vssd1 vccd1 vccd1 _04393_ sky130_fd_sc_hd__mux2_1
Xhold1147 top.CPU.registers.data\[753\] vssd1 vssd1 vccd1 vccd1 net3704 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1158 top.I2C.bit_timer_counter\[7\] vssd1 vssd1 vccd1 vccd1 net3715 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1169 top.CPU.addressnew\[24\] vssd1 vssd1 vccd1 vccd1 net3726 sky130_fd_sc_hd__dlygate4sd3_1
X_07705_ top.CPU.registers.data\[831\] net999 vssd1 vssd1 vccd1 vccd1 _03344_ sky130_fd_sc_hd__or2_1
XANTENNA__08687__A0 _04324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08685_ net689 _04323_ _04296_ vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_68_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10031__Y _05670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_92_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_92_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout454_A net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1196_A net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07636_ net1279 _03158_ _03272_ _03263_ _03152_ vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__a32oi_1
XFILLER_54_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12894__B _05362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11038__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07567_ net1047 _03163_ net1038 net1308 vssd1 vssd1 vccd1 vccd1 _03206_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout621_A net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout242_X net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1363_A top.CPU.alu.immediate\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11290__S net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10246__B1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09306_ top.CPU.registers.data\[388\] net1299 net1020 top.CPU.registers.data\[420\]
+ net918 vssd1 vssd1 vccd1 vccd1 _04945_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout719_A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07498_ net2617 vssd1 vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__inv_2
XFILLER_167_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11994__B1 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09237_ top.CPU.registers.data\[965\] net1310 net841 top.CPU.registers.data\[997\]
+ net713 vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout507_X net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09168_ top.CPU.registers.data\[70\] net1317 net847 top.CPU.registers.data\[102\]
+ net767 vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout990_A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11746__B1 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08119_ top.CPU.registers.data\[693\] top.CPU.registers.data\[661\] net993 vssd1
+ vssd1 vccd1 vccd1 _03758_ sky130_fd_sc_hd__mux2_1
XFILLER_134_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09099_ top.CPU.registers.data\[167\] top.CPU.registers.data\[135\] net832 vssd1
+ vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__mux2_1
XFILLER_162_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11130_ net572 net524 _06213_ vssd1 vssd1 vccd1 vccd1 _06623_ sky130_fd_sc_hd__and3_1
XFILLER_150_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13499__B1 _02968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold970 top.CPU.registers.data\[777\] vssd1 vssd1 vccd1 vccd1 net3527 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold981 top.CPU.registers.data\[354\] vssd1 vssd1 vccd1 vccd1 net3538 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout876_X net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11061_ net3613 net366 _06587_ net323 vssd1 vssd1 vccd1 vccd1 _02321_ sky130_fd_sc_hd__a22o_1
Xhold992 top.CPU.registers.data\[57\] vssd1 vssd1 vccd1 vccd1 net3549 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08375__C1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10012_ _03476_ _03544_ net379 vssd1 vssd1 vccd1 vccd1 _05651_ sky130_fd_sc_hd__mux2_1
X_14019__189 clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 net1658 sky130_fd_sc_hd__inv_2
XANTENNA__07943__S net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11513__A3 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07515__Y _03154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input15_A DAT_I[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11963_ _06512_ net344 net230 net3382 vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__a22o_1
XANTENNA__13671__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_83_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_clk sky130_fd_sc_hd__clkbuf_8
X_13702_ top.SPI.timem\[4\] _03054_ vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__and2_1
X_10914_ net479 net456 _06502_ net220 net3059 vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__a32o_1
X_11894_ net149 net3522 net190 vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__mux2_1
XFILLER_32_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16421_ clknet_leaf_56_clk _00003_ net1141 vssd1 vssd1 vccd1 vccd1 top.I2C.I2C_state\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10845_ net549 net370 net444 _05267_ vssd1 vssd1 vccd1 vccd1 _06453_ sky130_fd_sc_hd__a31o_1
X_13633_ net3855 _07154_ net664 vssd1 vssd1 vccd1 vccd1 _02567_ sky130_fd_sc_hd__mux2_1
XFILLER_32_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14676__846 clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 net2315 sky130_fd_sc_hd__inv_2
X_16352_ clknet_leaf_68_clk _02561_ net1167 vssd1 vssd1 vccd1 vccd1 top.CPU.addressnew\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_13564_ top.CPU.alu.program_counter\[6\] _06352_ net1348 vssd1 vssd1 vccd1 vccd1
+ _03005_ sky130_fd_sc_hd__mux2_1
X_10776_ net511 _05555_ _06387_ _06383_ _06377_ vssd1 vssd1 vccd1 vccd1 _06388_ sky130_fd_sc_hd__a311o_1
XFILLER_158_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11985__B1 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15303_ net1637 _01513_ net1192 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[103\]
+ sky130_fd_sc_hd__dfrtp_1
X_12515_ _07018_ _07023_ vssd1 vssd1 vccd1 vccd1 _07024_ sky130_fd_sc_hd__nor2_1
X_14420__590 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 net2059 sky130_fd_sc_hd__inv_2
X_16283_ clknet_leaf_62_clk _02493_ net1161 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.toreg\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13495_ net1400 net874 _03248_ _02965_ vssd1 vssd1 vccd1 vccd1 _02966_ sky130_fd_sc_hd__a31oi_4
XANTENNA__08850__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14717__887 clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 net2356 sky130_fd_sc_hd__inv_2
XFILLER_145_418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12446_ net898 _06959_ vssd1 vssd1 vccd1 vccd1 _00049_ sky130_fd_sc_hd__nor2_1
X_15234_ net1568 _01444_ net1175 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11737__B1 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12377_ top.I2C.byte_manager_state\[0\] top.I2C.byte_manager_done vssd1 vssd1 vccd1
+ vccd1 _06916_ sky130_fd_sc_hd__nor2_1
XFILLER_153_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15165_ net1502 _01375_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r1_prev\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_154_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_26_Left_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11328_ net3082 net289 net357 net130 vssd1 vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__a22o_1
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15096_ net1478 _01309_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r2_prev\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10116__Y _05754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11259_ net471 _06685_ vssd1 vssd1 vccd1 vccd1 _06686_ sky130_fd_sc_hd__nor2_1
XFILLER_68_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10712__A1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08381__A2 _04019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15998_ net2332 _02208_ net1237 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[798\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09005__S1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_167_Right_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14949_ clknet_leaf_52_clk _01195_ net1133 vssd1 vssd1 vccd1 vccd1 top.I2C.bit_timer_counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11268__A2 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08669__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_74_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_35_Left_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08133__A2 net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08470_ net943 _04108_ vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__or2_1
XFILLER_35_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16619_ net1347 vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12217__A1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10779__A1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11976__B1 net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11440__A2 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09022_ net452 _04660_ vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__nand2_1
XFILLER_108_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10962__B net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09397__A1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold200 top.SPI.parameters\[29\] vssd1 vssd1 vccd1 vccd1 net2757 sky130_fd_sc_hd__dlygate4sd3_1
Xhold211 top.SPI.paroutput\[17\] vssd1 vssd1 vccd1 vccd1 net2768 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09087__Y _04726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10307__X _05939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout202_A _06753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold222 top.CPU.registers.data\[291\] vssd1 vssd1 vccd1 vccd1 net2779 sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 top.SPI.counter\[1\] vssd1 vssd1 vccd1 vccd1 net2790 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 top.SPI.paroutput\[13\] vssd1 vssd1 vccd1 vccd1 net2801 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14934__RESET_B net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11743__A3 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold255 top.CPU.registers.data\[190\] vssd1 vssd1 vccd1 vccd1 net2812 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold266 top.CPU.addressnew\[28\] vssd1 vssd1 vccd1 vccd1 net2823 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10026__Y _05665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold277 top.CPU.registers.data\[136\] vssd1 vssd1 vccd1 vccd1 net2834 sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 top.CPU.registers.data\[629\] vssd1 vssd1 vccd1 vccd1 net2845 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09924_ _04765_ _04795_ vssd1 vssd1 vccd1 vccd1 _05563_ sky130_fd_sc_hd__and2_1
Xfanout702 net703 vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__buf_4
Xhold299 top.CPU.registers.data\[839\] vssd1 vssd1 vccd1 vccd1 net2856 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout713 net736 vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__clkbuf_4
XFILLER_172_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout724 net735 vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1111_A net1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1209_A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout735 net736 vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__clkbuf_4
Xfanout746 net747 vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__buf_2
XFILLER_113_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input7_A DAT_I[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout757 net759 vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__clkbuf_4
X_09855_ top.CPU.registers.data\[474\] net1305 net1027 top.CPU.registers.data\[506\]
+ net922 vssd1 vssd1 vccd1 vccd1 _05494_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_142_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout192_X net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout768 net771 vssd1 vssd1 vccd1 vccd1 net768 sky130_fd_sc_hd__clkbuf_4
XFILLER_100_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout779 net780 vssd1 vssd1 vccd1 vccd1 net779 sky130_fd_sc_hd__clkbuf_4
X_13901__71 clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 net1540 sky130_fd_sc_hd__inv_2
XANTENNA_fanout669_A _00000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08372__A2 net1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08806_ net617 _04437_ _04443_ _04444_ vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__o22a_1
X_09786_ net939 _05400_ _05401_ net956 vssd1 vssd1 vccd1 vccd1 _05425_ sky130_fd_sc_hd__o211a_1
XFILLER_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08109__C1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07580__B1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_134_Right_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12456__A1 _03405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08737_ _04374_ _04375_ net673 vssd1 vssd1 vccd1 vccd1 _04376_ sky130_fd_sc_hd__o21ai_1
XFILLER_38_170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_65_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout457_X net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout836_A net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14363__533 clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 net2002 sky130_fd_sc_hd__inv_2
XANTENNA__08124__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08594__S net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08668_ _04305_ _04306_ net675 vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_83_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_1007 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07619_ top.CPU.control_unit.instruction\[26\] top.CPU.control_unit.instruction\[25\]
+ _03257_ vssd1 vssd1 vccd1 vccd1 _03258_ sky130_fd_sc_hd__nor3_2
XFILLER_42_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09609__C1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08599_ _04236_ _04237_ net673 vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout624_X net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08607__B net1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1366_X net1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10630_ net548 _05283_ _06248_ vssd1 vssd1 vccd1 vccd1 _06249_ sky130_fd_sc_hd__o21ai_1
X_14404__574 clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 net2043 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_157_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11967__B1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10561_ _04330_ _05569_ _06156_ vssd1 vssd1 vccd1 vccd1 _06183_ sky130_fd_sc_hd__o21a_1
XFILLER_128_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11033__B net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12300_ net2622 _04697_ net1098 vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__mux2_1
XANTENNA__07938__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13280_ top.CPU.handler.state\[5\] _02825_ vssd1 vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_118_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10492_ _03315_ _05293_ _05918_ _05981_ _06116_ vssd1 vssd1 vccd1 vccd1 _06117_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout993_X net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10872__B _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11719__B1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12231_ net566 net363 _06696_ net170 top.CPU.registers.data\[35\] vssd1 vssd1 vccd1
+ vccd1 _06882_ sky130_fd_sc_hd__a32o_1
XFILLER_136_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11195__B2 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12162_ top.CPU.registers.data\[71\] net652 vssd1 vssd1 vccd1 vccd1 _06849_ sky130_fd_sc_hd__or2_1
XANTENNA__08060__A1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_420 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11113_ net490 net467 _06614_ net303 net2993 vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__a32o_1
XFILLER_123_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12093_ _06628_ net244 net176 top.CPU.registers.data\[106\] vssd1 vssd1 vccd1 vccd1
+ _06815_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_4_15_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07526__X _03165_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15921_ net2255 _02131_ net1178 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[721\]
+ sky130_fd_sc_hd__dfrtp_1
X_11044_ _05934_ net539 vssd1 vssd1 vccd1 vccd1 _06581_ sky130_fd_sc_hd__and2_1
XANTENNA__08899__B1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11498__A2 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13971__141 clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 net1610 sky130_fd_sc_hd__inv_2
X_15852_ net2186 _02062_ net1078 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[652\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_92_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10170__A2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07571__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11208__B net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15783_ net2117 _01993_ net1197 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[583\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_56_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_clk sky130_fd_sc_hd__clkbuf_8
X_12995_ top.SPI.register\[2\] net1354 top.SPI.register\[0\] _07117_ _07423_ vssd1
+ vssd1 vccd1 vccd1 _07424_ sky130_fd_sc_hd__o311a_1
XANTENNA__09848__C1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10458__B1 _03167_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11946_ _06035_ net3679 net231 vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10539__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11877_ _06056_ net3311 net189 vssd1 vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__mux2_1
X_16404_ clknet_leaf_64_clk _00075_ net1145 vssd1 vssd1 vccd1 vccd1 top.wm.curr_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11224__A net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13616_ net2637 _03036_ net581 vssd1 vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__mux2_1
XFILLER_60_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10828_ _05195_ _05547_ vssd1 vssd1 vccd1 vccd1 _06437_ sky130_fd_sc_hd__or2_1
XANTENNA__09615__A2 net1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11958__B1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16335_ clknet_leaf_66_clk _02544_ net1166 vssd1 vssd1 vccd1 vccd1 top.CPU.addressnew\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13547_ _07056_ _02993_ vssd1 vssd1 vccd1 vccd1 _02994_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_41_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11422__A2 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10759_ net600 _06371_ vssd1 vssd1 vccd1 vccd1 _06372_ sky130_fd_sc_hd__nor2_1
XFILLER_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16266_ clknet_leaf_44_clk _02476_ net1124 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.toreg\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13478_ net3978 _02960_ net124 vssd1 vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__mux2_1
XANTENNA__09379__B2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15217_ net1551 _01427_ net1189 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_12429_ net1340 top.I2C.output_state\[13\] net3117 vssd1 vssd1 vccd1 vccd1 _06951_
+ sky130_fd_sc_hd__a21oi_1
X_16197_ net2531 _02407_ net1083 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[997\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07929__A2 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15148_ clknet_leaf_48_clk _01358_ net1130 vssd1 vssd1 vccd1 vccd1 top.I2C.data_out\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_126_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10933__A1 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07970_ top.CPU.registers.data_out_r1_prev\[24\] net874 net636 _03595_ vssd1 vssd1
+ vccd1 vccd1 _03609_ sky130_fd_sc_hd__o22a_1
X_15079_ clknet_leaf_51_clk _00057_ net1132 vssd1 vssd1 vccd1 vccd1 top.I2C.output_state\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_142_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08339__C1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11489__A2 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12502__B _04855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14050__220 clknet_leaf_140_clk vssd1 vssd1 vccd1 vccd1 net1689 sky130_fd_sc_hd__inv_2
XANTENNA__08354__A2 net1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09640_ _04664_ _04666_ vssd1 vssd1 vccd1 vccd1 _05279_ sky130_fd_sc_hd__nand2_2
XFILLER_68_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14347__517 clknet_leaf_135_clk vssd1 vssd1 vccd1 vccd1 net1986 sky130_fd_sc_hd__inv_2
X_09571_ top.CPU.registers.data\[96\] net1005 net951 _05196_ vssd1 vssd1 vccd1 vccd1
+ _05210_ sky130_fd_sc_hd__a211o_1
XANTENNA__11118__B net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_47_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09303__A1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10449__B1 _05670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08522_ top.CPU.registers.data\[400\] net1291 net1011 top.CPU.registers.data\[432\]
+ net909 vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__a221o_1
XANTENNA__09854__A2 net1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08453_ _03117_ net1033 vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__or2_1
XANTENNA__11661__A2 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout152_A net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11134__A net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08384_ top.CPU.registers.data\[306\] top.CPU.registers.data\[274\] net982 vssd1
+ vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__mux2_1
XFILLER_51_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11949__B1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11413__A2 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10973__A net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout417_A _03242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1061_A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1159_A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09005_ _04640_ _04641_ _04642_ _04643_ net672 net900 vssd1 vssd1 vccd1 vccd1 _04644_
+ sky130_fd_sc_hd__mux4_1
XFILLER_117_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout205_X net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11177__A1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1326_A net1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09826__X _05465_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10924__A1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout786_A net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09790__A1 top.CPU.control_unit.instruction\[27\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_160_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13955__125 clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 net1594 sky130_fd_sc_hd__inv_2
Xfanout510 _05669_ vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__clkbuf_4
X_13878__48 clknet_leaf_175_clk vssd1 vssd1 vccd1 vccd1 net1517 sky130_fd_sc_hd__inv_2
XANTENNA__12126__B1 _06749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09274__A net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout521 net522 vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__buf_2
XFILLER_104_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09907_ net372 _05266_ vssd1 vssd1 vccd1 vccd1 _05546_ sky130_fd_sc_hd__nor2_1
Xfanout532 net533 vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__buf_4
XFILLER_76_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13508__B _02966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout543 net544 vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__buf_2
Xfanout554 _02847_ vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout953_A net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout565 net569 vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__buf_4
XANTENNA_fanout574_X net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09542__A1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout576 _03169_ vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__buf_4
Xfanout587 net589 vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__clkbuf_4
X_09838_ top.CPU.registers.data\[602\] net1305 net1027 top.CPU.registers.data\[634\]
+ net946 vssd1 vssd1 vccd1 vccd1 _05477_ sky130_fd_sc_hd__a221o_1
Xfanout598 _07088_ vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10213__A net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12839__S net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09769_ top.CPU.registers.data\[59\] top.CPU.registers.data\[27\] net991 vssd1 vssd1
+ vccd1 vccd1 _05408_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout741_X net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_38_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout839_X net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11800_ _06646_ net235 _06764_ vssd1 vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_159_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _07218_ _07235_ _07223_ vssd1 vssd1 vccd1 vccd1 _07236_ sky130_fd_sc_hd__a21o_1
XFILLER_61_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09845__A2 net1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11101__B2 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08502__C1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11731_ _06578_ net499 net193 net3762 vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_25_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11652__A2 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ net435 net196 vssd1 vssd1 vccd1 vccd1 _06757_ sky130_fd_sc_hd__nand2_8
XFILLER_42_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13401_ top.CPU.control_unit.instruction\[25\] _02918_ net671 vssd1 vssd1 vccd1 vccd1
+ _02459_ sky130_fd_sc_hd__mux2_1
X_10613_ net573 net515 net439 _06231_ vssd1 vssd1 vccd1 vccd1 _06233_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_172_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08805__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11593_ _03184_ _06751_ vssd1 vssd1 vccd1 vccd1 _06752_ sky130_fd_sc_hd__or2_4
XANTENNA__10883__A net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11404__A2 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16120_ net2454 _02330_ net1150 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[920\]
+ sky130_fd_sc_hd__dfrtp_1
X_10544_ _05668_ _05673_ vssd1 vssd1 vccd1 vccd1 _06167_ sky130_fd_sc_hd__or2_1
X_13332_ top.mmio.mem_data_i\[7\] net592 net1343 vssd1 vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__a21o_1
XANTENNA__09449__A _05087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08353__A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16051_ net2385 _02261_ net1177 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[851\]
+ sky130_fd_sc_hd__dfrtp_1
X_14491__661 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 net2130 sky130_fd_sc_hd__inv_2
X_10475_ _05297_ _05584_ _06061_ vssd1 vssd1 vccd1 vccd1 _06101_ sky130_fd_sc_hd__or3_1
X_13263_ net3885 _02814_ _02816_ net1053 vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__a22o_1
XFILLER_157_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14788__958 clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 net2427 sky130_fd_sc_hd__inv_2
X_15002_ clknet_leaf_97_clk net3667 net1253 vssd1 vssd1 vccd1 vccd1 top.SPI.parameters\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08569__C1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12214_ top.CPU.registers.data\[44\] net646 vssd1 vssd1 vccd1 vccd1 _06874_ sky130_fd_sc_hd__or2_1
XANTENNA__08033__A1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13194_ top.I2C.within_byte_counter_reading\[0\] top.I2C.within_byte_counter_reading\[1\]
+ top.I2C.within_byte_counter_reading\[2\] vssd1 vssd1 vccd1 vccd1 _02774_ sky130_fd_sc_hd__and3b_2
XANTENNA__09230__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10107__B net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09781__A1 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12145_ net146 net356 net236 _06840_ vssd1 vssd1 vccd1 vccd1 _01490_ sky130_fd_sc_hd__a31o_1
XFILLER_151_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14034__204 clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 net1673 sky130_fd_sc_hd__inv_2
XFILLER_123_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07792__B1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14829__999 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 net2468 sky130_fd_sc_hd__inv_2
X_12076_ _06617_ net244 _06806_ net178 net3671 vssd1 vssd1 vccd1 vccd1 _01525_ sky130_fd_sc_hd__a32o_1
XANTENNA__07659__C_N _03292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15904_ net2238 _02114_ net1090 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[704\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11027_ net3725 net219 _06571_ net319 vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__a22o_1
XANTENNA__09533__A1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10123__A net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08741__C1 net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13617__A0 top.CPU.alu.program_counter\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15835_ net2169 _02045_ net1209 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[635\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_29_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_8
X_13892__62 clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 net1531 sky130_fd_sc_hd__inv_2
XANTENNA__09297__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15766_ net2100 _01976_ net1231 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[566\]
+ sky130_fd_sc_hd__dfrtp_1
X_12978_ _07411_ top.I2C.bit_timer_state\[0\] _07410_ vssd1 vssd1 vccd1 vccd1 _01199_
+ sky130_fd_sc_hd__and3b_1
XFILLER_45_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11929_ net3319 net185 net348 _06413_ vssd1 vssd1 vccd1 vccd1 _01637_ sky130_fd_sc_hd__a22o_1
XANTENNA__11643__A2 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15697_ net2031 _01907_ net1175 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[497\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14732__902 clknet_leaf_189_clk vssd1 vssd1 vccd1 vccd1 net2371 sky130_fd_sc_hd__inv_2
X_16318_ clknet_leaf_95_clk _02527_ net1246 vssd1 vssd1 vccd1 vccd1 top.CPU.data_out\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08272__A1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16253__Q top.CPU.control_unit.instruction\[29\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16249_ clknet_leaf_60_clk _02459_ net1139 vssd1 vssd1 vccd1 vccd1 top.CPU.control_unit.instruction\[25\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_11_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09078__B net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput102 net102 vssd1 vssd1 vccd1 vccd1 SEL_O[2] sky130_fd_sc_hd__buf_2
Xoutput113 net113 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_58_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13939__109 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 net1578 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_58_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08024__A1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08550__X _04189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12108__B1 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10382__A2 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07783__B1 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09094__A top.CPU.alu.program_counter\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08202__S net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07953_ net793 _03586_ _03587_ net744 vssd1 vssd1 vccd1 vccd1 _03592_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_71_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07884_ top.CPU.registers.data\[988\] net1332 net863 top.CPU.registers.data\[1020\]
+ net729 vssd1 vssd1 vccd1 vccd1 _03523_ sky130_fd_sc_hd__a221o_1
XFILLER_110_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09623_ net741 _05255_ _05256_ net765 vssd1 vssd1 vccd1 vccd1 _05262_ sky130_fd_sc_hd__o211a_1
XANTENNA__13608__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout367_A net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09554_ net381 _05192_ vssd1 vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__nand2_1
XANTENNA__09288__B1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11095__B1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08505_ top.CPU.registers.data\[976\] net1322 net853 top.CPU.registers.data\[1008\]
+ net721 vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__a221o_1
XANTENNA__07838__A1 top.CPU.control_unit.instruction\[29\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_52_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09485_ net394 _05123_ vssd1 vssd1 vccd1 vccd1 _05124_ sky130_fd_sc_hd__nand2_2
XANTENNA__11634__A2 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout534_A net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout155_X net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1276_A net1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08436_ _04071_ _04074_ net637 vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__a21o_1
XFILLER_24_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08872__S net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08367_ net792 _04005_ vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout322_X net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14475__645 clknet_leaf_163_clk vssd1 vssd1 vccd1 vccd1 net2114 sky130_fd_sc_hd__inv_2
XANTENNA__08263__A1 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08298_ net796 _03926_ _03927_ net725 vssd1 vssd1 vccd1 vccd1 _03937_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_115_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11311__B net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1329_X net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10260_ _05731_ _05747_ net390 vssd1 vssd1 vccd1 vccd1 _05894_ sky130_fd_sc_hd__mux2_1
XFILLER_11_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14516__686 clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 net2155 sky130_fd_sc_hd__inv_2
XANTENNA__09212__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout691_X net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout789_X net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13519__A _04048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08566__A2 net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10191_ net390 _05826_ vssd1 vssd1 vccd1 vccd1 _05827_ sky130_fd_sc_hd__nand2_1
XANTENNA__07774__B1 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1305 net1306 vssd1 vssd1 vccd1 vccd1 net1305 sky130_fd_sc_hd__buf_2
XFILLER_121_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1316 net1317 vssd1 vssd1 vccd1 vccd1 net1316 sky130_fd_sc_hd__clkbuf_4
Xfanout1327 _03109_ vssd1 vssd1 vccd1 vccd1 net1327 sky130_fd_sc_hd__buf_2
Xfanout340 _02978_ vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout956_X net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1338 _03109_ vssd1 vssd1 vccd1 vccd1 net1338 sky130_fd_sc_hd__clkbuf_4
Xfanout1349 top.CPU.handler.state\[3\] vssd1 vssd1 vccd1 vccd1 net1349 sky130_fd_sc_hd__buf_2
Xfanout351 net352 vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__clkbuf_4
XFILLER_120_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout362 net364 vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11039__A _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout373 net376 vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__clkbuf_4
Xfanout384 net385 vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__buf_2
XFILLER_101_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout395 net398 vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__buf_2
XANTENNA__11322__B2 _06373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12901_ top.CPU.alu.program_counter\[26\] _07337_ vssd1 vssd1 vccd1 vccd1 _07345_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__11873__A2 net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10878__A _05693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15620_ net1954 _01830_ net1221 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[420\]
+ sky130_fd_sc_hd__dfrtp_1
X_12832_ top.CPU.alu.program_counter\[18\] _07283_ net1359 vssd1 vssd1 vccd1 vccd1
+ _01181_ sky130_fd_sc_hd__mux2_1
XFILLER_27_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15551_ net1885 _01761_ net1222 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[351\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07829__A1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ top.CPU.alu.program_counter\[12\] _07208_ vssd1 vssd1 vccd1 vccd1 _07221_
+ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_174_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _06551_ net197 net420 net2885 vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__a22o_1
X_15482_ net1816 _01692_ net1250 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[282\]
+ sky130_fd_sc_hd__dfrtp_1
X_12694_ _07156_ _07157_ vssd1 vssd1 vccd1 vccd1 _07158_ sky130_fd_sc_hd__nand2_1
XANTENNA__13378__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11645_ _06151_ net200 net425 net3139 vssd1 vssd1 vccd1 vccd1 _01906_ sky130_fd_sc_hd__a22o_1
XANTENNA__11389__A1 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput15 DAT_I[21] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
XFILLER_167_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput26 DAT_I[31] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
X_11576_ _06687_ net259 net246 net2798 vssd1 vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__a22o_1
XANTENNA__12050__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput37 gpio_in[2] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_1
X_16103_ net2437 _02313_ net1203 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[903\]
+ sky130_fd_sc_hd__dfrtp_1
X_13315_ net4018 _02855_ net669 vssd1 vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__mux2_1
XFILLER_171_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10527_ net527 _06150_ vssd1 vssd1 vccd1 vccd1 _06151_ sky130_fd_sc_hd__nor2_1
X_16034_ net2368 _02244_ net1174 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[834\]
+ sky130_fd_sc_hd__dfrtp_1
X_13246_ net3900 _02805_ _02807_ _02803_ vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__a22o_1
XFILLER_6_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09203__B1 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10458_ _06082_ _06083_ _03167_ vssd1 vssd1 vccd1 vccd1 _06085_ sky130_fd_sc_hd__a21oi_4
XANTENNA__12889__A1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08557__A2 net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13177_ _03124_ _06911_ vssd1 vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__nand2_1
X_10389_ net548 _03789_ _06017_ vssd1 vssd1 vccd1 vccd1 _06018_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_36_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13148__B _05232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12128_ top.CPU.registers.data\[88\] net650 _03187_ _05962_ net355 vssd1 vssd1 vccd1
+ vccd1 _06832_ sky130_fd_sc_hd__o2111a_1
XFILLER_123_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08309__A2 net1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12059_ top.CPU.registers.data\[123\] net178 vssd1 vssd1 vccd1 vccd1 _06798_ sky130_fd_sc_hd__and2_1
XFILLER_42_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08714__C1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11313__B2 _06212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07714__X _03353_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10788__A _05672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08190__B1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15818_ net2152 _02028_ net1085 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[618\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_92_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09809__A2 net1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16248__Q top.CPU.control_unit.instruction\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15749_ net2083 _01959_ net1062 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[549\]
+ sky130_fd_sc_hd__dfrtp_1
X_09270_ net950 _04908_ _04907_ net611 vssd1 vssd1 vccd1 vccd1 _04909_ sky130_fd_sc_hd__a211o_1
X_14162__332 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 net1801 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14459__629 clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 net2098 sky130_fd_sc_hd__inv_2
X_08221_ top.CPU.alu.program_counter\[22\] net1035 vssd1 vssd1 vccd1 vccd1 _03860_
+ sky130_fd_sc_hd__nor2_1
XFILLER_159_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08152_ top.CPU.registers.data\[343\] net1325 net856 top.CPU.registers.data\[375\]
+ net773 vssd1 vssd1 vccd1 vccd1 _03791_ sky130_fd_sc_hd__a221o_1
XFILLER_158_170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08245__A1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09442__B1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12041__A2 _06779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14203__373 clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 net1842 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_95_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_3_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08083_ _03720_ _03721_ vssd1 vssd1 vccd1 vccd1 _03722_ sky130_fd_sc_hd__nor2_1
XANTENNA__10028__A net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12942__S net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_9_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_174_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09536__B net1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1024_A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07756__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08953__C1 _03342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11552__B2 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08985_ net783 _04622_ _04623_ net713 vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__o211a_1
X_13848__18 clknet_leaf_166_clk vssd1 vssd1 vccd1 vccd1 net1487 sky130_fd_sc_hd__inv_2
XANTENNA_fanout484_A net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07936_ _03559_ _03574_ vssd1 vssd1 vccd1 vccd1 _03575_ sky130_fd_sc_hd__or2_4
XANTENNA__11304__B2 _06033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09552__A _05190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout651_A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11855__A2 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10698__A net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout272_X net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07867_ net952 _03500_ _03502_ _03505_ vssd1 vssd1 vccd1 vccd1 _03506_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout1393_A net1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout749_A net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09606_ net787 _05240_ _05241_ net741 vssd1 vssd1 vccd1 vccd1 _05245_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_108_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07798_ net628 _03435_ _03436_ net608 vssd1 vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__a31o_1
XANTENNA__11068__B1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09537_ top.CPU.registers.data\[193\] net835 net779 _05175_ vssd1 vssd1 vccd1 vccd1
+ _05176_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout916_A net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout537_X net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08484__A1 top.CPU.control_unit.instruction\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09468_ top.CPU.registers.data\[738\] net1393 net823 top.CPU.registers.data\[706\]
+ net723 vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__a221o_1
XFILLER_24_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09681__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08419_ _03924_ _04057_ vssd1 vssd1 vccd1 vccd1 _04058_ sky130_fd_sc_hd__nand2b_1
XFILLER_12_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout704_X net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09399_ net696 _05036_ _05037_ vssd1 vssd1 vccd1 vccd1 _05038_ sky130_fd_sc_hd__or3_1
XFILLER_11_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11430_ net1401 _03189_ _06575_ vssd1 vssd1 vccd1 vccd1 _06717_ sky130_fd_sc_hd__or3_1
XANTENNA__09433__B1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10043__A1 _03315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11361_ net3203 net288 net284 _06449_ vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__a22o_1
XANTENNA__12852__S net1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10594__A2 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13100_ top.SPI.count\[1\] top.SPI.count\[0\] vssd1 vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__or2_1
X_10312_ _05943_ vssd1 vssd1 vccd1 vccd1 _05944_ sky130_fd_sc_hd__inv_2
XANTENNA__09727__A _05332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11292_ net357 vssd1 vssd1 vccd1 vccd1 _06705_ sky130_fd_sc_hd__inv_2
XFILLER_153_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08631__A net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11468__S net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08539__A2 net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13031_ top.SPI.parameters\[17\] top.SPI.paroutput\[9\] net1357 vssd1 vssd1 vccd1
+ vccd1 _07441_ sky130_fd_sc_hd__mux2_1
X_10243_ net602 _05876_ _05877_ vssd1 vssd1 vccd1 vccd1 _05878_ sky130_fd_sc_hd__a21oi_4
XANTENNA__13532__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11695__C net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11543__A1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07747__B1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_52 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08944__C1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1102 net1103 vssd1 vssd1 vccd1 vccd1 net1102 sky130_fd_sc_hd__clkbuf_4
X_10174_ net515 _05810_ vssd1 vssd1 vccd1 vccd1 _05811_ sky130_fd_sc_hd__and2_1
XFILLER_160_390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1113 net1147 vssd1 vssd1 vccd1 vccd1 net1113 sky130_fd_sc_hd__clkbuf_4
XFILLER_152_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1124 net1127 vssd1 vssd1 vccd1 vccd1 net1124 sky130_fd_sc_hd__clkbuf_4
Xfanout1135 net1136 vssd1 vssd1 vccd1 vccd1 net1135 sky130_fd_sc_hd__clkbuf_4
XANTENNA__15236__RESET_B net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1146 net1147 vssd1 vssd1 vccd1 vccd1 net1146 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_128_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14982_ clknet_leaf_98_clk _01227_ net1254 vssd1 vssd1 vccd1 vccd1 top.SPI.paroutput\[21\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1157 net1170 vssd1 vssd1 vccd1 vccd1 net1157 sky130_fd_sc_hd__buf_2
XANTENNA__08777__S net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12099__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1168 net1169 vssd1 vssd1 vccd1 vccd1 net1168 sky130_fd_sc_hd__buf_2
Xfanout170 net171 vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__buf_6
Xfanout1179 net1205 vssd1 vssd1 vccd1 vccd1 net1179 sky130_fd_sc_hd__buf_2
Xfanout181 _06777_ vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__buf_4
XANTENNA__09462__A net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout192 net193 vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__clkbuf_8
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13862__32 clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 net1501 sky130_fd_sc_hd__inv_2
XANTENNA__08078__A _03716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14146__316 clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 net1785 sky130_fd_sc_hd__inv_2
X_15603_ net1937 _01813_ net1184 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[403\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11059__B1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12815_ _07251_ _07257_ _07264_ _07266_ vssd1 vssd1 vccd1 vccd1 _07268_ sky130_fd_sc_hd__o22a_1
XFILLER_34_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11216__B net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13795_ net25 net1052 net887 net4010 vssd1 vssd1 vccd1 vccd1 _02676_ sky130_fd_sc_hd__a22o_1
XANTENNA__09121__C1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15534_ net1868 _01744_ net1104 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[334\]
+ sky130_fd_sc_hd__dfrtp_1
X_12746_ _07203_ _07204_ vssd1 vssd1 vccd1 vccd1 _07205_ sky130_fd_sc_hd__nand2_1
XANTENNA__08475__A1 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07710__A top.CPU.control_unit.instruction\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10282__A1 _05793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15465_ net1799 _01675_ net1055 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[265\]
+ sky130_fd_sc_hd__dfrtp_1
X_12677_ top.CPU.alu.program_counter\[2\] top.CPU.alu.program_counter\[3\] top.CPU.alu.program_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _07143_ sky130_fd_sc_hd__a21oi_1
XANTENNA__16024__RESET_B net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11232__A net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11628_ net563 _06598_ vssd1 vssd1 vccd1 vccd1 _06755_ sky130_fd_sc_hd__nor2_1
X_15396_ net1730 _01606_ net1210 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[196\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08017__S net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08322__S1 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08778__A2 net1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11559_ net3018 net248 _06741_ net488 vssd1 vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__a22o_1
XFILLER_144_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold607 top.CPU.addressnew\[20\] vssd1 vssd1 vccd1 vccd1 net3164 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07856__S net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold618 top.CPU.registers.data\[811\] vssd1 vssd1 vccd1 vccd1 net3175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold629 top.CPU.registers.data\[194\] vssd1 vssd1 vccd1 vccd1 net3186 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_170_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16017_ net2351 _02227_ net1189 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[817\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_90_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13229_ _02755_ _02792_ vssd1 vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_90_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1307 top.CPU.registers.data\[884\] vssd1 vssd1 vccd1 vccd1 net3864 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1318 top.mmio.mem_data_i\[26\] vssd1 vssd1 vccd1 vccd1 net3875 sky130_fd_sc_hd__dlygate4sd3_1
X_08770_ top.CPU.registers.data\[972\] net1316 net847 top.CPU.registers.data\[1004\]
+ net718 vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__a221o_1
XFILLER_84_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08687__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1329 top.CPU.registers.data\[98\] vssd1 vssd1 vccd1 vccd1 net3886 sky130_fd_sc_hd__dlygate4sd3_1
X_07721_ net923 _03358_ _03359_ net628 vssd1 vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__o211a_1
XANTENNA__09360__C1 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07652_ net1038 _03288_ _03289_ _03290_ vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__a211oi_4
XFILLER_92_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07910__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11126__B net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07583_ net779 _03220_ _03221_ net731 vssd1 vssd1 vccd1 vccd1 _03222_ sky130_fd_sc_hd__a211o_1
X_09322_ top.CPU.registers.data\[260\] net1329 net860 top.CPU.registers.data\[292\]
+ net696 vssd1 vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__a221o_1
XFILLER_34_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10965__B _05933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09253_ _04891_ vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__inv_2
XANTENNA__11470__B1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout232_A _06772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08204_ net937 _03841_ _03842_ net954 vssd1 vssd1 vccd1 vccd1 _03843_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_32_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09184_ net790 _04820_ _04821_ _04822_ net692 vssd1 vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__a311o_1
X_08135_ top.CPU.registers.data\[757\] net1381 net991 top.CPU.registers.data\[725\]
+ net916 vssd1 vssd1 vccd1 vccd1 _03774_ sky130_fd_sc_hd__a221o_1
XANTENNA__08769__A2 net1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10981__A _03167_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07977__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11796__B net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08066_ net932 _03703_ _03704_ net952 vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__o211a_1
XFILLER_146_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09718__A1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout699_A net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09179__C1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14290__460 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 net1929 sky130_fd_sc_hd__inv_2
XANTENNA__10328__A2 _05958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1406_A net1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07729__B1 _03342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11525__A1 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14587__757 clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 net2226 sky130_fd_sc_hd__inv_2
XFILLER_0_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout866_A net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout487_X net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12701__A top.CPU.alu.program_counter\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08968_ top.CPU.registers.data\[681\] top.CPU.registers.data\[649\] net805 vssd1
+ vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__mux2_1
XANTENNA__09282__A _04891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_162_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07919_ net683 _03553_ _03554_ _03557_ net614 vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_162_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14628__798 clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 net2267 sky130_fd_sc_hd__inv_2
XANTENNA__11828__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08154__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08899_ top.CPU.registers.data\[586\] net1313 net844 top.CPU.registers.data\[618\]
+ net765 vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout654_X net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1396_X net1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10930_ net659 _06354_ net436 vssd1 vssd1 vccd1 vccd1 _06512_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_123_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07901__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10861_ net524 _06466_ vssd1 vssd1 vccd1 vccd1 _06468_ sky130_fd_sc_hd__or2_1
XFILLER_72_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout821_X net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09103__C1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout919_X net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12600_ _03139_ top.SPI.count\[3\] _07100_ vssd1 vssd1 vccd1 vccd1 _07101_ sky130_fd_sc_hd__a21oi_1
XFILLER_140_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13580_ top.CPU.alu.program_counter\[12\] net1350 net582 vssd1 vssd1 vccd1 vccd1
+ _03015_ sky130_fd_sc_hd__o21a_1
XFILLER_71_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10792_ _05124_ _05270_ _06402_ vssd1 vssd1 vccd1 vccd1 _06403_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10264__A1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11461__A0 _06253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07530__A top.CPU.control_unit.instruction\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12531_ _07031_ _07032_ _07039_ _07021_ vssd1 vssd1 vccd1 vccd1 _07040_ sky130_fd_sc_hd__a22o_1
XFILLER_9_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10367__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15250_ net1584 _01460_ net1099 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_157_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12462_ net448 _05428_ vssd1 vssd1 vccd1 vccd1 _06971_ sky130_fd_sc_hd__or2_1
XANTENNA__09957__A1 _03650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11213__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11413_ _06547_ net279 net268 net2964 vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__a22o_1
XFILLER_172_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09728__Y _05367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15181_ net1518 _01391_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r1_prev\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_12393_ _06922_ _06925_ _06927_ _06930_ vssd1 vssd1 vccd1 vccd1 _06931_ sky130_fd_sc_hd__nor4b_1
XFILLER_138_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10891__A net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10567__A2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12961__B1 net1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14531__701 clknet_leaf_170_clk vssd1 vssd1 vccd1 vccd1 net2170 sky130_fd_sc_hd__inv_2
XANTENNA__08090__C1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11344_ net3598 net286 net277 _06107_ vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__a22o_1
XFILLER_99_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11275_ net522 _06565_ vssd1 vssd1 vccd1 vccd1 _06695_ sky130_fd_sc_hd__nor2_1
XFILLER_165_84 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08917__C1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_148_Right_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13014_ net2690 _07432_ net895 vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__mux2_1
XFILLER_140_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10226_ net395 net308 _05654_ _05860_ vssd1 vssd1 vccd1 vccd1 _05861_ sky130_fd_sc_hd__a31oi_2
XFILLER_3_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10115__B _05643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10157_ _05792_ _05793_ net224 vssd1 vssd1 vccd1 vccd1 _05794_ sky130_fd_sc_hd__a21o_1
XFILLER_121_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13269__B2 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold4 top.CPU.registers.data_out_r1_prev\[0\] vssd1 vssd1 vccd1 vccd1 net2561 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10088_ _05725_ vssd1 vssd1 vccd1 vccd1 _05726_ sky130_fd_sc_hd__inv_2
X_14965_ clknet_leaf_97_clk net3439 net1248 vssd1 vssd1 vccd1 vccd1 top.SPI.paroutput\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08145__A0 _03783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09342__C1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08448__A1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13778_ net6 net1049 net884 net3850 vssd1 vssd1 vccd1 vccd1 _02659_ sky130_fd_sc_hd__o22a_1
XFILLER_31_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15517_ net1851 _01727_ net1122 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[317\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_148_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12729_ _07189_ _07188_ net127 vssd1 vssd1 vccd1 vccd1 _07190_ sky130_fd_sc_hd__mux2_1
X_16497_ clknet_leaf_41_clk _02659_ net1115 vssd1 vssd1 vccd1 vccd1 top.mmio.mem_data_i\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_148_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15448_ net1782 _01658_ net1148 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[248\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11204__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15379_ net1713 _01589_ net1187 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[179\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_129_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12952__A0 _07391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07959__B1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold404 top.SPI.paroutput\[28\] vssd1 vssd1 vccd1 vccd1 net2961 sky130_fd_sc_hd__dlygate4sd3_1
Xhold415 _02696_ vssd1 vssd1 vccd1 vccd1 net2972 sky130_fd_sc_hd__dlygate4sd3_1
X_14274__444 clknet_leaf_143_clk vssd1 vssd1 vccd1 vccd1 net1913 sky130_fd_sc_hd__inv_2
XFILLER_171_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold426 top.CPU.registers.data\[989\] vssd1 vssd1 vccd1 vccd1 net2983 sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 top.SPI.paroutput\[25\] vssd1 vssd1 vccd1 vccd1 net2994 sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 top.CPU.registers.data\[281\] vssd1 vssd1 vccd1 vccd1 net3005 sky130_fd_sc_hd__dlygate4sd3_1
X_09940_ _03723_ _03789_ vssd1 vssd1 vccd1 vccd1 _05579_ sky130_fd_sc_hd__nand2_1
Xhold459 top.CPU.registers.data\[271\] vssd1 vssd1 vccd1 vccd1 net3016 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10306__A net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11507__A1 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_115_Right_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09176__A2 net1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout906 net909 vssd1 vssd1 vccd1 vccd1 net906 sky130_fd_sc_hd__buf_2
X_09871_ _03476_ _03509_ vssd1 vssd1 vccd1 vccd1 _05510_ sky130_fd_sc_hd__nand2_1
Xfanout917 net918 vssd1 vssd1 vccd1 vccd1 net917 sky130_fd_sc_hd__clkbuf_4
Xfanout928 net929 vssd1 vssd1 vccd1 vccd1 net928 sky130_fd_sc_hd__clkbuf_4
X_14315__485 clknet_leaf_134_clk vssd1 vssd1 vccd1 vccd1 net1954 sky130_fd_sc_hd__inv_2
Xfanout939 net942 vssd1 vssd1 vccd1 vccd1 net939 sky130_fd_sc_hd__clkbuf_4
XFILLER_97_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12180__A1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08822_ net689 _04459_ _04432_ vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09581__C1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1104 top.CPU.registers.data\[668\] vssd1 vssd1 vccd1 vccd1 net3661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1115 top.SPI.paroutput\[22\] vssd1 vssd1 vccd1 vccd1 net3672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1126 top.CPU.registers.data\[268\] vssd1 vssd1 vccd1 vccd1 net3683 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1137 top.CPU.registers.data\[950\] vssd1 vssd1 vccd1 vccd1 net3694 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08753_ net1398 _03160_ _03985_ vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__o21a_1
Xhold1148 top.CPU.registers.data\[374\] vssd1 vssd1 vccd1 vccd1 net3705 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08136__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout182_A _06777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1159 top.CPU.registers.data\[993\] vssd1 vssd1 vccd1 vccd1 net3716 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07704_ top.CPU.control_unit.instruction\[24\] net685 vssd1 vssd1 vccd1 vccd1 _03343_
+ sky130_fd_sc_hd__nand2_1
XFILLER_94_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10041__A net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08687__A1 _04325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08684_ _03342_ _04309_ _04322_ vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__o21ai_2
XANTENNA__10494__A1 _05733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07635_ _03151_ _03162_ net1033 vssd1 vssd1 vccd1 vccd1 _03274_ sky130_fd_sc_hd__nand3_1
XANTENNA__11691__B1 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07895__C1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10976__A net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12235__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07566_ net1048 _03164_ net1039 top.CPU.control_unit.instruction\[16\] vssd1 vssd1
+ vccd1 vccd1 _03205_ sky130_fd_sc_hd__o31a_1
X_09305_ top.CPU.registers.data_out_r2_prev\[4\] net687 net620 _04936_ _04943_ vssd1
+ vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__o2111ai_2
XANTENNA__09100__A2 net1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07497_ net1353 vssd1 vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout235_X net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout614_A net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1356_A top.SPI.state\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09236_ net739 _04871_ _04874_ _04868_ vssd1 vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__a31o_1
XFILLER_10_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold1464_A top.CPU.registers.data_out_r1_prev\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout402_X net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09167_ top.CPU.registers.data\[38\] top.CPU.registers.data\[6\] net815 vssd1 vssd1
+ vccd1 vccd1 _04806_ sky130_fd_sc_hd__mux2_1
XANTENNA__12943__A0 top.CPU.alu.program_counter\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10549__A2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15581__RESET_B net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08118_ top.CPU.registers.data\[565\] top.CPU.registers.data\[533\] net992 vssd1
+ vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__mux2_1
XFILLER_79_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08072__C1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08181__A _03819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09098_ top.CPU.registers.data\[71\] net1332 net864 top.CPU.registers.data\[103\]
+ net778 vssd1 vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout983_A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08049_ top.CPU.registers.data\[180\] net1008 net905 vssd1 vssd1 vccd1 vccd1 _03688_
+ sky130_fd_sc_hd__a21o_1
XFILLER_123_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13499__A1 top.CPU.data_out\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1311_X net1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold960 top.CPU.registers.data\[232\] vssd1 vssd1 vccd1 vccd1 net3517 sky130_fd_sc_hd__dlygate4sd3_1
Xhold971 top.CPU.registers.data\[879\] vssd1 vssd1 vccd1 vccd1 net3528 sky130_fd_sc_hd__dlygate4sd3_1
X_11060_ net143 net535 vssd1 vssd1 vccd1 vccd1 _06587_ sky130_fd_sc_hd__and2_1
Xhold982 top.CPU.registers.data\[275\] vssd1 vssd1 vccd1 vccd1 net3539 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_164_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold993 top.CPU.registers.data\[355\] vssd1 vssd1 vccd1 vccd1 net3550 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout771_X net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10011_ _05646_ _05649_ net389 vssd1 vssd1 vccd1 vccd1 _05650_ sky130_fd_sc_hd__mux2_1
XFILLER_135_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13527__A _03915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08914__A2 net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09324__C1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08222__S0 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11962_ net519 _06510_ net350 _06776_ vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__a31o_1
XANTENNA__08678__A1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13701_ _03054_ net3474 vssd1 vssd1 vccd1 vccd1 _02622_ sky130_fd_sc_hd__nor2_1
XFILLER_17_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10913_ _06213_ net435 vssd1 vssd1 vccd1 vccd1 _06502_ sky130_fd_sc_hd__and2_1
XANTENNA__11682__B1 net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07886__C1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11893_ net147 net3546 net190 vssd1 vssd1 vccd1 vccd1 _01670_ sky130_fd_sc_hd__mux2_1
X_16420_ clknet_leaf_57_clk _00002_ net1145 vssd1 vssd1 vccd1 vccd1 top.I2C.I2C_state\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09627__A0 top.CPU.alu.program_counter\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13632_ net3039 _07144_ net664 vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__mux2_1
XANTENNA__07531__Y _03170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10844_ net377 _05266_ vssd1 vssd1 vccd1 vccd1 _06452_ sky130_fd_sc_hd__nor2_1
XANTENNA__12226__A2 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11434__A0 _05808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16351_ clknet_leaf_68_clk _02560_ net1167 vssd1 vssd1 vccd1 vccd1 top.CPU.addressnew\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_158_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_4_11_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13563_ top.CPU.addressnew\[5\] net579 _03003_ _03004_ vssd1 vssd1 vccd1 vccd1 _02535_
+ sky130_fd_sc_hd__a22o_1
X_10775_ _05545_ _05554_ _04991_ vssd1 vssd1 vccd1 vccd1 _06387_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15302_ net1636 _01512_ net1074 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[102\]
+ sky130_fd_sc_hd__dfrtp_1
X_12514_ _07017_ _07019_ _07020_ vssd1 vssd1 vccd1 vccd1 _07023_ sky130_fd_sc_hd__o21ai_1
X_16282_ clknet_leaf_62_clk _02492_ net1161 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.toreg\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13494_ _03108_ _03200_ _03263_ vssd1 vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__nor3_2
X_14258__428 clknet_leaf_201_clk vssd1 vssd1 vccd1 vccd1 net1897 sky130_fd_sc_hd__inv_2
X_15233_ net1567 _01443_ net1230 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[33\]
+ sky130_fd_sc_hd__dfrtp_1
X_12445_ net1339 top.I2C.output_state\[2\] net3543 vssd1 vssd1 vccd1 vccd1 _06959_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_138_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09187__A net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15164_ clknet_leaf_62_clk _01374_ net1161 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.readout
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08063__C1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12376_ top.I2C.byte_manager_state\[2\] _06914_ _06915_ top.I2C.byte_manager_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00041_ sky130_fd_sc_hd__a22o_1
XFILLER_126_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14002__172 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 net1641 sky130_fd_sc_hd__inv_2
XFILLER_141_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07810__C1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11327_ net3071 net292 _06711_ net495 vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__a22o_1
XFILLER_126_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15095_ net1477 _01308_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r2_prev\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11258_ net514 _06553_ vssd1 vssd1 vccd1 vccd1 _06685_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09563__C1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10209_ net512 _05611_ _05844_ _05843_ _05813_ vssd1 vssd1 vccd1 vccd1 _05845_ sky130_fd_sc_hd__a311o_1
X_11189_ net3706 net299 _06653_ net325 vssd1 vssd1 vccd1 vccd1 _02259_ sky130_fd_sc_hd__a22o_1
XANTENNA__10712__A2 _06317_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12060__B net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15997_ net2331 _02207_ net1119 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[797\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_76_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14948_ clknet_leaf_62_clk _01194_ net1163 vssd1 vssd1 vccd1 vccd1 top.CPU.alu.program_counter\[31\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08669__A1 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08965__S net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07877__C1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16618_ net1347 vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07892__A2 net1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14700__870 clknet_leaf_195_clk vssd1 vssd1 vccd1 vccd1 net2339 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10228__A1 _03315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16549_ clknet_4_15_0_clk _02711_ net1263 vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10228__B2 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11425__B1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09021_ top.CPU.control_unit.instruction\[29\] _04596_ _04597_ vssd1 vssd1 vccd1
+ vccd1 _04660_ sky130_fd_sc_hd__o21a_1
XFILLER_129_471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold201 top.CPU.registers.data\[9\] vssd1 vssd1 vccd1 vccd1 net2758 sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 top.SPI.paroutput\[11\] vssd1 vssd1 vccd1 vccd1 net2769 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold223 top.I2C.I2C_state\[5\] vssd1 vssd1 vccd1 vccd1 net2780 sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 top.I2C.output_state\[5\] vssd1 vssd1 vccd1 vccd1 net2791 sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 net93 vssd1 vssd1 vccd1 vccd1 net2802 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold256 top.CPU.registers.data\[912\] vssd1 vssd1 vccd1 vccd1 net2813 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold267 top.CPU.registers.data\[563\] vssd1 vssd1 vccd1 vccd1 net2824 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09384__X _05023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold278 top.CPU.registers.data\[729\] vssd1 vssd1 vccd1 vccd1 net2835 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09923_ _05541_ _05561_ vssd1 vssd1 vccd1 vccd1 _05562_ sky130_fd_sc_hd__nand2_1
XANTENNA__09149__A2 net1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09825__A net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout703 _03212_ vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__clkbuf_4
Xhold289 top.CPU.registers.data\[830\] vssd1 vssd1 vccd1 vccd1 net2846 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout714 net736 vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__clkbuf_4
XFILLER_160_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13350__A0 top.CPU.control_unit.instruction\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout397_A net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout725 net735 vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__clkbuf_2
Xfanout736 _03209_ vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__clkbuf_4
Xfanout747 net760 vssd1 vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__buf_2
X_09854_ top.CPU.registers.data\[346\] net1305 net1028 top.CPU.registers.data\[378\]
+ net945 vssd1 vssd1 vccd1 vccd1 _05493_ sky130_fd_sc_hd__a221o_1
Xfanout758 net759 vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1104_A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout769 net770 vssd1 vssd1 vccd1 vccd1 net769 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_142_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08805_ net952 _04440_ net625 vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__a21o_1
XFILLER_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09785_ net679 _05404_ _05405_ _05423_ net607 vssd1 vssd1 vccd1 vccd1 _05424_ sky130_fd_sc_hd__a311o_1
XFILLER_58_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout564_A net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08109__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout185_X net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_0_Left_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_192_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09306__C1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08736_ top.CPU.registers.data\[205\] net1371 net967 top.CPU.registers.data\[237\]
+ net926 vssd1 vssd1 vccd1 vccd1 _04375_ sky130_fd_sc_hd__o221a_1
XANTENNA__12456__A2 _03439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08875__S net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_72_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11664__B1 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14699__869 clknet_leaf_149_clk vssd1 vssd1 vccd1 vccd1 net2338 sky130_fd_sc_hd__inv_2
X_08667_ top.CPU.registers.data\[206\] net1376 net981 top.CPU.registers.data\[238\]
+ net934 vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout731_A net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout352_X net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout829_A net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07618_ top.CPU.control_unit.instruction\[28\] top.CPU.control_unit.instruction\[27\]
+ top.CPU.control_unit.instruction\[29\] net1363 vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__or4_1
XFILLER_53_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12208__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08598_ top.CPU.registers.data\[207\] net1375 net974 top.CPU.registers.data\[239\]
+ net929 vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__o221a_1
XANTENNA__07883__A2 net1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11416__B1 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09085__A1 net1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07549_ top.CPU.control_unit.instruction\[11\] net648 _03184_ vssd1 vssd1 vccd1 vccd1
+ _03188_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_87_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout617_X net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1359_X net1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10560_ net415 _06180_ _06181_ vssd1 vssd1 vccd1 vccd1 _06182_ sky130_fd_sc_hd__o21ba_1
XANTENNA__11033__C net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08904__A net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_130_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09219_ _04857_ vssd1 vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__inv_2
XFILLER_154_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10491_ _04125_ net509 net503 _05291_ vssd1 vssd1 vccd1 vccd1 _06116_ sky130_fd_sc_hd__o22ai_1
XTAP_TAPCELL_ROW_118_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13021__S net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10872__C net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12230_ net3872 net654 _06881_ vssd1 vssd1 vccd1 vccd1 _01446_ sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_10_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout986_X net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11195__A2 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12161_ net3941 net645 _06848_ vssd1 vssd1 vccd1 vccd1 _01482_ sky130_fd_sc_hd__o21a_1
XFILLER_146_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_145_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11112_ net574 net530 _06010_ vssd1 vssd1 vccd1 vccd1 _06614_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_131_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08348__A0 _03984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12092_ net3956 net645 _06814_ vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__o21a_1
Xhold790 top.CPU.registers.data\[593\] vssd1 vssd1 vccd1 vccd1 net3347 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_25_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11329__X _06712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15920_ net2254 _02130_ net1154 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[720\]
+ sky130_fd_sc_hd__dfrtp_1
X_11043_ net3848 net368 _06580_ net320 vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__a22o_1
XANTENNA__16550__RESET_B net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15851_ net2185 _02061_ net1065 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[651\]
+ sky130_fd_sc_hd__dfrtp_1
X_14643__813 clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 net2282 sky130_fd_sc_hd__inv_2
XFILLER_65_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_3_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_3_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_92_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15782_ net2116 _01992_ net1074 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[582\]
+ sky130_fd_sc_hd__dfrtp_1
X_12994_ net1357 net1410 _07422_ vssd1 vssd1 vccd1 vccd1 _07423_ sky130_fd_sc_hd__or3b_1
XFILLER_17_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10458__A1 _06082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11945_ net520 _06488_ net351 _06774_ vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__a31o_1
XANTENNA__11655__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07859__C1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11876_ _06033_ net3248 net190 vssd1 vssd1 vccd1 vccd1 _01687_ sky130_fd_sc_hd__mux2_1
XANTENNA__11670__A3 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16403_ clknet_leaf_57_clk _00074_ net1162 vssd1 vssd1 vccd1 vccd1 top.wm.curr_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_13615_ top.CPU.alu.program_counter\[26\] _05904_ net1351 vssd1 vssd1 vccd1 vccd1
+ _03036_ sky130_fd_sc_hd__mux2_1
XANTENNA__11407__B1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10827_ net549 _05195_ _06434_ _06435_ vssd1 vssd1 vccd1 vccd1 _06436_ sky130_fd_sc_hd__o211a_1
XANTENNA__11224__B net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16334_ clknet_leaf_68_clk _02543_ net1167 vssd1 vssd1 vccd1 vccd1 top.CPU.addressnew\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_158_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13546_ net1353 top.CPU.done top.CPU.handler.state\[0\] vssd1 vssd1 vccd1 vccd1 _02993_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12080__B1 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08823__A1 net1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10758_ _05557_ _06370_ _06369_ _06359_ vssd1 vssd1 vccd1 vccd1 _06371_ sky130_fd_sc_hd__o211a_2
XTAP_TAPCELL_ROW_41_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10630__A1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11511__Y _06734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16265_ clknet_leaf_44_clk _02475_ net1126 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.toreg\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_13477_ net1397 net872 _02927_ net419 vssd1 vssd1 vccd1 vccd1 _02960_ sky130_fd_sc_hd__a31o_1
XANTENNA__10555__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10689_ _04797_ _05276_ _04732_ vssd1 vssd1 vccd1 vccd1 _06305_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11240__A net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15216_ net1550 _01426_ net1234 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_12428_ top.I2C.initiate_read_bit _06903_ _06905_ net1054 top.I2C.output_state\[28\]
+ vssd1 vssd1 vccd1 vccd1 _00059_ sky130_fd_sc_hd__a32o_1
XFILLER_127_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08036__C1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16196_ net2530 _02406_ net1212 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[996\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_154_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15147_ clknet_leaf_48_clk _01357_ net1130 vssd1 vssd1 vccd1 vccd1 top.I2C.data_out\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09784__C1 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12359_ top.I2C.byte_manager_state\[2\] _06901_ vssd1 vssd1 vccd1 vccd1 _06902_ sky130_fd_sc_hd__or2_1
XFILLER_142_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08820__Y _04459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10933__A2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15078_ clknet_leaf_49_clk _00056_ net1129 vssd1 vssd1 vccd1 vccd1 top.I2C.output_state\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_39_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09000__A1 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09551__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14386__556 clknet_leaf_201_clk vssd1 vssd1 vccd1 vccd1 net2025 sky130_fd_sc_hd__inv_2
X_09570_ _05207_ _05208_ net611 vssd1 vssd1 vccd1 vccd1 _05209_ sky130_fd_sc_hd__a21o_1
XANTENNA__11118__C net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10449__A1 _03315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09380__A _05018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08521_ top.CPU.registers.data\[304\] top.CPU.registers.data\[272\] net984 vssd1
+ vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__mux2_1
XANTENNA__11646__B1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14427__597 clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 net2066 sky130_fd_sc_hd__inv_2
XANTENNA__08511__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08452_ _04090_ vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__inv_2
XANTENNA__12010__S net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07865__A2 net1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1030 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08383_ top.CPU.registers.data\[178\] top.CPU.registers.data\[146\] top.CPU.registers.data\[50\]
+ top.CPU.registers.data\[18\] net982 net908 vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout145_A _06270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09379__X _05018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12071__B1 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08814__A1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08275__C1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10621__A1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08290__A2 net1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout312_A net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09004_ top.CPU.registers.data\[873\] top.CPU.registers.data\[841\] net965 vssd1
+ vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_152_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13571__A0 top.CPU.alu.program_counter\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1221_A net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10924__A2 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1319_A net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13994__164 clknet_leaf_148_clk vssd1 vssd1 vccd1 vccd1 net1633 sky130_fd_sc_hd__inv_2
X_14330__500 clknet_leaf_163_clk vssd1 vssd1 vccd1 vccd1 net1969 sky130_fd_sc_hd__inv_2
XFILLER_78_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout500 _06755_ vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__buf_6
XANTENNA_fanout681_A net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout511 _05520_ vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__buf_4
XFILLER_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout779_A net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09906_ _05544_ vssd1 vssd1 vccd1 vccd1 _05545_ sky130_fd_sc_hd__inv_2
Xfanout522 net523 vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10053__X _05692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout533 _03196_ vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__buf_4
XANTENNA__10137__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12677__A2 top.CPU.alu.program_counter\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout544 _06523_ vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__buf_4
Xfanout555 net556 vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__buf_2
XANTENNA__11228__A_N _05933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout566 net569 vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__buf_2
XANTENNA__11885__A0 _06230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09837_ top.CPU.registers.data\[762\] net1384 net1001 top.CPU.registers.data\[730\]
+ net921 vssd1 vssd1 vccd1 vccd1 _05476_ sky130_fd_sc_hd__a221o_1
XFILLER_59_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout577 _03169_ vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__clkbuf_4
XFILLER_101_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout588 net589 vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10213__B net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout946_A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout567_X net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08750__B1 _03342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11028__C net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09768_ top.CPU.registers.data\[987\] net1298 net1019 top.CPU.registers.data\[1019\]
+ net915 vssd1 vssd1 vccd1 vccd1 _05407_ sky130_fd_sc_hd__a221o_1
XFILLER_132_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07803__A _03407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08719_ net784 _04354_ _04355_ net714 vssd1 vssd1 vccd1 vccd1 _04358_ sky130_fd_sc_hd__o211a_1
XANTENNA__11637__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ top.CPU.registers.data\[985\] net1306 net1029 top.CPU.registers.data\[1017\]
+ net922 vssd1 vssd1 vccd1 vccd1 _05338_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout734_X net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11101__A2 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08502__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11730_ _06577_ net207 net194 net3817 vssd1 vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__a22o_1
XFILLER_26_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11044__B net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11661_ _06465_ net198 net424 net3348 vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout901_X net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13400_ net890 _02917_ vssd1 vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_54_Left_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10612_ net439 _06231_ vssd1 vssd1 vccd1 vccd1 _06232_ sky130_fd_sc_hd__nand2_1
XANTENNA__07608__A2 net1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08805__A1 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08266__C1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12062__B1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11592_ net648 net360 vssd1 vssd1 vccd1 vccd1 _06751_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_172_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13331_ top.CPU.control_unit.instruction\[6\] _02867_ net669 vssd1 vssd1 vccd1 vccd1
+ _02440_ sky130_fd_sc_hd__mux2_1
XFILLER_10_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11331__Y _06713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10543_ _05673_ _06141_ _06164_ net407 _06165_ vssd1 vssd1 vccd1 vccd1 _06166_ sky130_fd_sc_hd__o221a_1
XFILLER_127_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11060__A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16050_ net2384 _02260_ net1098 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[850\]
+ sky130_fd_sc_hd__dfrtp_1
X_13262_ net891 top.I2C.data_out\[5\] _02785_ vssd1 vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__mux2_1
XFILLER_109_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08018__C1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10474_ _06092_ _06096_ _06097_ _06099_ vssd1 vssd1 vccd1 vccd1 _06100_ sky130_fd_sc_hd__or4_2
X_15001_ clknet_leaf_96_clk _01246_ net1248 vssd1 vssd1 vccd1 vccd1 top.SPI.parameters\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13562__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09766__C1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12213_ net3865 net646 _06873_ vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__o21a_1
XFILLER_123_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13193_ top.I2C.which_data_address\[0\] _02772_ vssd1 vssd1 vccd1 vccd1 _02773_ sky130_fd_sc_hd__and2b_2
XANTENNA__12003__A_N net1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09465__A net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12144_ top.CPU.registers.data\[80\] net174 vssd1 vssd1 vccd1 vccd1 _06840_ sky130_fd_sc_hd__and2_1
XFILLER_151_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14073__243 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 net1712 sky130_fd_sc_hd__inv_2
XANTENNA__07792__A1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Left_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10128__B1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12075_ top.CPU.registers.data\[115\] net651 vssd1 vssd1 vccd1 vccd1 _06806_ sky130_fd_sc_hd__or2_1
XFILLER_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11876__A0 _06033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15903_ net2237 _02113_ net1220 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[703\]
+ sky130_fd_sc_hd__dfrtp_1
X_11026_ net531 _06570_ vssd1 vssd1 vccd1 vccd1 _06571_ sky130_fd_sc_hd__nor2_1
XANTENNA__10123__B net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11340__A2 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14114__284 clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 net1753 sky130_fd_sc_hd__inv_2
XFILLER_49_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15834_ net2168 _02044_ net1244 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[634\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_64_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08809__A net1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12977_ top.I2C.bit_timer_counter\[3\] top.I2C.bit_timer_counter\[4\] _07407_ vssd1
+ vssd1 vccd1 vccd1 _07411_ sky130_fd_sc_hd__and3_1
XANTENNA__09297__A1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15765_ net2099 _01975_ net1228 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[565\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15684__RESET_B net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11928_ net3707 net185 net348 _06393_ vssd1 vssd1 vccd1 vccd1 _01638_ sky130_fd_sc_hd__a22o_1
XANTENNA__07847__A2 net1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15696_ net2030 _01906_ net1108 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[496\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_75_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_72_Left_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12765__S net1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11859_ _06695_ net203 net154 net2852 vssd1 vssd1 vccd1 vccd1 _01702_ sky130_fd_sc_hd__a22o_1
XFILLER_159_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08257__C1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12053__B1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14771__941 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 net2410 sky130_fd_sc_hd__inv_2
XFILLER_9_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10603__A1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16317_ clknet_leaf_83_clk _02526_ net1263 vssd1 vssd1 vccd1 vccd1 top.CPU.data_out\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_13529_ _03854_ net584 vssd1 vssd1 vccd1 vccd1 _02985_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_97_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16248_ clknet_leaf_60_clk _02458_ net1139 vssd1 vssd1 vccd1 vccd1 top.CPU.control_unit.instruction\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_11_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14812__982 clknet_leaf_139_clk vssd1 vssd1 vccd1 vccd1 net2451 sky130_fd_sc_hd__inv_2
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 SEL_O[3] sky130_fd_sc_hd__buf_2
X_13978__148 clknet_leaf_159_clk vssd1 vssd1 vccd1 vccd1 net1617 sky130_fd_sc_hd__inv_2
Xoutput114 net114 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
XANTENNA__10367__A0 _03822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16179_ net2513 _02389_ net1184 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[979\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_58_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_81_Left_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12513__B _04531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12108__A1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09509__C1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07952_ net793 _03584_ _03585_ net721 vssd1 vssd1 vccd1 vccd1 _03591_ sky130_fd_sc_hd__o211a_1
XFILLER_87_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12659__A2 _05232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11867__A0 _05808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09524__A2 net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_71_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07883_ top.CPU.registers.data\[860\] net1332 net863 top.CPU.registers.data\[892\]
+ net754 vssd1 vssd1 vccd1 vccd1 _03522_ sky130_fd_sc_hd__a221o_1
X_09622_ net788 _05251_ _05252_ vssd1 vssd1 vccd1 vccd1 _05261_ sky130_fd_sc_hd__and3_1
XANTENNA__13608__A1 top.CPU.alu.program_counter\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11619__A0 _06311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09553_ net880 _05190_ _05159_ vssd1 vssd1 vccd1 vccd1 _05192_ sky130_fd_sc_hd__o21ai_4
XANTENNA__11145__A net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08504_ top.CPU.registers.data\[848\] net1321 net852 top.CPU.registers.data\[880\]
+ net745 vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__a221o_1
XANTENNA__11095__A1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_90_Left_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09484_ net1034 _05120_ _05122_ vssd1 vssd1 vccd1 vccd1 _05123_ sky130_fd_sc_hd__a21oi_2
XANTENNA__08496__C1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08435_ net697 _04072_ _04073_ vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__or3_1
XFILLER_23_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10984__A net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout148_X net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1171_A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout527_A net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12044__B1 _06781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08366_ top.CPU.registers.data\[178\] top.CPU.registers.data\[146\] net818 vssd1
+ vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__mux2_1
XANTENNA__11799__B net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11398__A2 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13792__B1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14889__1059 clknet_leaf_154_clk vssd1 vssd1 vccd1 vccd1 net2528 sky130_fd_sc_hd__inv_2
XANTENNA__10048__X _05687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09460__A1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08297_ net707 _03934_ _03935_ vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout315_X net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11311__C _05694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09748__C1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10358__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14057__227 clknet_leaf_156_clk vssd1 vssd1 vccd1 vccd1 net1696 sky130_fd_sc_hd__inv_2
XFILLER_133_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12704__A top.CPU.alu.program_counter\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10190_ _05737_ _05825_ net309 vssd1 vssd1 vccd1 vccd1 _05826_ sky130_fd_sc_hd__mux2_1
XFILLER_2_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout684_X net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11570__A2 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1306 net1307 vssd1 vssd1 vccd1 vccd1 net1306 sky130_fd_sc_hd__clkbuf_4
Xfanout1317 net1323 vssd1 vssd1 vccd1 vccd1 net1317 sky130_fd_sc_hd__clkbuf_4
Xfanout330 _03048_ vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__buf_2
Xfanout1328 net1331 vssd1 vssd1 vccd1 vccd1 net1328 sky130_fd_sc_hd__clkbuf_4
Xfanout1339 net1342 vssd1 vssd1 vccd1 vccd1 net1339 sky130_fd_sc_hd__buf_2
Xfanout341 net343 vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__clkbuf_8
XFILLER_59_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout352 net353 vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11039__B net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11858__B1 net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout363 net364 vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout851_X net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout374 net375 vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout385 _05157_ vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__clkbuf_4
XFILLER_19_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11322__A2 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout949_X net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12900_ top.CPU.alu.program_counter\[25\] _07344_ net1362 vssd1 vssd1 vccd1 vccd1
+ _01188_ sky130_fd_sc_hd__mux2_1
Xfanout396 net397 vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__clkbuf_2
XFILLER_4_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13535__A _05498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09224__S net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07533__A net1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12831_ _07274_ _07282_ net126 vssd1 vssd1 vccd1 vccd1 _07283_ sky130_fd_sc_hd__mux2_1
XFILLER_36_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11055__A net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15550_ net1884 _01760_ net1237 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[350\]
+ sky130_fd_sc_hd__dfrtp_1
X_12762_ _07218_ _07219_ vssd1 vssd1 vccd1 vccd1 _07220_ sky130_fd_sc_hd__and2_1
XANTENNA__11086__B2 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11713_ _06550_ net200 net421 net2720 vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__a22o_1
X_15481_ net1815 _01691_ net1244 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[281\]
+ sky130_fd_sc_hd__dfrtp_1
X_12693_ top.CPU.alu.program_counter\[6\] _04856_ vssd1 vssd1 vccd1 vccd1 _07157_
+ sky130_fd_sc_hd__or2_1
XFILLER_43_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14755__925 clknet_leaf_170_clk vssd1 vssd1 vccd1 vccd1 net2394 sky130_fd_sc_hd__inv_2
X_11644_ _06127_ net205 net426 net3488 vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__a22o_1
XANTENNA__08239__C1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput16 DAT_I[22] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10597__A0 _04363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11575_ net2914 net246 _06745_ net478 vssd1 vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__a22o_1
XANTENNA__08254__A2 net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput27 DAT_I[3] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16102_ net2436 _02312_ net1080 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[902\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_167_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13314_ _02830_ _02854_ vssd1 vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__nor2_1
Xinput38 nrst vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_2
X_10526_ net551 net501 net146 vssd1 vssd1 vccd1 vccd1 _06150_ sky130_fd_sc_hd__or3b_1
XFILLER_7_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12338__A1 _05084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09739__C1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16033_ net2367 _02243_ net1243 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[833\]
+ sky130_fd_sc_hd__dfrtp_1
X_13245_ net891 top.I2C.data_out\[13\] _02785_ vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__mux2_1
XANTENNA__09907__B _05266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10457_ _06082_ _06083_ vssd1 vssd1 vccd1 vccd1 _06084_ sky130_fd_sc_hd__nand2_2
XANTENNA__10349__B1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13176_ _06911_ _02757_ _02758_ _02756_ net3989 vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__a32o_1
X_10388_ _03787_ net509 net504 _03786_ _06016_ vssd1 vssd1 vccd1 vccd1 _06017_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_36_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07765__A1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11561__A2 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12127_ net3957 net175 _06831_ _06483_ vssd1 vssd1 vccd1 vccd1 _01499_ sky130_fd_sc_hd__a22o_1
XANTENNA__10134__A net1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12052__C net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11849__B1 net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12058_ net477 _06608_ _06797_ net179 net3794 vssd1 vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__a32o_1
XFILLER_78_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12510__A1 _04291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08714__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11313__A2 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12510__B2 _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11009_ _06333_ net541 vssd1 vssd1 vccd1 vccd1 _06560_ sky130_fd_sc_hd__or2_1
XFILLER_37_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15817_ net2151 _02027_ net1056 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[617\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15748_ net2082 _01958_ net1219 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[548\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07730__X _03369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15679_ net2013 _01889_ net1219 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[479\]
+ sky130_fd_sc_hd__dfrtp_1
X_14498__668 clknet_leaf_146_clk vssd1 vssd1 vccd1 vccd1 net2137 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08220_ _03857_ _03858_ vssd1 vssd1 vccd1 vccd1 _03859_ sky130_fd_sc_hd__and2_2
XANTENNA__12026__A0 _06056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08151_ top.CPU.registers.data\[311\] top.CPU.registers.data\[279\] net823 vssd1
+ vssd1 vccd1 vccd1 _03790_ sky130_fd_sc_hd__mux2_1
XFILLER_158_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10052__A2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08082_ _03683_ _03718_ vssd1 vssd1 vccd1 vccd1 _03721_ sky130_fd_sc_hd__nor2_1
XANTENNA__10028__B _05665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13526__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09745__A2 net1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11552__A2 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08984_ top.CPU.registers.data\[329\] net1309 net840 top.CPU.registers.data\[361\]
+ net761 vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__a221o_1
XFILLER_87_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10760__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13829__B2 top.CPU.data_out\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1017_A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07935_ net628 _03565_ _03573_ vssd1 vssd1 vccd1 vccd1 _03574_ sky130_fd_sc_hd__and3_1
XFILLER_87_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10979__A net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11304__A2 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout477_A _03193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_748 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07866_ net674 _03503_ _03504_ net604 vssd1 vssd1 vccd1 vccd1 _03505_ sky130_fd_sc_hd__a31o_1
XANTENNA__10698__B net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09605_ net788 _05238_ _05239_ net717 vssd1 vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__o211a_1
XANTENNA__09044__S net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14442__612 clknet_leaf_152_clk vssd1 vssd1 vccd1 vccd1 net2081 sky130_fd_sc_hd__inv_2
XFILLER_43_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07797_ top.CPU.registers.data\[478\] net1303 net1025 top.CPU.registers.data\[510\]
+ net920 vssd1 vssd1 vccd1 vccd1 _03436_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout265_X net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1386_A net1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11068__A1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14739__909 clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 net2378 sky130_fd_sc_hd__inv_2
X_09536_ top.CPU.registers.data\[225\] net1395 vssd1 vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__and2_1
XANTENNA__10815__A1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09467_ top.CPU.registers.data\[578\] net1324 net855 top.CPU.registers.data\[610\]
+ net748 vssd1 vssd1 vccd1 vccd1 _05106_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout432_X net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout811_A net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout909_A net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08418_ _03719_ _03787_ _03786_ vssd1 vssd1 vccd1 vccd1 _04057_ sky130_fd_sc_hd__o21ai_1
X_09398_ net797 _05031_ _05032_ net751 vssd1 vssd1 vccd1 vccd1 _05037_ sky130_fd_sc_hd__o211a_1
X_08349_ _03958_ _03987_ vssd1 vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__or2_1
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08236__A2 net1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_129_Right_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_128_Left_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11360_ net3507 net287 net280 _06430_ vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__a22o_1
XFILLER_137_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout899_X net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07995__A1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10311_ _05826_ _05942_ net389 vssd1 vssd1 vccd1 vccd1 _05943_ sky130_fd_sc_hd__mux2_1
XANTENNA__11791__A2 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11291_ net570 _03183_ net486 vssd1 vssd1 vccd1 vccd1 _06704_ sky130_fd_sc_hd__and3_2
XFILLER_98_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13030_ net3038 _07440_ net895 vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__mux2_1
XFILLER_4_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10242_ top.CPU.fetch.current_ra\[27\] net1043 net882 top.CPU.handler.toreg\[27\]
+ vssd1 vssd1 vccd1 vccd1 _05877_ sky130_fd_sc_hd__a22o_1
XANTENNA__07528__A _03148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10200__C1 _05754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11543__A2 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1103 net1109 vssd1 vssd1 vccd1 vccd1 net1103 sky130_fd_sc_hd__clkbuf_4
X_10173_ net659 net573 net439 _05808_ vssd1 vssd1 vccd1 vccd1 _05810_ sky130_fd_sc_hd__and4_1
XFILLER_154_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1114 net1147 vssd1 vssd1 vccd1 vccd1 net1114 sky130_fd_sc_hd__clkbuf_2
Xfanout1125 net1127 vssd1 vssd1 vccd1 vccd1 net1125 sky130_fd_sc_hd__clkbuf_4
Xfanout1136 net1146 vssd1 vssd1 vccd1 vccd1 net1136 sky130_fd_sc_hd__buf_2
Xfanout1147 net1277 vssd1 vssd1 vccd1 vccd1 net1147 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_128_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input38_A nrst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14981_ clknet_leaf_96_clk _01226_ net1247 vssd1 vssd1 vccd1 vccd1 top.SPI.paroutput\[20\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1158 net1170 vssd1 vssd1 vccd1 vccd1 net1158 sky130_fd_sc_hd__clkbuf_4
Xfanout160 _06760_ vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10889__A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_137_Left_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout171 _06857_ vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__buf_4
Xfanout1169 net1170 vssd1 vssd1 vccd1 vccd1 net1169 sky130_fd_sc_hd__clkbuf_4
Xfanout182 _06777_ vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__clkbuf_8
Xfanout193 net195 vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10503__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11846__A3 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14185__355 clknet_leaf_157_clk vssd1 vssd1 vccd1 vccd1 net1824 sky130_fd_sc_hd__inv_2
X_12814_ _07251_ _07257_ _07264_ _07266_ vssd1 vssd1 vccd1 vccd1 _07267_ sky130_fd_sc_hd__nor4_1
XFILLER_16_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15602_ net1936 _01812_ net1102 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[402\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11059__A1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13794_ net23 net1050 net885 net3270 vssd1 vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__o22a_1
XANTENNA__11216__C net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12745_ top.CPU.alu.program_counter\[11\] _07202_ vssd1 vssd1 vccd1 vccd1 _07204_
+ sky130_fd_sc_hd__or2_1
X_15533_ net1867 _01743_ net1057 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[333\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09672__A1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14226__396 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 net1865 sky130_fd_sc_hd__inv_2
X_15464_ net1798 _01674_ net1087 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[264\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12008__B1 net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07710__B _03331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12676_ top.CPU.alu.program_counter\[2\] top.CPU.alu.program_counter\[3\] top.CPU.alu.program_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _07142_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_13_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08094__A net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08880__C1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_146_Left_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11232__B net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11627_ net130 net3322 net212 vssd1 vssd1 vccd1 vccd1 _01922_ sky130_fd_sc_hd__mux2_1
X_15395_ net1729 _01605_ net1207 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[195\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09424__A1 net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08381__X _04020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11558_ _06731_ _05990_ net440 net546 vssd1 vssd1 vccd1 vccd1 _06741_ sky130_fd_sc_hd__and4b_1
XANTENNA__08632__C1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11231__B2 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11782__A2 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold608 top.CPU.registers.data\[624\] vssd1 vssd1 vccd1 vccd1 net3165 sky130_fd_sc_hd__dlygate4sd3_1
X_10509_ net399 _05939_ _06132_ net412 vssd1 vssd1 vccd1 vccd1 _06133_ sky130_fd_sc_hd__o211a_1
XFILLER_171_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold619 top.CPU.registers.data\[510\] vssd1 vssd1 vccd1 vccd1 net3176 sky130_fd_sc_hd__dlygate4sd3_1
X_11489_ net487 net474 _06619_ net256 net3162 vssd1 vssd1 vccd1 vccd1 _02035_ sky130_fd_sc_hd__a32o_1
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09188__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16016_ net2350 _02226_ net1155 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[816\]
+ sky130_fd_sc_hd__dfrtp_1
X_13228_ net3486 _02776_ _02797_ vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_90_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11534__A2 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13159_ _06891_ _02747_ _02748_ vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08968__S net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_155_Left_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1308 top.CPU.registers.data\[45\] vssd1 vssd1 vccd1 vccd1 net3865 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1319 top.CPU.registers.data\[782\] vssd1 vssd1 vccd1 vccd1 net3876 sky130_fd_sc_hd__dlygate4sd3_1
X_07720_ net959 _03347_ _03348_ net947 vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__a211o_1
X_14888__1058 clknet_leaf_126_clk vssd1 vssd1 vccd1 vccd1 net2527 sky130_fd_sc_hd__inv_2
XANTENNA__08699__C1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11837__A3 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08163__A1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09360__B1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07651_ top.CPU.control_unit.instruction\[12\] _03245_ _03258_ _03260_ _03256_ vssd1
+ vssd1 vccd1 vccd1 _03290_ sky130_fd_sc_hd__a221oi_2
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11126__C net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07582_ top.CPU.registers.data\[1023\] net1334 net865 top.CPU.registers.data\[991\]
+ net802 vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__o221a_1
X_09321_ net708 _04959_ vssd1 vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_66_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10965__C net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07620__B net1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09252_ top.CPU.alu.program_counter\[5\] _04889_ net1033 vssd1 vssd1 vccd1 vccd1
+ _04891_ sky130_fd_sc_hd__mux2_2
XFILLER_33_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08871__C1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08203_ top.CPU.registers.data\[919\] net1295 net1014 top.CPU.registers.data\[951\]
+ net911 vssd1 vssd1 vccd1 vccd1 _03842_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_32_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09183_ net742 _04814_ _04815_ net767 vssd1 vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__o211a_1
XANTENNA__12953__S net1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10039__A top.CPU.alu.immediate\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12014__A3 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout225_A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10025__A2 _03292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08134_ top.CPU.registers.data\[597\] net1300 net1021 top.CPU.registers.data\[629\]
+ net941 vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__a221o_1
XANTENNA__09966__A2 _03407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08623__C1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10981__B net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11773__A2 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13908__78 clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 net1547 sky130_fd_sc_hd__inv_2
XFILLER_88_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08065_ top.CPU.registers.data\[916\] net1289 net1009 top.CPU.registers.data\[948\]
+ net906 vssd1 vssd1 vccd1 vccd1 _03704_ sky130_fd_sc_hd__a221o_1
XANTENNA__09179__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08926__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1301_A _03113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08878__S net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08967_ net783 _04604_ _04605_ net713 vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__o211a_1
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout761_A net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12701__B top.CPU.alu.program_counter\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout859_A net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07918_ net944 _03555_ _03556_ net958 vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__o211a_1
XANTENNA__11289__B2 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08898_ top.CPU.registers.data\[554\] top.CPU.registers.data\[522\] net809 vssd1
+ vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__mux2_1
XANTENNA__10502__A net1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14169__339 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 net1808 sky130_fd_sc_hd__inv_2
XFILLER_72_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07849_ top.CPU.registers.data\[573\] top.CPU.registers.data\[541\] net980 vssd1
+ vssd1 vccd1 vccd1 _03488_ sky130_fd_sc_hd__mux2_1
XANTENNA__10221__B net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1291_X net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout647_X net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1389_X net1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12238__B1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10860_ net525 _06466_ vssd1 vssd1 vccd1 vccd1 _06467_ sky130_fd_sc_hd__nor2_4
XFILLER_71_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09519_ net384 vssd1 vssd1 vccd1 vccd1 _05158_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_140_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10791_ _05057_ _05058_ vssd1 vssd1 vccd1 vccd1 _06402_ sky130_fd_sc_hd__nand2_1
XANTENNA__08457__A2 net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout814_X net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13024__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12530_ _07030_ _07038_ vssd1 vssd1 vccd1 vccd1 _07039_ sky130_fd_sc_hd__nor2_1
XANTENNA__10264__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07530__B net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08118__S net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12461_ _05466_ _05498_ vssd1 vssd1 vccd1 vccd1 _06970_ sky130_fd_sc_hd__and2_1
XANTENNA__08209__A2 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09406__A1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11412_ _06545_ net283 net269 net3448 vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__a22o_1
XANTENNA__11213__A1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15180_ net1517 _01390_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r1_prev\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_12392_ _06928_ _06929_ vssd1 vssd1 vccd1 vccd1 _06930_ sky130_fd_sc_hd__nor2_1
XANTENNA__08614__C1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10891__B net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07968__A1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12961__A1 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14570__740 clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 net2209 sky130_fd_sc_hd__inv_2
XANTENNA__11764__A2 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11343_ net3757 net287 net280 _06086_ vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__a22o_1
XANTENNA__08090__B1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11274_ net3081 net293 _06694_ net311 vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__a22o_1
X_13013_ top.SPI.parameters\[8\] top.SPI.paroutput\[0\] net1357 vssd1 vssd1 vccd1
+ vccd1 _07432_ sky130_fd_sc_hd__mux2_1
XANTENNA__08917__B1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11516__A2 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10225_ net390 _05859_ vssd1 vssd1 vccd1 vccd1 _05860_ sky130_fd_sc_hd__and2_1
X_14611__781 clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 net2250 sky130_fd_sc_hd__inv_2
XFILLER_121_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09590__B1 net1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13922__92 clknet_leaf_140_clk vssd1 vssd1 vccd1 vccd1 net1561 sky130_fd_sc_hd__inv_2
X_10156_ net411 _05757_ vssd1 vssd1 vccd1 vccd1 _05793_ sky130_fd_sc_hd__and2_2
Xhold5 top.CPU.registers.data_out_r1_prev\[21\] vssd1 vssd1 vccd1 vccd1 net2562 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11508__A net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12477__B1 _03955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10087_ _05723_ _05724_ net383 vssd1 vssd1 vccd1 vccd1 _05725_ sky130_fd_sc_hd__mux2_1
X_14964_ clknet_leaf_98_clk net2684 net1258 vssd1 vssd1 vccd1 vccd1 top.SPI.paroutput\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08145__A1 _03756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09342__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09893__A1 _04634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10131__B net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08696__A2 net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload3_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12229__B1 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08817__A net1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16456__D net1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13777_ net5 net1049 net884 net3925 vssd1 vssd1 vccd1 vccd1 _02658_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_48_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10989_ net513 net439 net143 net543 vssd1 vssd1 vccd1 vccd1 _06548_ sky130_fd_sc_hd__and4_1
X_15516_ net1850 _01726_ net1235 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[316\]
+ sky130_fd_sc_hd__dfrtp_1
X_12728_ top.CPU.alu.program_counter\[9\] _07173_ vssd1 vssd1 vccd1 vccd1 _07189_
+ sky130_fd_sc_hd__xor2_1
XFILLER_30_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08853__C1 net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16496_ clknet_leaf_41_clk _02658_ net1115 vssd1 vssd1 vccd1 vccd1 top.mmio.mem_data_i\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_148_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12659_ _03106_ _05232_ _07125_ _07124_ vssd1 vssd1 vccd1 vccd1 _07127_ sky130_fd_sc_hd__o31ai_2
X_15447_ net1781 _01657_ net1182 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[247\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_157_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11204__A1 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08552__A _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15378_ net1712 _01588_ net1100 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[178\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11755__A2 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10293__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold405 top.CPU.registers.data\[822\] vssd1 vssd1 vccd1 vccd1 net2962 sky130_fd_sc_hd__dlygate4sd3_1
Xhold416 top.I2C.output_state\[12\] vssd1 vssd1 vccd1 vccd1 net2973 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold427 top.CPU.registers.data\[6\] vssd1 vssd1 vccd1 vccd1 net2984 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12489__A1_N net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold438 top.CPU.registers.data\[570\] vssd1 vssd1 vccd1 vccd1 net2995 sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 top.CPU.registers.data\[985\] vssd1 vssd1 vccd1 vccd1 net3006 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10306__B _05616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09256__S0 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11507__A2 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09870_ _05506_ _05508_ _03581_ vssd1 vssd1 vccd1 vccd1 _05509_ sky130_fd_sc_hd__a21o_1
Xfanout907 net908 vssd1 vssd1 vccd1 vccd1 net907 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09030__C1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout918 net925 vssd1 vssd1 vccd1 vccd1 net918 sky130_fd_sc_hd__clkbuf_4
XFILLER_140_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout929 net949 vssd1 vssd1 vccd1 vccd1 net929 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09383__A _05021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08821_ _03099_ _04459_ net685 vssd1 vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__mux2_1
XFILLER_98_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wire448_X net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1105 top.I2C.I2C_state\[10\] vssd1 vssd1 vccd1 vccd1 net3662 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15127__RESET_B net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1116 top.CPU.registers.data\[250\] vssd1 vssd1 vccd1 vccd1 net3673 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1127 top.CPU.registers.data\[461\] vssd1 vssd1 vccd1 vccd1 net3684 sky130_fd_sc_hd__dlygate4sd3_1
X_08752_ net689 _04390_ _04365_ vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__o21ai_2
Xhold1138 top.CPU.registers.data\[37\] vssd1 vssd1 vccd1 vccd1 net3695 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12468__B1 _03887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08136__A1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1149 top.CPU.registers.data\[849\] vssd1 vssd1 vccd1 vccd1 net3706 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09333__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07703_ top.CPU.control_unit.instruction\[24\] net685 vssd1 vssd1 vccd1 vccd1 _03342_
+ sky130_fd_sc_hd__and2_4
X_08683_ _03116_ _04317_ _04320_ _04321_ net616 vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_105_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout175_A _06825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07634_ _03162_ net1037 vssd1 vssd1 vccd1 vccd1 _03273_ sky130_fd_sc_hd__nand2_1
XANTENNA__07902__Y _03541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_85_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07565_ net1047 _03163_ net1038 net1321 vssd1 vssd1 vccd1 vccd1 _03204_ sky130_fd_sc_hd__a31o_2
XANTENNA_fanout342_A net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11153__A net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09304_ net680 _04937_ _04938_ _04942_ net612 vssd1 vssd1 vccd1 vccd1 _04943_ sky130_fd_sc_hd__a311o_1
XANTENNA__10246__A2 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07496_ top.SPI.state\[4\] vssd1 vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__inv_2
XANTENNA__08844__C1 _03342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09235_ _04872_ _04873_ net635 vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__a21o_1
XANTENNA__11994__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10992__A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1251_A net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout607_A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout228_X net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14554__724 clknet_leaf_163_clk vssd1 vssd1 vccd1 vccd1 net2193 sky130_fd_sc_hd__inv_2
XANTENNA_fanout1349_A top.CPU.handler.state\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09166_ _04801_ _04804_ net742 vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__o21a_1
XFILLER_5_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08117_ net1368 net1045 net899 vssd1 vssd1 vccd1 vccd1 _03756_ sky130_fd_sc_hd__o21a_2
XANTENNA__11746__A2 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09097_ top.CPU.registers.data\[39\] top.CPU.registers.data\[7\] net832 vssd1 vssd1
+ vccd1 vccd1 _04736_ sky130_fd_sc_hd__mux2_1
XANTENNA__08611__A2 net1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08048_ top.CPU.registers.data\[20\] net979 _03686_ vssd1 vssd1 vccd1 vccd1 _03687_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__15068__Q top.I2C.output_state\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold950 top.CPU.registers.data\[738\] vssd1 vssd1 vccd1 vccd1 net3507 sky130_fd_sc_hd__dlygate4sd3_1
Xhold961 top.CPU.registers.data\[651\] vssd1 vssd1 vccd1 vccd1 net3518 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout976_A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold972 top.CPU.registers.data\[960\] vssd1 vssd1 vccd1 vccd1 net3529 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_164_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold983 top.CPU.registers.data\[350\] vssd1 vssd1 vccd1 vccd1 net3540 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12712__A top.CPU.alu.program_counter\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold994 top.CPU.registers.data\[165\] vssd1 vssd1 vccd1 vccd1 net3551 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1304_X net1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08375__A1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10010_ _05647_ _05648_ net385 vssd1 vssd1 vccd1 vccd1 _05649_ sky130_fd_sc_hd__mux2_1
XANTENNA__12171__A2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09999_ _04363_ _04430_ net378 vssd1 vssd1 vccd1 vccd1 _05638_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout764_X net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07583__C1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10232__A net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09324__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11961_ top.CPU.registers.data\[199\] net231 vssd1 vssd1 vccd1 vccd1 _06776_ sky130_fd_sc_hd__and2_1
XANTENNA__12858__S net1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout931_X net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11131__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08222__S1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13700_ top.SPI.timem\[2\] _03052_ net3473 vssd1 vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__a21oi_1
X_10912_ net3681 net221 _06501_ net461 vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__a22o_1
XFILLER_45_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11682__A1 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11892_ _06373_ net3360 net188 vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__mux2_1
XFILLER_71_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13631_ net3372 _07135_ net664 vssd1 vssd1 vccd1 vccd1 _02565_ sky130_fd_sc_hd__mux2_1
X_10843_ _03323_ _05609_ _06450_ _03322_ vssd1 vssd1 vccd1 vccd1 _06451_ sky130_fd_sc_hd__a22oi_1
XFILLER_44_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09627__A1 _05265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16350_ clknet_leaf_68_clk _02559_ net1167 vssd1 vssd1 vccd1 vccd1 top.CPU.addressnew\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13562_ top.CPU.alu.program_counter\[5\] net1348 net583 vssd1 vssd1 vccd1 vccd1 _03004_
+ sky130_fd_sc_hd__o21a_1
X_10774_ _03315_ _04990_ _05680_ _04988_ _06385_ vssd1 vssd1 vccd1 vccd1 _06386_ sky130_fd_sc_hd__a221o_1
XANTENNA__08835__C1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12513_ _04499_ _04531_ vssd1 vssd1 vccd1 vccd1 _07022_ sky130_fd_sc_hd__nand2_1
X_15301_ net1635 _01511_ net1087 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[101\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11985__A2 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16281_ clknet_leaf_58_clk _02491_ net1144 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.toreg\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13493_ top.CPU.data_out\[7\] _04792_ net587 vssd1 vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_160_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_160_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_173_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12444_ _06894_ _06958_ vssd1 vssd1 vccd1 vccd1 _00050_ sky130_fd_sc_hd__nor2_1
X_15232_ net1566 _01442_ net1175 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[32\]
+ sky130_fd_sc_hd__dfrtp_1
X_14297__467 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 net1936 sky130_fd_sc_hd__inv_2
X_14887__1057 clknet_leaf_185_clk vssd1 vssd1 vccd1 vccd1 net2526 sky130_fd_sc_hd__inv_2
XANTENNA__11737__A2 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15163_ clknet_leaf_91_clk _01373_ vssd1 vssd1 vccd1 vccd1 top.SPI.percount\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_12375_ top.I2C.I2C_state\[23\] top.I2C.I2C_state\[20\] top.I2C.I2C_state\[25\] vssd1
+ vssd1 vccd1 vccd1 _06915_ sky130_fd_sc_hd__or3_1
XFILLER_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09260__C1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10407__A net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08602__A2 net1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11326_ net475 _06519_ net428 vssd1 vssd1 vccd1 vccd1 _06711_ sky130_fd_sc_hd__and3_1
XFILLER_119_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15094_ net1476 _01307_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r2_prev\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07810__B1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13899__69 clknet_leaf_135_clk vssd1 vssd1 vccd1 vccd1 net1538 sky130_fd_sc_hd__inv_2
X_11257_ net2967 net293 _06684_ net483 vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__a22o_1
X_10208_ _03580_ _05602_ _05603_ vssd1 vssd1 vccd1 vccd1 _05844_ sky130_fd_sc_hd__nand3_1
XANTENNA__09563__B1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09407__S net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11188_ net139 net430 vssd1 vssd1 vccd1 vccd1 _06653_ sky130_fd_sc_hd__and2_1
XANTENNA__11370__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10139_ _05621_ _05630_ net305 vssd1 vssd1 vccd1 vccd1 _05776_ sky130_fd_sc_hd__mux2_1
XFILLER_39_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15996_ net2330 _02206_ net1235 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[796\]
+ sky130_fd_sc_hd__dfrtp_1
X_14947_ clknet_leaf_65_clk _01193_ net1163 vssd1 vssd1 vccd1 vccd1 top.CPU.alu.program_counter\[30\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_36_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07877__B1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16617_ net1347 vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__clkbuf_1
X_13829_ net2899 net335 net328 top.CPU.data_out\[31\] vssd1 vssd1 vccd1 vccd1 _02709_
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14241__411 clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 net1880 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_63_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16548_ clknet_leaf_63_clk _02710_ net1161 vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__dfrtp_2
X_14538__708 clknet_leaf_145_clk vssd1 vssd1 vccd1 vccd1 net2177 sky130_fd_sc_hd__inv_2
XANTENNA__11976__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16479_ clknet_leaf_89_clk _02641_ net1273 vssd1 vssd1 vccd1 vccd1 top.SPI.timem\[22\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_151_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_151_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_15_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09020_ top.CPU.registers.data_out_r2_prev\[9\] net688 _04657_ vssd1 vssd1 vccd1
+ vccd1 _04659_ sky130_fd_sc_hd__o21a_1
XFILLER_163_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08282__A _03889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16272__Q top.CPU.handler.toreg\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold202 top.CPU.registers.data\[255\] vssd1 vssd1 vccd1 vccd1 net2759 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold213 net89 vssd1 vssd1 vccd1 vccd1 net2770 sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 _00035_ vssd1 vssd1 vccd1 vccd1 net2781 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07801__A0 _03439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold235 top.SPI.parameters\[10\] vssd1 vssd1 vccd1 vccd1 net2792 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold246 top.CPU.registers.data\[175\] vssd1 vssd1 vccd1 vccd1 net2803 sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 top.CPU.registers.data\[826\] vssd1 vssd1 vccd1 vccd1 net2814 sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 top.CPU.registers.data\[172\] vssd1 vssd1 vccd1 vccd1 net2825 sky130_fd_sc_hd__dlygate4sd3_1
Xhold279 net74 vssd1 vssd1 vccd1 vccd1 net2836 sky130_fd_sc_hd__dlygate4sd3_1
X_09922_ _04862_ _05559_ _05560_ vssd1 vssd1 vccd1 vccd1 _05561_ sky130_fd_sc_hd__a21o_1
Xfanout704 net706 vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__clkbuf_4
Xfanout715 net717 vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__clkbuf_4
Xfanout726 net728 vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12153__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout737 net739 vssd1 vssd1 vccd1 vccd1 net737 sky130_fd_sc_hd__clkbuf_4
X_09853_ top.CPU.registers.data\[282\] net1000 _05491_ vssd1 vssd1 vccd1 vccd1 _05492_
+ sky130_fd_sc_hd__a21o_1
Xfanout748 net749 vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11361__B1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout759 net760 vssd1 vssd1 vccd1 vccd1 net759 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_142_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08804_ _04441_ _04442_ net674 vssd1 vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__o21a_1
XFILLER_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09784_ net942 _05402_ _05403_ net956 vssd1 vssd1 vccd1 vccd1 _05423_ sky130_fd_sc_hd__o211a_1
XFILLER_86_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09306__B1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07580__A2 net1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08735_ top.CPU.registers.data\[77\] net1371 net967 top.CPU.registers.data\[109\]
+ net910 vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__o221a_1
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11113__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10987__A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09857__A1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout557_A _07418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout178_X net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1299_A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08666_ top.CPU.registers.data\[78\] net1375 net981 top.CPU.registers.data\[110\]
+ net908 vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__o221a_1
XFILLER_82_952 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11664__A1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07617_ net1408 net1278 _03154_ vssd1 vssd1 vccd1 vccd1 _03256_ sky130_fd_sc_hd__or3_1
XFILLER_121_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09609__A1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08597_ top.CPU.registers.data\[79\] net1375 net974 top.CPU.registers.data\[111\]
+ net903 vssd1 vssd1 vccd1 vccd1 _04236_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout724_A net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout345_X net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10219__A2 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07548_ _03186_ vssd1 vssd1 vccd1 vccd1 _03187_ sky130_fd_sc_hd__inv_2
XANTENNA__11020__C_N net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11967__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07479_ top.I2C.output_state\[0\] vssd1 vssd1 vccd1 vccd1 _03119_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_142_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_142_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_167_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09218_ _04855_ _04856_ net452 vssd1 vssd1 vccd1 vccd1 _04857_ sky130_fd_sc_hd__mux2_1
X_10490_ net414 _06114_ net224 vssd1 vssd1 vccd1 vccd1 _06115_ sky130_fd_sc_hd__o21bai_1
XFILLER_155_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14025__195 clknet_leaf_156_clk vssd1 vssd1 vccd1 vccd1 net1664 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_20_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_101_Left_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11719__A2 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09149_ top.CPU.registers.data\[839\] net1304 net1024 top.CPU.registers.data\[871\]
+ net943 vssd1 vssd1 vccd1 vccd1 _04788_ sky130_fd_sc_hd__a221o_1
XANTENNA__10227__A _05667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12160_ _06311_ net360 net354 net172 top.CPU.registers.data\[72\] vssd1 vssd1 vccd1
+ vccd1 _06848_ sky130_fd_sc_hd__a32o_1
XFILLER_123_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout881_X net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11111_ net488 net464 _06613_ net303 net3094 vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__a32o_1
XANTENNA__11757__S net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout979_X net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10661__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12091_ _06627_ net244 net176 top.CPU.registers.data\[107\] vssd1 vssd1 vccd1 vccd1
+ _06814_ sky130_fd_sc_hd__a22o_1
XANTENNA__12442__A net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold780 top.CPU.registers.data\[661\] vssd1 vssd1 vccd1 vccd1 net3337 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08348__A1 _03986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold791 top.CPU.registers.data\[480\] vssd1 vssd1 vccd1 vccd1 net3348 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07536__A net1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11042_ net531 _05694_ _06479_ vssd1 vssd1 vccd1 vccd1 _06580_ sky130_fd_sc_hd__and3_1
XFILLER_49_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08899__A2 net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11352__B1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15850_ net2184 _02060_ net1084 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[650\]
+ sky130_fd_sc_hd__dfrtp_1
X_14682__852 clknet_leaf_165_clk vssd1 vssd1 vccd1 vccd1 net2321 sky130_fd_sc_hd__inv_2
XFILLER_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_110_Left_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07571__A2 net1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input20_A DAT_I[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15781_ net2115 _01991_ net1087 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[581\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09848__A1 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12993_ _03127_ top.SPI.state\[1\] _07421_ vssd1 vssd1 vccd1 vccd1 _07422_ sky130_fd_sc_hd__nor3_1
XANTENNA__10897__A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11944_ top.CPU.registers.data\[214\] net232 vssd1 vssd1 vccd1 vccd1 _06774_ sky130_fd_sc_hd__and2_1
X_14723__893 clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 net2362 sky130_fd_sc_hd__inv_2
XANTENNA__08367__A net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08520__A1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11875_ _06708_ net239 net190 net3245 vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_28_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16402_ clknet_leaf_62_clk _00025_ net1163 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.state\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13614_ net2827 _03035_ net580 vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__mux2_1
X_10826_ _05193_ net504 _05678_ vssd1 vssd1 vccd1 vccd1 _06435_ sky130_fd_sc_hd__o21a_1
XANTENNA__08808__C1 net1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11958__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16333_ clknet_leaf_68_clk _02542_ net1167 vssd1 vssd1 vccd1 vccd1 top.CPU.addressnew\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13545_ top.CPU.data_out\[31\] _03370_ net589 vssd1 vssd1 vccd1 vccd1 _02529_ sky130_fd_sc_hd__mux2_1
X_10757_ _05543_ _05556_ net511 vssd1 vssd1 vccd1 vccd1 _06370_ sky130_fd_sc_hd__o21ai_1
XFILLER_13_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_133_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_133_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_158_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13476_ net3906 _02959_ net124 vssd1 vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__mux2_1
X_16264_ clknet_leaf_44_clk _02474_ net1124 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.toreg\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_173_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10688_ _04731_ _05670_ _06302_ _06303_ vssd1 vssd1 vccd1 vccd1 _06304_ sky130_fd_sc_hd__a211o_1
XFILLER_145_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12427_ _03129_ net3206 _06950_ vssd1 vssd1 vccd1 vccd1 _00067_ sky130_fd_sc_hd__a21oi_1
X_15215_ net1549 _01425_ net1099 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11240__B net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09233__C1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16195_ net2529 _02405_ net1206 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[995\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10918__B1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13580__A1 top.CPU.alu.program_counter\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12358_ top.I2C.I2C_state\[15\] top.I2C.I2C_state\[14\] top.I2C.I2C_state\[17\] top.I2C.I2C_state\[18\]
+ vssd1 vssd1 vccd1 vccd1 _06901_ sky130_fd_sc_hd__or4_1
X_15146_ clknet_leaf_48_clk _01356_ net1130 vssd1 vssd1 vccd1 vccd1 top.I2C.data_out\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_126_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11667__S net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07795__C1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11309_ net3449 net290 net358 net146 vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__a22o_1
X_15077_ clknet_leaf_49_clk _00055_ net1129 vssd1 vssd1 vccd1 vccd1 top.I2C.output_state\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_113_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12289_ net2626 _04019_ net1106 vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__mux2_1
XANTENNA__08339__A1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12135__A2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11343__B1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13096__A0 top.CPU.data_out\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15979_ net2313 _02189_ net1064 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[779\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11118__D net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08520_ net880 _04155_ _04157_ vssd1 vssd1 vccd1 vccd1 _04159_ sky130_fd_sc_hd__o21a_1
XANTENNA__10600__A net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08511__A1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08451_ top.CPU.registers.data_out_r1_prev\[17\] net875 _04075_ _04089_ vssd1 vssd1
+ vccd1 vccd1 _04090_ sky130_fd_sc_hd__o211ai_4
XANTENNA__13399__B2 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08382_ net880 _04019_ _03990_ vssd1 vssd1 vccd1 vccd1 _04021_ sky130_fd_sc_hd__o21ai_2
XFILLER_91_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11949__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14009__179 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 net1648 sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_124_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_124_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10973__C net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11431__A net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout138_A _05692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08216__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09003_ top.CPU.registers.data\[809\] top.CPU.registers.data\[777\] net965 vssd1
+ vssd1 vccd1 vccd1 _04642_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_152_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08027__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08122__S0 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13571__A1 _06288_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11177__A3 _06648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1214_A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout501 _05696_ vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__buf_4
XANTENNA__13323__A1 _02861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14666__836 clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 net2305 sky130_fd_sc_hd__inv_2
XANTENNA__09047__S net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12126__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout512 _05520_ vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__clkbuf_2
X_09905_ net401 _05055_ vssd1 vssd1 vccd1 vccd1 _05544_ sky130_fd_sc_hd__nor2_1
Xfanout523 _03197_ vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__buf_2
Xfanout534 net537 vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__buf_4
XANTENNA_fanout295_X net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout545 net546 vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__buf_4
XANTENNA__11334__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout674_A net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout556 _02847_ vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10688__A2 _05670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09836_ net960 _05469_ _05471_ _05474_ vssd1 vssd1 vccd1 vccd1 _05475_ sky130_fd_sc_hd__a31o_1
Xfanout567 net569 vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__buf_4
XFILLER_100_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout578 net579 vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__clkbuf_4
XFILLER_112_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1002_X net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout589 net590 vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__buf_2
X_14410__580 clknet_leaf_152_clk vssd1 vssd1 vccd1 vccd1 net2049 sky130_fd_sc_hd__inv_2
XFILLER_86_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10213__C net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14707__877 clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 net2346 sky130_fd_sc_hd__inv_2
XANTENNA_fanout841_A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09767_ top.CPU.registers.data\[859\] net1298 net1019 top.CPU.registers.data\[891\]
+ net942 vssd1 vssd1 vccd1 vccd1 _05406_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout462_X net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout939_A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14886__1056 clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 net2525 sky130_fd_sc_hd__inv_2
XFILLER_73_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08718_ net784 _04347_ _04348_ net738 vssd1 vssd1 vccd1 vccd1 _04357_ sky130_fd_sc_hd__o211a_1
XFILLER_132_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09698_ top.CPU.registers.data\[857\] net1306 net1029 top.CPU.registers.data\[889\]
+ net946 vssd1 vssd1 vccd1 vccd1 _05337_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_159_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08649_ net792 _04287_ _04286_ net744 vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__o211a_1
XFILLER_70_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout727_X net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11660_ _06449_ net208 net427 net3294 vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__a22o_1
XFILLER_25_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10611_ net660 _06230_ vssd1 vssd1 vccd1 vccd1 _06231_ sky130_fd_sc_hd__and2_2
XANTENNA__08266__B1 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12062__A1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11591_ net653 net363 vssd1 vssd1 vccd1 vccd1 _06750_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_115_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_115_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_137_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09463__C1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13330_ net888 _02866_ vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__and2_1
X_10542_ net404 _05977_ vssd1 vssd1 vccd1 vccd1 _06165_ sky130_fd_sc_hd__or2_1
XFILLER_128_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08126__S net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13261_ net3980 _02814_ _02815_ net1053 vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__a22o_1
XANTENNA__11060__B net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08018__B1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10473_ _05741_ _06098_ vssd1 vssd1 vccd1 vccd1 _06099_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_133_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13011__B1 _07431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15000_ clknet_leaf_98_clk _01245_ net1258 vssd1 vssd1 vccd1 vccd1 top.SPI.parameters\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_124_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12212_ _06213_ net542 _06796_ net168 top.CPU.registers.data\[45\] vssd1 vssd1 vccd1
+ vccd1 _06873_ sky130_fd_sc_hd__a32o_1
XFILLER_136_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13562__A1 top.CPU.alu.program_counter\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13192_ top.I2C.which_data_address\[1\] top.I2C.which_data_address\[2\] vssd1 vssd1
+ vccd1 vccd1 _02772_ sky130_fd_sc_hd__and2b_1
XFILLER_108_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08650__A net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12143_ net3940 net174 _06839_ _06653_ vssd1 vssd1 vccd1 vccd1 _01491_ sky130_fd_sc_hd__a22o_1
XFILLER_151_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09518__A0 _05154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13869__39 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 net1508 sky130_fd_sc_hd__inv_2
XANTENNA__12117__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12074_ net473 _06616_ _06805_ net177 net3861 vssd1 vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__a32o_1
XFILLER_132_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11325__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11025_ _06447_ net541 vssd1 vssd1 vccd1 vccd1 _06570_ sky130_fd_sc_hd__or2_1
X_15902_ net2236 _02112_ net1239 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[702\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13078__A0 top.CPU.data_out\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15833_ net2167 _02043_ net1223 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[633\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_64_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15764_ net2098 _01974_ net1082 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[564\]
+ sky130_fd_sc_hd__dfrtp_1
X_12976_ top.I2C.bit_timer_counter\[4\] _07409_ vssd1 vssd1 vccd1 vccd1 _07410_ sky130_fd_sc_hd__or2_1
XFILLER_73_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11927_ net3464 net184 net342 _06375_ vssd1 vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__a22o_1
XANTENNA__13153__D top.I2C.output_state\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10300__A1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15695_ net2029 _01905_ net1097 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[495\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11858_ _06694_ net197 net152 net2895 vssd1 vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__a22o_1
XFILLER_32_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10809_ _05672_ _06091_ _06098_ _05665_ _06141_ vssd1 vssd1 vccd1 vccd1 _06419_ sky130_fd_sc_hd__a221oi_2
Xclkbuf_leaf_106_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_106_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_14_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11789_ net467 _06635_ net239 net162 net3072 vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__a32o_1
XFILLER_41_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11251__A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08352__S0 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16316_ clknet_leaf_83_clk _02525_ net1262 vssd1 vssd1 vccd1 vccd1 top.CPU.data_out\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13528_ top.CPU.data_out\[22\] net589 net339 _02984_ vssd1 vssd1 vccd1 vccd1 _02520_
+ sky130_fd_sc_hd__o22a_1
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16247_ clknet_leaf_43_clk _02457_ net1123 vssd1 vssd1 vccd1 vccd1 top.CPU.control_unit.instruction\[23\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_9_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_191_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13459_ net1396 net873 _02903_ net418 vssd1 vssd1 vccd1 vccd1 _02951_ sky130_fd_sc_hd__a31o_1
XFILLER_63_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09206__C1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 STB_O sky130_fd_sc_hd__buf_2
X_14353__523 clknet_leaf_190_clk vssd1 vssd1 vccd1 vccd1 net1992 sky130_fd_sc_hd__inv_2
Xoutput115 net115 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__buf_2
XANTENNA__10367__A1 _03889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_71_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16178_ net2512 _02388_ net1101 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[978\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_58_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11564__B1 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15129_ clknet_leaf_57_clk _01339_ net1145 vssd1 vssd1 vccd1 vccd1 top.I2C.within_byte_counter_writing\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_126_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13305__A1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12108__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09509__B1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07783__A2 net1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07951_ top.CPU.registers.data\[472\] net1321 net852 top.CPU.registers.data\[504\]
+ net771 vssd1 vssd1 vccd1 vccd1 _03590_ sky130_fd_sc_hd__a221o_1
XANTENNA__11316__B1 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_86_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07882_ net700 _03519_ _03520_ vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_71_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08193__C1 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13069__A0 top.CPU.data_out\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09621_ net788 _05253_ _05254_ net691 vssd1 vssd1 vccd1 vccd1 _05260_ sky130_fd_sc_hd__a31o_1
X_13883__53 clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 net1522 sky130_fd_sc_hd__inv_2
X_09552_ _05190_ vssd1 vssd1 vccd1 vccd1 _05191_ sky130_fd_sc_hd__inv_2
XANTENNA__10330__A _05697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09288__A2 net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08503_ top.CPU.registers.data\[752\] net1390 net821 top.CPU.registers.data\[720\]
+ net721 vssd1 vssd1 vccd1 vccd1 _04142_ sky130_fd_sc_hd__a221o_1
X_09483_ top.CPU.alu.program_counter\[2\] net1033 vssd1 vssd1 vccd1 vccd1 _05122_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__11095__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout255_A _06728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_144_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08434_ net796 _04067_ _04068_ net750 vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__o211a_1
XFILLER_169_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10984__B net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13360__B net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08365_ net769 _03992_ _03996_ _04003_ vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_154_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_24_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout422_A net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1164_A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11161__A net1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13961__131 clknet_leaf_158_clk vssd1 vssd1 vccd1 vccd1 net1600 sky130_fd_sc_hd__inv_2
X_08296_ net796 _03930_ _03931_ net749 vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_115_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_159_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12691__S net1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_2_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_2_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout210_X net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1331_A _03109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13544__A1 top.CPU.data_out\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09748__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_250 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_39_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14096__266 clknet_leaf_199_clk vssd1 vssd1 vccd1 vccd1 net1735 sky130_fd_sc_hd__inv_2
XANTENNA__08470__A net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09212__A2 net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout791_A net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12704__B _04793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10358__B2 top.CPU.handler.toreg\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11555__B1 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout889_A net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07774__A2 net1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1307 _03113_ vssd1 vssd1 vccd1 vccd1 net1307 sky130_fd_sc_hd__clkbuf_4
Xfanout320 net322 vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__buf_2
XFILLER_114_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout677_X net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11307__B1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1318 net1319 vssd1 vssd1 vccd1 vccd1 net1318 sky130_fd_sc_hd__buf_2
Xfanout331 net332 vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__buf_2
XFILLER_132_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1329 net1331 vssd1 vssd1 vccd1 vccd1 net1329 sky130_fd_sc_hd__clkbuf_4
Xfanout342 net343 vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__buf_4
Xfanout353 _06771_ vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__buf_2
Xfanout364 net365 vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__clkbuf_8
Xfanout375 net376 vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__buf_2
Xfanout386 net393 vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__clkbuf_4
XFILLER_19_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout397 net398 vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__buf_2
X_09819_ top.CPU.registers.data\[90\] net1337 net868 top.CPU.registers.data\[122\]
+ net757 vssd1 vssd1 vccd1 vccd1 _05458_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout844_X net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07931__C1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12830_ _07280_ _07281_ vssd1 vssd1 vccd1 vccd1 _07282_ sky130_fd_sc_hd__nor2_1
XANTENNA__07533__B net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11055__B net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12761_ _07203_ _07215_ _07217_ vssd1 vssd1 vccd1 vccd1 _07219_ sky130_fd_sc_hd__nand3_1
XANTENNA__11086__A2 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09684__C1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _06548_ net199 net420 net2960 vssd1 vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__a22o_1
X_12692_ top.CPU.alu.program_counter\[6\] _04856_ vssd1 vssd1 vccd1 vccd1 _07156_
+ sky130_fd_sc_hd__nand2_1
X_14794__964 clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 net2433 sky130_fd_sc_hd__inv_2
X_15480_ net1814 _01690_ net1150 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[280\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08239__B1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11643_ _06107_ net200 net425 net3278 vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__a22o_1
XFILLER_52_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11071__A _06311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11574_ net570 _06685_ vssd1 vssd1 vccd1 vccd1 _06745_ sky130_fd_sc_hd__nor2_1
X_14040__210 clknet_leaf_166_clk vssd1 vssd1 vccd1 vccd1 net1679 sky130_fd_sc_hd__inv_2
XFILLER_156_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10597__A1 _04430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput17 DAT_I[23] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
XFILLER_168_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput28 DAT_I[4] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
X_16101_ net2435 _02311_ net1062 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[901\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_155_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10525_ net602 _06147_ _06148_ vssd1 vssd1 vccd1 vccd1 _06149_ sky130_fd_sc_hd__a21o_1
X_13313_ top.I2C.data_out\[2\] net553 _02853_ vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__a21oi_1
X_14337__507 clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 net1976 sky130_fd_sc_hd__inv_2
XFILLER_155_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13244_ net3837 _02805_ _02806_ _02803_ vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__a22o_1
XANTENNA__09739__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16032_ net2366 _02242_ net1093 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[832\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10456_ top.CPU.fetch.current_ra\[19\] net1041 net881 top.CPU.handler.toreg\[19\]
+ vssd1 vssd1 vccd1 vccd1 _06083_ sky130_fd_sc_hd__a22oi_4
XANTENNA__09203__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10349__B2 _03823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11546__B1 _06734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13175_ top.I2C.within_byte_counter_writing\[0\] top.I2C.within_byte_counter_writing\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__or2_1
XFILLER_124_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10387_ _03756_ net506 vssd1 vssd1 vccd1 vccd1 _06016_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_36_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12126_ top.CPU.registers.data\[89\] net655 _06749_ vssd1 vssd1 vccd1 vccd1 _06831_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_36_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10134__B net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11849__A1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12057_ top.CPU.registers.data\[124\] net657 _03185_ vssd1 vssd1 vccd1 vccd1 _06797_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__10702__X _06317_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11008_ net3559 net216 _06559_ net312 vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__a22o_1
XANTENNA__12510__A2 _04324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07922__C1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08190__A2 net1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11246__A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15816_ net2150 _02026_ net1100 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[616\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10809__C1 _06141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15747_ net2081 _01957_ net1206 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[547\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12274__A1 _03241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12959_ _07393_ _07394_ _07395_ _07397_ net128 vssd1 vssd1 vccd1 vccd1 _07398_ sky130_fd_sc_hd__o311a_1
XANTENNA__13471__B1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15678_ net2012 _01888_ net1238 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[478\]
+ sky130_fd_sc_hd__dfrtp_1
X_13945__115 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 net1584 sky130_fd_sc_hd__inv_2
XFILLER_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09427__C1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08150_ _03786_ _03788_ vssd1 vssd1 vccd1 vccd1 _03789_ sky130_fd_sc_hd__nand2_2
XANTENNA__09442__A2 net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11785__B1 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08081_ _03719_ vssd1 vssd1 vccd1 vccd1 _03720_ sky130_fd_sc_hd__inv_2
XFILLER_119_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14885__1055 clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 net2524 sky130_fd_sc_hd__inv_2
XFILLER_134_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11537__B1 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16280__Q top.CPU.handler.toreg\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07618__B top.CPU.control_unit.instruction\[27\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_114_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08953__A1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07756__A2 net1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08983_ top.CPU.registers.data\[297\] top.CPU.registers.data\[265\] net805 vssd1
+ vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__mux2_1
XFILLER_130_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07905__Y _03544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07934_ net961 _03567_ _03569_ _03572_ vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__a31o_1
XFILLER_102_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_147_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08166__C1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10979__B net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07865_ top.CPU.registers.data\[477\] net1289 net1007 top.CPU.registers.data\[509\]
+ net905 vssd1 vssd1 vccd1 vccd1 _03504_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout372_A net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11156__A net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09604_ top.CPU.registers.data\[448\] net1313 net844 top.CPU.registers.data\[480\]
+ net766 vssd1 vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_108_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07796_ top.CPU.registers.data\[350\] net1303 net1025 top.CPU.registers.data\[382\]
+ net944 vssd1 vssd1 vccd1 vccd1 _03435_ sky130_fd_sc_hd__a221o_1
XFILLER_113_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481__651 clknet_leaf_187_clk vssd1 vssd1 vccd1 vccd1 net2120 sky130_fd_sc_hd__inv_2
XANTENNA__11068__A2 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14778__948 clknet_leaf_158_clk vssd1 vssd1 vccd1 vccd1 net2417 sky130_fd_sc_hd__inv_2
XANTENNA__12265__A1 _06354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09535_ _05166_ _05173_ net642 vssd1 vssd1 vccd1 vccd1 _05174_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout160_X net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1281_A net1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout637_A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout258_X net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10276__B1 _05367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1379_A net1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09466_ _05101_ _05104_ net637 vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__a21o_1
XFILLER_19_1038 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14522__692 clknet_leaf_158_clk vssd1 vssd1 vccd1 vccd1 net2161 sky130_fd_sc_hd__inv_2
XFILLER_40_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09681__A2 net1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08417_ _04055_ vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__inv_2
X_09397_ net797 _05025_ _05026_ net727 vssd1 vssd1 vccd1 vccd1 _05036_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout425_X net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14819__989 clknet_leaf_114_clk vssd1 vssd1 vccd1 vccd1 net2458 sky130_fd_sc_hd__inv_2
XANTENNA_fanout804_A _03205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08348_ _03984_ _03986_ net454 vssd1 vssd1 vccd1 vccd1 _03987_ sky130_fd_sc_hd__mux2_1
XANTENNA__09433__A2 net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11776__B1 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08279_ _03917_ vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__inv_2
XFILLER_20_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08641__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13832__2 clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 net1471 sky130_fd_sc_hd__inv_2
XANTENNA__12715__A top.CPU.alu.program_counter\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1334_X net1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10310_ _05885_ _05941_ net308 vssd1 vssd1 vccd1 vccd1 _05942_ sky130_fd_sc_hd__mux2_1
XFILLER_4_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11290_ net137 net2911 net291 vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__mux2_1
XFILLER_164_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11528__B1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout794_X net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10241_ _05853_ _05855_ _05875_ vssd1 vssd1 vccd1 vccd1 _05876_ sky130_fd_sc_hd__a21o_1
XANTENNA__07528__B net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07747__A2 net1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10172_ net659 _05808_ vssd1 vssd1 vccd1 vccd1 _05809_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout961_X net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1104 net1105 vssd1 vssd1 vccd1 vccd1 net1104 sky130_fd_sc_hd__clkbuf_4
XFILLER_105_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1115 net1118 vssd1 vssd1 vccd1 vccd1 net1115 sky130_fd_sc_hd__clkbuf_4
XFILLER_105_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1126 net1127 vssd1 vssd1 vccd1 vccd1 net1126 sky130_fd_sc_hd__buf_2
XFILLER_121_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14980_ clknet_leaf_93_clk _01225_ net1267 vssd1 vssd1 vccd1 vccd1 top.SPI.paroutput\[19\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1137 net1140 vssd1 vssd1 vccd1 vccd1 net1137 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_128_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout150 _06780_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__buf_6
Xfanout1148 net1151 vssd1 vssd1 vccd1 vccd1 net1148 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_128_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1159 net1170 vssd1 vssd1 vccd1 vccd1 net1159 sky130_fd_sc_hd__buf_2
Xfanout161 _06760_ vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10889__B _06010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout172 _06825_ vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__buf_4
XANTENNA__07544__A _03180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout183 _06777_ vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__clkbuf_4
Xfanout194 net195 vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__buf_6
XFILLER_47_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11700__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15601_ net1935 _01811_ net1189 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[401\]
+ sky130_fd_sc_hd__dfrtp_1
X_12813_ top.CPU.alu.program_counter\[17\] _04123_ vssd1 vssd1 vccd1 vccd1 _07266_
+ sky130_fd_sc_hd__and2_1
XANTENNA__12256__A1 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11059__A2 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13793_ net22 net1050 net885 net3755 vssd1 vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__o22a_1
XANTENNA__13453__B1 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09121__A1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15532_ net1866 _01742_ net1069 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[332\]
+ sky130_fd_sc_hd__dfrtp_1
X_12744_ top.CPU.alu.program_counter\[11\] _07202_ vssd1 vssd1 vccd1 vccd1 _07203_
+ sky130_fd_sc_hd__nand2_1
XFILLER_72_1007 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12008__A1 _06577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09409__C1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15463_ net1797 _01673_ net1201 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[263\]
+ sky130_fd_sc_hd__dfrtp_1
X_12675_ _07139_ _07140_ vssd1 vssd1 vccd1 vccd1 _07141_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_13_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10019__A0 _03613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11626_ _06519_ _06701_ net209 net215 net2930 vssd1 vssd1 vccd1 vccd1 _01923_ sky130_fd_sc_hd__a32o_1
X_15394_ net1728 _01604_ net1173 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[194\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11767__B1 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11231__A2 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08632__B1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11557_ _06670_ net258 net247 net2773 vssd1 vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__a22o_1
XFILLER_156_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10508_ net399 _05946_ vssd1 vssd1 vccd1 vccd1 _06132_ sky130_fd_sc_hd__nand2_1
Xhold609 top.CPU.registers.data\[16\] vssd1 vssd1 vccd1 vccd1 net3166 sky130_fd_sc_hd__dlygate4sd3_1
X_11488_ _06618_ net258 net255 net3664 vssd1 vssd1 vccd1 vccd1 _02036_ sky130_fd_sc_hd__a22o_1
XANTENNA__11519__B1 _06734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10990__B2 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16015_ net2349 _02225_ net1095 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[815\]
+ sky130_fd_sc_hd__dfrtp_1
X_13227_ _02782_ _02793_ vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__nor2_1
X_10439_ _05585_ _06062_ net444 vssd1 vssd1 vccd1 vccd1 _06066_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_55_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12192__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13158_ _07414_ _07416_ net1411 net1342 vssd1 vssd1 vccd1 vccd1 _02748_ sky130_fd_sc_hd__a211o_1
XFILLER_111_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12109_ net3886 net651 _06822_ vssd1 vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__o21a_1
X_13089_ top.CPU.data_out\[24\] net2882 net560 vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__mux2_1
XFILLER_100_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1309 top.CPU.registers.data\[898\] vssd1 vssd1 vccd1 vccd1 net3866 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09145__S net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08699__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14465__635 clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 net2104 sky130_fd_sc_hd__inv_2
X_07650_ top.CPU.control_unit.instruction\[5\] _03146_ _03154_ _03263_ net1398 vssd1
+ vssd1 vccd1 vccd1 _03289_ sky130_fd_sc_hd__o311a_1
XANTENNA__08794__S0 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13853__23 clknet_leaf_133_clk vssd1 vssd1 vccd1 vccd1 net1492 sky130_fd_sc_hd__inv_2
XANTENNA__07910__A2 net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07581_ top.CPU.registers.data\[959\] top.CPU.registers.data\[927\] net836 vssd1
+ vssd1 vccd1 vccd1 _03220_ sky130_fd_sc_hd__mux2_1
X_14506__676 clknet_leaf_148_clk vssd1 vssd1 vccd1 vccd1 net2145 sky130_fd_sc_hd__inv_2
XANTENNA__11126__D net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09320_ top.CPU.registers.data\[36\] top.CPU.registers.data\[4\] net829 vssd1 vssd1
+ vccd1 vccd1 _04959_ sky130_fd_sc_hd__mux2_1
XANTENNA__07460__Y _03100_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09663__A2 net1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_103_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16275__Q top.CPU.handler.toreg\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09251_ _04889_ vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11470__A2 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08871__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08202_ top.CPU.registers.data\[823\] top.CPU.registers.data\[791\] net987 vssd1
+ vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__mux2_1
XFILLER_166_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09182_ top.CPU.registers.data\[966\] net1316 net847 top.CPU.registers.data\[998\]
+ net718 vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__a221o_1
XANTENNA__09415__A2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10039__B net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11758__B1 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08133_ top.CPU.registers.data\[853\] net1299 net1020 top.CPU.registers.data\[885\]
+ net941 vssd1 vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__a221o_1
XFILLER_146_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout120_A net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08623__B1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout218_A net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10981__C net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07977__A2 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08064_ top.CPU.registers.data\[820\] top.CPU.registers.data\[788\] net980 vssd1
+ vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__mux2_1
XANTENNA__10326__Y _05958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10055__A net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1127_A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08926__A1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08387__C1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11525__A3 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10733__A1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11930__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08966_ top.CPU.registers.data\[585\] net1309 net840 top.CPU.registers.data\[617\]
+ net761 vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__a221o_1
XANTENNA__08139__C1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11289__A2 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07917_ top.CPU.registers.data\[668\] net1303 net1026 top.CPU.registers.data\[700\]
+ net924 vssd1 vssd1 vccd1 vccd1 _03556_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_162_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout375_X net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08897_ top.CPU.alu.program_counter\[10\] net1033 vssd1 vssd1 vccd1 vccd1 _04536_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__10502__B net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout754_A net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_95_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_95_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08154__A2 net1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07848_ top.CPU.registers.data\[605\] net1288 net1007 top.CPU.registers.data\[637\]
+ net932 vssd1 vssd1 vccd1 vccd1 _03487_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_162_Right_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout921_A net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout542_X net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07779_ top.CPU.registers.data\[574\] net1025 net628 _03417_ vssd1 vssd1 vccd1 vccd1
+ _03418_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout1284_X net1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09103__A1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10249__B1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09518_ _05154_ _05156_ net454 vssd1 vssd1 vccd1 vccd1 _05157_ sky130_fd_sc_hd__mux2_1
X_10790_ _06140_ _06399_ _06400_ _06398_ net411 vssd1 vssd1 vccd1 vccd1 _06401_ sky130_fd_sc_hd__a32o_1
XFILLER_71_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11997__B1 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07665__A1 _03262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09449_ _05087_ vssd1 vssd1 vccd1 vccd1 _05088_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout807_X net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12460_ net448 _05428_ vssd1 vssd1 vccd1 vccd1 _06969_ sky130_fd_sc_hd__and2_1
XANTENNA__11749__B1 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11411_ _06544_ net278 net268 net3138 vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__a22o_1
X_12391_ top.CPU.addressnew\[5\] top.CPU.addressnew\[6\] top.CPU.addressnew\[15\]
+ top.CPU.addressnew\[14\] vssd1 vssd1 vccd1 vccd1 _06929_ sky130_fd_sc_hd__or4_1
XFILLER_138_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13040__S net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16544__RESET_B net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11342_ net3759 net286 net278 _06058_ vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__a22o_1
XFILLER_125_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10972__B2 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11273_ net524 _06374_ net542 vssd1 vssd1 vccd1 vccd1 _06694_ sky130_fd_sc_hd__and3_1
XFILLER_134_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08378__C1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12174__B1 _06749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10224_ _05784_ _05858_ net308 vssd1 vssd1 vccd1 vccd1 _05859_ sky130_fd_sc_hd__mux2_1
X_13012_ top.SPI.paroutput\[7\] _07429_ _07431_ net3064 vssd1 vssd1 vccd1 vccd1 _01213_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09754__A net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14152__322 clknet_leaf_129_clk vssd1 vssd1 vccd1 vccd1 net1791 sky130_fd_sc_hd__inv_2
XANTENNA__11921__B1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10155_ net402 _05791_ vssd1 vssd1 vccd1 vccd1 _05792_ sky130_fd_sc_hd__nand2_1
XFILLER_121_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14449__619 clknet_leaf_186_clk vssd1 vssd1 vccd1 vccd1 net2088 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_50_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10086_ _04158_ _04225_ net378 vssd1 vssd1 vccd1 vccd1 _05724_ sky130_fd_sc_hd__mux2_1
X_14963_ clknet_leaf_93_clk net2703 net1268 vssd1 vssd1 vccd1 vccd1 top.SPI.paroutput\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold6 top.CPU.registers.data_out_r2_prev\[10\] vssd1 vssd1 vccd1 vccd1 net2563 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11508__B net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13674__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12477__B2 _03984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_86_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_86_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09760__Y _05399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07561__X _03200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14884__1054 clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 net2523 sky130_fd_sc_hd__inv_2
X_13776_ net4 net1049 net884 net3846 vssd1 vssd1 vccd1 vccd1 _02657_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_48_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08302__C1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10988_ net3634 net217 _06547_ net315 vssd1 vssd1 vccd1 vccd1 _02354_ sky130_fd_sc_hd__a22o_1
XANTENNA__11988__B1 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15515_ net1849 _01725_ net1214 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[315\]
+ sky130_fd_sc_hd__dfrtp_1
X_12727_ _07186_ _07187_ vssd1 vssd1 vccd1 vccd1 _07188_ sky130_fd_sc_hd__xnor2_1
X_16495_ clknet_leaf_41_clk _02657_ net1116 vssd1 vssd1 vccd1 vccd1 top.mmio.mem_data_i\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10660__B1 _06276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15446_ net1780 _01656_ net1227 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[246\]
+ sky130_fd_sc_hd__dfrtp_1
X_12658_ _03106_ _05232_ vssd1 vssd1 vccd1 vccd1 _07126_ sky130_fd_sc_hd__nor2_1
X_11609_ net141 net3241 net213 vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__mux2_1
XFILLER_129_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15377_ net1711 _01587_ net1191 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[177\]
+ sky130_fd_sc_hd__dfrtp_1
X_12589_ top.CPU.handler.readout _07054_ _07090_ _03132_ vssd1 vssd1 vccd1 vccd1 _07091_
+ sky130_fd_sc_hd__a211o_1
XANTENNA__09802__C1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_10_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__16285__RESET_B net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07959__A2 net1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold406 top.CPU.registers.data\[389\] vssd1 vssd1 vccd1 vccd1 net2963 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold417 top.CPU.registers.data\[818\] vssd1 vssd1 vccd1 vccd1 net2974 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold428 top.CPU.registers.data\[339\] vssd1 vssd1 vccd1 vccd1 net2985 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold439 top.CPU.registers.data\[422\] vssd1 vssd1 vccd1 vccd1 net2996 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09256__S1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10306__C _05937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09030__B1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout908 net909 vssd1 vssd1 vccd1 vccd1 net908 sky130_fd_sc_hd__clkbuf_4
Xfanout919 net920 vssd1 vssd1 vccd1 vccd1 net919 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11912__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09581__A1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08820_ _03342_ _04445_ _04458_ vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__o21ai_4
XFILLER_140_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12180__A3 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07592__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1106 top.CPU.registers.data\[620\] vssd1 vssd1 vccd1 vccd1 net3663 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1117 top.CPU.registers.data\[329\] vssd1 vssd1 vccd1 vccd1 net3674 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1128 top.CPU.registers.data\[835\] vssd1 vssd1 vccd1 vccd1 net3685 sky130_fd_sc_hd__dlygate4sd3_1
X_08751_ _03342_ _04378_ _04389_ vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__o21a_2
XANTENNA__12468__A1 _03754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12468__B2 _03915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1139 top.CPU.registers.data\[522\] vssd1 vssd1 vccd1 vccd1 net3696 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_77_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09333__A1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10479__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07702_ top.CPU.registers.data\[639\] top.CPU.registers.data\[607\] net999 vssd1
+ vssd1 vccd1 vccd1 _03341_ sky130_fd_sc_hd__mux2_1
XFILLER_39_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08682_ net1368 _04313_ _04312_ top.CPU.control_unit.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 _04321_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_68_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09603__S net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07633_ top.CPU.control_unit.instruction\[14\] _03108_ net1400 vssd1 vssd1 vccd1
+ vccd1 _03272_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07895__A1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13417__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11691__A2 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout168_A net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07564_ net1048 _03164_ net1039 net1390 vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__o31a_4
XFILLER_110_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11979__B1 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09303_ net940 _04939_ _04941_ net957 vssd1 vssd1 vccd1 vccd1 _04942_ sky130_fd_sc_hd__o211a_1
XANTENNA__11153__B net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07495_ net4012 vssd1 vssd1 vccd1 vccd1 _03135_ sky130_fd_sc_hd__inv_2
XFILLER_21_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout335_A _03047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10651__B1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09234_ top.CPU.registers.data\[421\] net1386 net806 top.CPU.registers.data\[389\]
+ net690 vssd1 vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14593__763 clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 net2232 sky130_fd_sc_hd__inv_2
XFILLER_148_952 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09165_ net789 _04802_ _04803_ net704 vssd1 vssd1 vccd1 vccd1 _04804_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout123_X net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout502_A _05696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1244_A net1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08116_ net1035 _03754_ _03724_ vssd1 vssd1 vccd1 vccd1 _03755_ sky130_fd_sc_hd__a21oi_4
XANTENNA__10403__B1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09096_ top.CPU.registers.data\[327\] net1333 net863 top.CPU.registers.data\[359\]
+ net778 vssd1 vssd1 vccd1 vccd1 _04735_ sky130_fd_sc_hd__a221o_1
XANTENNA__10954__B2 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08047_ top.CPU.registers.data\[52\] net1008 net931 vssd1 vssd1 vccd1 vccd1 _03686_
+ sky130_fd_sc_hd__a21o_1
Xhold940 _02702_ vssd1 vssd1 vccd1 vccd1 net3497 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1032_X net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14136__306 clknet_leaf_167_clk vssd1 vssd1 vccd1 vccd1 net1775 sky130_fd_sc_hd__inv_2
XFILLER_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12156__B1 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold951 top.CPU.registers.data\[920\] vssd1 vssd1 vccd1 vccd1 net3508 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold962 top.CPU.registers.data\[373\] vssd1 vssd1 vccd1 vccd1 net3519 sky130_fd_sc_hd__dlygate4sd3_1
Xhold973 top.CPU.registers.data\[627\] vssd1 vssd1 vccd1 vccd1 net3530 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_164_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold984 top.CPU.registers.data\[196\] vssd1 vssd1 vccd1 vccd1 net3541 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_164_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold995 top.CPU.handler.toreg\[9\] vssd1 vssd1 vccd1 vccd1 net3552 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout492_X net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout871_A net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout969_A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11903__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09998_ _04225_ _04294_ net378 vssd1 vssd1 vccd1 vccd1 _05637_ sky130_fd_sc_hd__mux2_1
XFILLER_95_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08780__C1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08949_ top.CPU.registers.data\[1002\] top.CPU.registers.data\[970\] net971 vssd1
+ vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_68_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout757_X net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13120__A2 net1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10800__X _06411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11960_ _06507_ net341 net229 net3434 vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__a22o_1
XANTENNA__11131__A1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_174_Left_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10911_ net486 net516 _06500_ vssd1 vssd1 vccd1 vccd1 _06501_ sky130_fd_sc_hd__and3_1
XANTENNA__07886__A1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11891_ _06354_ net3252 net189 vssd1 vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout924_X net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13630_ net3908 _03100_ net663 vssd1 vssd1 vccd1 vccd1 _02564_ sky130_fd_sc_hd__mux2_1
X_10842_ _03374_ _05609_ _05604_ vssd1 vssd1 vccd1 vccd1 _06450_ sky130_fd_sc_hd__a21o_1
XFILLER_44_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13561_ net1348 _06371_ vssd1 vssd1 vccd1 vccd1 _03003_ sky130_fd_sc_hd__nand2_1
X_10773_ _04989_ _05685_ net443 vssd1 vssd1 vccd1 vccd1 _06385_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08835__B1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15300_ net1634 _01510_ net1185 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[100\]
+ sky130_fd_sc_hd__dfrtp_1
X_12512_ net450 _04461_ _07018_ _07019_ _07020_ vssd1 vssd1 vccd1 vccd1 _07021_ sky130_fd_sc_hd__o2111a_1
X_16280_ clknet_leaf_60_clk _02490_ net1139 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.toreg\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_13492_ top.CPU.data_out\[6\] _04855_ net587 vssd1 vssd1 vccd1 vccd1 _02504_ sky130_fd_sc_hd__mux2_1
XANTENNA__08653__A _04291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15231_ net1565 _01441_ net1203 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_12443_ net1339 top.I2C.output_state\[3\] net3053 vssd1 vssd1 vccd1 vccd1 _06958_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_23_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11198__B2 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15162_ clknet_leaf_44_clk _01372_ net1124 vssd1 vssd1 vccd1 vccd1 top.I2C.data_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11737__A3 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12374_ top.I2C.output_state\[14\] _06912_ vssd1 vssd1 vccd1 vccd1 _06914_ sky130_fd_sc_hd__nand2_1
XANTENNA__09260__B1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11510__C _06731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10407__B net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10945__B2 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11325_ net3470 net291 net359 _06428_ vssd1 vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__a22o_1
X_15093_ net1475 _01306_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r2_prev\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08799__S net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12147__B1 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11256_ net473 _06683_ vssd1 vssd1 vccd1 vccd1 _06684_ sky130_fd_sc_hd__nor2_1
X_10207_ _05618_ _05824_ _05842_ vssd1 vssd1 vccd1 vccd1 _05843_ sky130_fd_sc_hd__o21ai_1
X_11187_ net1401 net485 _06652_ net298 net3350 vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__a32o_1
XANTENNA__11370__A1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10138_ net381 _05546_ _05622_ vssd1 vssd1 vccd1 vccd1 _05775_ sky130_fd_sc_hd__or3_1
XANTENNA__11238__B net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15995_ net2329 _02205_ net1213 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[795\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_59_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_94_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14946_ clknet_leaf_65_clk _01192_ net1163 vssd1 vssd1 vccd1 vccd1 top.CPU.alu.program_counter\[29\]
+ sky130_fd_sc_hd__dfrtp_2
X_10069_ net382 _05705_ _05706_ vssd1 vssd1 vccd1 vccd1 _05707_ sky130_fd_sc_hd__or3_1
XFILLER_85_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16616_ net1347 vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__clkbuf_1
X_13828_ net2927 net337 net329 top.CPU.data_out\[30\] vssd1 vssd1 vccd1 vccd1 _02708_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09079__B1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12069__B net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14280__450 clknet_leaf_129_clk vssd1 vssd1 vccd1 vccd1 net1919 sky130_fd_sc_hd__inv_2
X_16547_ clknet_leaf_92_clk _02709_ net1270 vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13759_ _02803_ _03089_ _03091_ top.I2C.which_data_address\[1\] vssd1 vssd1 vccd1
+ vccd1 _02644_ sky130_fd_sc_hd__o22a_1
XANTENNA__11425__A2 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14577__747 clknet_leaf_186_clk vssd1 vssd1 vccd1 vccd1 net2216 sky130_fd_sc_hd__inv_2
XFILLER_93_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16478_ clknet_leaf_89_clk _02640_ net1274 vssd1 vssd1 vccd1 vccd1 top.SPI.timem\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_15429_ net1763 _01639_ net1083 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[229\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14321__491 clknet_leaf_180_clk vssd1 vssd1 vccd1 vccd1 net1960 sky130_fd_sc_hd__inv_2
XANTENNA__11189__B2 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14618__788 clknet_leaf_162_clk vssd1 vssd1 vccd1 vccd1 net2257 sky130_fd_sc_hd__inv_2
XANTENNA__08054__A1 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold203 top.CPU.registers.data\[684\] vssd1 vssd1 vccd1 vccd1 net2760 sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 top.CPU.registers.data\[415\] vssd1 vssd1 vccd1 vccd1 net2771 sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 top.I2C.I2C_state\[12\] vssd1 vssd1 vccd1 vccd1 net2782 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07801__A1 _03409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold236 top.CPU.registers.data\[168\] vssd1 vssd1 vccd1 vccd1 net2793 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_160_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12138__B1 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold247 top.CPU.registers.data\[537\] vssd1 vssd1 vccd1 vccd1 net2804 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold258 top.CPU.registers.data\[699\] vssd1 vssd1 vccd1 vccd1 net2815 sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ _04829_ _04858_ vssd1 vssd1 vccd1 vccd1 _05560_ sky130_fd_sc_hd__and2_1
Xhold269 top.CPU.registers.data\[472\] vssd1 vssd1 vccd1 vccd1 net2826 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_113_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout705 net706 vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__clkbuf_2
Xfanout716 net717 vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__clkbuf_4
Xfanout727 net735 vssd1 vssd1 vccd1 vccd1 net727 sky130_fd_sc_hd__clkbuf_4
X_09852_ top.CPU.registers.data\[314\] net1027 net945 vssd1 vssd1 vccd1 vccd1 _05491_
+ sky130_fd_sc_hd__a21o_1
Xfanout738 net739 vssd1 vssd1 vccd1 vccd1 net738 sky130_fd_sc_hd__clkbuf_4
XFILLER_58_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07565__B1 net1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout749 net760 vssd1 vssd1 vccd1 vccd1 net749 sky130_fd_sc_hd__clkbuf_4
XFILLER_105_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08762__C1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08803_ top.CPU.registers.data\[204\] net1372 net977 top.CPU.registers.data\[236\]
+ net926 vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_142_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ net607 _05419_ _05420_ _05421_ net623 vssd1 vssd1 vccd1 vccd1 _05422_ sky130_fd_sc_hd__o311a_1
XANTENNA__08109__A2 net1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout285_A _06712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08734_ _04371_ _04372_ net927 vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__mux2_1
XANTENNA__11113__A1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08514__C1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08665_ _04302_ _04303_ net934 vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout452_A net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11164__A net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07616_ net1400 _03148_ _03245_ net882 vssd1 vssd1 vccd1 vccd1 _03255_ sky130_fd_sc_hd__or4b_2
X_08596_ _04233_ _04234_ net929 vssd1 vssd1 vccd1 vccd1 _04235_ sky130_fd_sc_hd__mux2_1
XFILLER_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11416__A2 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07547_ top.CPU.control_unit.instruction\[11\] _03184_ vssd1 vssd1 vccd1 vccd1 _03186_
+ sky130_fd_sc_hd__and2_2
XANTENNA_fanout240_X net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1361_A net1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout338_X net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout717_A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07478_ net1361 vssd1 vssd1 vccd1 vccd1 _03118_ sky130_fd_sc_hd__inv_2
XFILLER_10_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09217_ top.CPU.control_unit.instruction\[26\] _04596_ _04597_ vssd1 vssd1 vccd1
+ vccd1 _04856_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout505_X net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_118_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08045__A1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09148_ top.CPU.registers.data\[967\] net1296 net1016 top.CPU.registers.data\[999\]
+ net913 vssd1 vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_135_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09242__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09079_ top.CPU.registers.data\[552\] net975 net903 _04717_ vssd1 vssd1 vccd1 vccd1
+ _04718_ sky130_fd_sc_hd__o211a_1
XFILLER_146_33 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12723__A top.CPU.alu.program_counter\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14883__1053 clknet_leaf_171_clk vssd1 vssd1 vccd1 vccd1 net2522 sky130_fd_sc_hd__inv_2
X_11110_ net1406 net577 net528 net134 vssd1 vssd1 vccd1 vccd1 _06613_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_9_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12090_ net3988 net646 _06813_ vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__o21a_1
XANTENNA__08412__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold770 top.CPU.registers.data\[533\] vssd1 vssd1 vccd1 vccd1 net3327 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout874_X net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold781 top.CPU.registers.data\[338\] vssd1 vssd1 vccd1 vccd1 net3338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold792 top.SPI.parameters\[12\] vssd1 vssd1 vccd1 vccd1 net3349 sky130_fd_sc_hd__dlygate4sd3_1
X_11041_ net325 net135 net538 net368 net2869 vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__a32o_1
XFILLER_77_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07536__B net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12869__S net1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15780_ net2114 _01990_ net1186 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[580\]
+ sky130_fd_sc_hd__dfrtp_1
X_12992_ top.SPI.state\[5\] top.SPI.state\[3\] top.SPI.state\[4\] vssd1 vssd1 vccd1
+ vccd1 _07421_ sky130_fd_sc_hd__or3_1
XFILLER_29_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10897__B net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08505__C1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1470 top.CPU.data_out\[5\] vssd1 vssd1 vccd1 vccd1 net4027 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input13_A DAT_I[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11943_ _06486_ net347 net231 net3305 vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__a22o_1
XANTENNA__07859__A1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11655__A2 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14264__434 clknet_leaf_168_clk vssd1 vssd1 vccd1 vccd1 net1903 sky130_fd_sc_hd__inv_2
XANTENNA__08520__A2 _04155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12488__A1_N _04566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11874_ net134 net3472 net190 vssd1 vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16401_ clknet_leaf_62_clk _00024_ net1161 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.state\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_28_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13613_ top.CPU.alu.program_counter\[25\] _05931_ net1351 vssd1 vssd1 vccd1 vccd1
+ _03035_ sky130_fd_sc_hd__mux2_1
X_10825_ _05194_ _05670_ vssd1 vssd1 vccd1 vccd1 _06434_ sky130_fd_sc_hd__nand2_1
XANTENNA__08808__B1 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11407__A2 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11224__D net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16332_ clknet_leaf_68_clk _02541_ net1167 vssd1 vssd1 vccd1 vccd1 top.CPU.addressnew\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_14305__475 clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 net1944 sky130_fd_sc_hd__inv_2
X_13544_ top.CPU.data_out\[30\] net590 _02992_ vssd1 vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__o21a_1
X_10756_ net549 _05543_ _06367_ _06368_ vssd1 vssd1 vccd1 vccd1 _06369_ sky130_fd_sc_hd__o211a_1
XANTENNA__12080__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16263_ clknet_leaf_44_clk _02473_ net1124 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.toreg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11521__B net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13475_ net1397 net873 _02924_ net418 vssd1 vssd1 vccd1 vccd1 _02959_ sky130_fd_sc_hd__a31o_1
X_10687_ _04730_ net503 net443 vssd1 vssd1 vccd1 vccd1 _06303_ sky130_fd_sc_hd__o21ai_1
XFILLER_139_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15214_ net1548 _01424_ net1190 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_12426_ top.I2C.read_byte_done top.I2C.reader_state\[0\] vssd1 vssd1 vccd1 vccd1
+ _06950_ sky130_fd_sc_hd__nor2_1
XFILLER_145_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08036__A1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16194_ net2528 _02404_ net1174 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[994\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09233__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11240__C net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10918__A1 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08587__A2 _04222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09784__A1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15145_ clknet_leaf_47_clk _01355_ net1130 vssd1 vssd1 vccd1 vccd1 top.I2C.data_out\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_12357_ net1054 _06900_ vssd1 vssd1 vccd1 vccd1 _00061_ sky130_fd_sc_hd__and2_1
XFILLER_127_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07795__B1 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08992__C1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11308_ net3157 net289 net359 net139 vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__a22o_1
X_15076_ clknet_leaf_51_clk _00054_ net1134 vssd1 vssd1 vccd1 vccd1 top.I2C.output_state\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12288_ net3863 _03956_ net1177 vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__mux2_1
XANTENNA__13332__A2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11249__A net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11239_ net3423 net294 _06674_ net485 vssd1 vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__a22o_1
XFILLER_110_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08744__C1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09942__A _03755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15441__RESET_B net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15978_ net2312 _02188_ net1084 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[778\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16548__Q net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14929_ clknet_leaf_63_clk _01175_ net1161 vssd1 vssd1 vccd1 vccd1 top.CPU.alu.program_counter\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_64_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11646__A2 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10854__B1 _06461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08450_ net800 _04081_ _04088_ net642 vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__a211o_1
XFILLER_36_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08381_ net880 _04019_ _03990_ vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__o21a_1
XFILLER_91_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10606__B1 _06223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08275__A1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12071__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11431__B net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09002_ top.CPU.registers.data\[1001\] top.CPU.registers.data\[969\] net965 vssd1
+ vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_152_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08122__S1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12543__A net1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout200_A net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07786__B1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11582__B2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09527__A1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09904_ _05542_ vssd1 vssd1 vccd1 vccd1 _05543_ sky130_fd_sc_hd__inv_2
Xfanout502 _05696_ vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__buf_2
XANTENNA__11159__A net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout513 net514 vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__clkbuf_4
Xfanout524 net533 vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__buf_4
XFILLER_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08735__C1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout535 net537 vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__clkbuf_4
XFILLER_101_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout546 _06523_ vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__buf_4
XFILLER_58_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout557 _07418_ vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input5_A DAT_I[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09835_ net682 _05472_ _05473_ net609 vssd1 vssd1 vccd1 vccd1 _05474_ sky130_fd_sc_hd__a31o_1
Xfanout568 net569 vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__clkbuf_4
Xfanout579 _02995_ vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__buf_2
XANTENNA__10998__A net1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout190_X net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout667_A net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout288_X net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09766_ top.CPU.registers.data\[475\] net1298 net1019 top.CPU.registers.data\[507\]
+ net916 vssd1 vssd1 vccd1 vccd1 _05405_ sky130_fd_sc_hd__a221o_1
XFILLER_101_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14248__418 clknet_leaf_126_clk vssd1 vssd1 vccd1 vccd1 net1887 sky130_fd_sc_hd__inv_2
XFILLER_67_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08717_ net784 _04352_ _04353_ net714 vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__o211a_1
XANTENNA__11637__A2 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout834_A net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09697_ top.CPU.registers.data\[921\] net1306 net1029 top.CPU.registers.data\[953\]
+ net922 vssd1 vssd1 vccd1 vccd1 _05336_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout455_X net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08502__A2 net1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10002__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08648_ top.CPU.registers.data\[430\] top.CPU.registers.data\[398\] net818 vssd1
+ vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__mux2_1
XFILLER_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16317__RESET_B net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08579_ top.CPU.registers.data\[431\] net1387 net812 top.CPU.registers.data\[399\]
+ net716 vssd1 vssd1 vccd1 vccd1 _04218_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout622_X net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1364_X net1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10610_ net600 _06228_ _06229_ vssd1 vssd1 vccd1 vccd1 _06230_ sky130_fd_sc_hd__o21ai_4
XTAP_TAPCELL_ROW_137_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11590_ net565 _03182_ net362 vssd1 vssd1 vccd1 vccd1 _06749_ sky130_fd_sc_hd__and3_4
XANTENNA__12062__A2 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10541_ net397 _06163_ _06161_ vssd1 vssd1 vccd1 vccd1 _06164_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_133_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13260_ net892 top.I2C.data_out\[6\] _02787_ vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__mux2_1
X_10472_ _05887_ _06090_ net403 vssd1 vssd1 vccd1 vccd1 _06098_ sky130_fd_sc_hd__mux2_1
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout991_X net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08569__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12211_ net3821 net647 _06872_ vssd1 vssd1 vccd1 vccd1 _01456_ sky130_fd_sc_hd__o21a_1
XFILLER_68_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13191_ _02770_ _02771_ net3882 vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__a21o_1
XANTENNA__10525__X _06149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11573__B2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12142_ top.CPU.registers.data\[81\] net652 net244 vssd1 vssd1 vccd1 vccd1 _06839_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__07547__A top.CPU.control_unit.instruction\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_29_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10244__Y _05879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09518__A1 _05156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11069__A net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12073_ top.CPU.registers.data\[116\] net649 net361 vssd1 vssd1 vccd1 vccd1 _06805_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__11325__B2 _06428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11024_ net3789 net216 _06569_ net316 vssd1 vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__a22o_1
X_15901_ net2235 _02111_ net1121 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[701\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15832_ net2166 _02042_ net1148 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[632\]
+ sky130_fd_sc_hd__dfrtp_1
X_15763_ net2097 _01973_ net1198 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[563\]
+ sky130_fd_sc_hd__dfrtp_1
X_12975_ _07409_ top.I2C.bit_timer_state\[0\] _07408_ vssd1 vssd1 vccd1 vccd1 _01198_
+ sky130_fd_sc_hd__and3b_1
XANTENNA__13571__X _03009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11926_ net3857 net184 net344 _06357_ vssd1 vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__a22o_1
X_15694_ net2028 _01904_ net1104 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[494\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1038 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11857_ net459 _06693_ net235 net153 net2651 vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__a32o_1
XFILLER_60_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11091__X _06602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10808_ net409 _06263_ _06417_ net416 vssd1 vssd1 vccd1 vccd1 _06418_ sky130_fd_sc_hd__a211oi_1
XANTENNA__12053__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13250__B2 _02803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11788_ _06634_ net198 net160 net3293 vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__a22o_1
XFILLER_14_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16315_ clknet_leaf_83_clk _02524_ net1261 vssd1 vssd1 vccd1 vccd1 top.CPU.data_out\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13527_ _03915_ net584 vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__and2_1
XANTENNA__08352__S1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10739_ top.CPU.fetch.current_ra\[6\] net1040 net881 top.CPU.handler.toreg\[6\] vssd1
+ vssd1 vccd1 vccd1 _06353_ sky130_fd_sc_hd__a22o_1
XFILLER_159_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11800__A2 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16246_ clknet_leaf_43_clk _02456_ net1123 vssd1 vssd1 vccd1 vccd1 top.CPU.control_unit.instruction\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_173_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13458_ top.CPU.handler.toreg\[18\] _02950_ net123 vssd1 vssd1 vccd1 vccd1 _02484_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09206__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09757__A1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12409_ _06918_ _06925_ _06934_ vssd1 vssd1 vccd1 vccd1 _06935_ sky130_fd_sc_hd__or3_1
X_14392__562 clknet_leaf_160_clk vssd1 vssd1 vccd1 vccd1 net2031 sky130_fd_sc_hd__inv_2
X_16177_ net2511 _02387_ net1176 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[977\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 WE_O sky130_fd_sc_hd__buf_2
X_13389_ net888 _02909_ vssd1 vssd1 vccd1 vccd1 _02910_ sky130_fd_sc_hd__and2_1
XFILLER_127_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput116 net116 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__buf_2
XFILLER_56_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14689__859 clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 net2328 sky130_fd_sc_hd__inv_2
XFILLER_126_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15128_ clknet_leaf_57_clk _01338_ net1144 vssd1 vssd1 vccd1 vccd1 top.I2C.within_byte_counter_writing\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_114_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15059_ clknet_leaf_50_clk _00063_ net1129 vssd1 vssd1 vccd1 vccd1 top.I2C.output_state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_07950_ top.CPU.registers.data\[408\] net820 net793 _03588_ vssd1 vssd1 vccd1 vccd1
+ _03589_ sky130_fd_sc_hd__a211o_1
XANTENNA__08987__S net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11316__B2 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08717__C1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07891__S net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07881_ top.CPU.registers.data\[764\] net1394 net832 top.CPU.registers.data\[732\]
+ net729 vssd1 vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_71_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08193__B1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09620_ net741 _05257_ _05258_ net765 vssd1 vssd1 vccd1 vccd1 _05259_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_71_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07904__B net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10611__A net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16278__Q top.CPU.handler.toreg\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09551_ top.CPU.registers.data_out_r1_prev\[1\] net876 net638 _05189_ _05174_ vssd1
+ vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__o221ai_4
XFILLER_83_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07623__C _03154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09142__C1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08502_ top.CPU.registers.data\[592\] net1321 net852 top.CPU.registers.data\[624\]
+ net745 vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__a221o_1
XFILLER_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08496__A1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09482_ _05120_ vssd1 vssd1 vccd1 vccd1 _05121_ sky130_fd_sc_hd__inv_2
XFILLER_63_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14882__1052 clknet_leaf_143_clk vssd1 vssd1 vccd1 vccd1 net2521 sky130_fd_sc_hd__inv_2
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08433_ net796 _04061_ _04062_ net725 vssd1 vssd1 vccd1 vccd1 _04072_ sky130_fd_sc_hd__o211a_1
XFILLER_24_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout150_A _06780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout248_A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08248__A1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08364_ net790 _03999_ _04002_ net641 vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__a31o_1
XANTENNA__12044__A2 _06779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08227__S net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09996__A1 _04634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11161__B net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11252__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13792__A2 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08295_ net796 _03928_ _03929_ net724 vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__o211a_1
XANTENNA__10058__A net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout415_A net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14633__803 clknet_leaf_154_clk vssd1 vssd1 vccd1 vccd1 net2272 sky130_fd_sc_hd__inv_2
XANTENNA_fanout1157_A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13544__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12273__A _06887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout203_X net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1324_A net1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15363__RESET_B net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout784_A net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout310 _05158_ vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__buf_2
Xfanout1308 _03110_ vssd1 vssd1 vccd1 vccd1 net1308 sky130_fd_sc_hd__clkbuf_8
Xfanout321 net322 vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__buf_4
XANTENNA__11307__B2 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1319 net1323 vssd1 vssd1 vccd1 vccd1 net1319 sky130_fd_sc_hd__clkbuf_4
Xfanout332 _03047_ vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__clkbuf_2
Xfanout343 _06771_ vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11858__A2 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout354 net356 vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout572_X net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout951_A net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08184__B1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout365 _06600_ vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__clkbuf_8
Xfanout376 _05235_ vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__clkbuf_4
Xfanout387 net393 vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__clkbuf_4
X_09818_ net698 _05454_ _05455_ _05456_ vssd1 vssd1 vccd1 vccd1 _05457_ sky130_fd_sc_hd__a31o_1
XFILLER_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout398 _05089_ vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07931__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09749_ net799 _05386_ _05387_ net727 vssd1 vssd1 vccd1 vccd1 _05388_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout837_X net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10818__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12760_ _07215_ _07216_ _07204_ vssd1 vssd1 vccd1 vccd1 _07218_ sky130_fd_sc_hd__or3b_2
XANTENNA__11055__C net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_6_Left_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09521__S net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _06547_ net202 net421 net2818 vssd1 vssd1 vccd1 vccd1 _01842_ sky130_fd_sc_hd__a22o_1
XANTENNA__07830__A net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07695__C1 net1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11491__B1 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12691_ top.CPU.alu.program_counter\[5\] _07155_ net1360 vssd1 vssd1 vccd1 vccd1
+ _01168_ sky130_fd_sc_hd__mux2_1
XFILLER_159_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12448__A net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11642_ _06086_ net205 net426 net3342 vssd1 vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__a22o_1
XANTENNA__12035__A2 _06780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11071__B net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11573_ net3001 net246 _06744_ net483 vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__a22o_1
Xinput18 DAT_I[24] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
X_16100_ net2434 _02310_ net1185 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[900\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_156_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13312_ net1343 top.mmio.mem_data_i\[2\] net596 vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__o21a_1
X_14376__546 clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 net2015 sky130_fd_sc_hd__inv_2
X_10524_ top.CPU.fetch.current_ra\[16\] net1043 net634 top.CPU.handler.toreg\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06148_ sky130_fd_sc_hd__a22o_1
Xinput29 DAT_I[5] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_168_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13929__99 clknet_leaf_159_clk vssd1 vssd1 vccd1 vccd1 net1568 sky130_fd_sc_hd__inv_2
XANTENNA__08661__A net1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16031_ net2365 _02241_ net1225 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[831\]
+ sky130_fd_sc_hd__dfrtp_1
X_13243_ net893 top.I2C.data_out\[14\] _02787_ vssd1 vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__mux2_1
X_10455_ _06067_ _06081_ net600 vssd1 vssd1 vccd1 vccd1 _06082_ sky130_fd_sc_hd__a21o_1
XANTENNA__10349__A2 _05670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12743__A0 top.CPU.control_unit.instruction\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14120__290 clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 net1759 sky130_fd_sc_hd__inv_2
X_13174_ _02757_ _02756_ top.I2C.within_byte_counter_writing\[0\] vssd1 vssd1 vccd1
+ vccd1 _01337_ sky130_fd_sc_hd__mux2_1
X_14417__587 clknet_leaf_186_clk vssd1 vssd1 vccd1 vccd1 net2056 sky130_fd_sc_hd__inv_2
X_10386_ _05674_ _06014_ net410 vssd1 vssd1 vccd1 vccd1 _06015_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_92_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13566__X _03006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12125_ net3971 net175 _06830_ _06480_ vssd1 vssd1 vccd1 vccd1 _01500_ sky130_fd_sc_hd__a22o_1
XFILLER_124_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10134__C net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07564__X _03203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12056_ _06729_ net235 net177 net3351 vssd1 vssd1 vccd1 vccd1 _01535_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_53_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11007_ net513 _06312_ net542 vssd1 vssd1 vccd1 vccd1 _06559_ sky130_fd_sc_hd__and3_1
XANTENNA__08714__A2 net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10521__A2 _05669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07922__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15815_ net2149 _02025_ net1197 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[615\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_37_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15746_ net2080 _01956_ net1171 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[546\]
+ sky130_fd_sc_hd__dfrtp_1
X_12958_ top.CPU.alu.program_counter\[30\] _03409_ _07386_ _07396_ vssd1 vssd1 vccd1
+ vccd1 _07397_ sky130_fd_sc_hd__a211o_1
XANTENNA__13471__A1 net1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11909_ net3933 net185 net347 _05991_ vssd1 vssd1 vccd1 vccd1 _01657_ sky130_fd_sc_hd__a22o_1
XANTENNA__11482__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10577__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15677_ net2011 _01887_ net1112 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[477\]
+ sky130_fd_sc_hd__dfrtp_1
X_12889_ net126 _07334_ net1359 vssd1 vssd1 vccd1 vccd1 _07335_ sky130_fd_sc_hd__o21a_1
X_13984__154 clknet_leaf_125_clk vssd1 vssd1 vccd1 vccd1 net1623 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12077__B net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08080_ _03683_ _03718_ vssd1 vssd1 vccd1 vccd1 _03719_ sky130_fd_sc_hd__nand2_1
X_16229_ clknet_leaf_31_clk _02439_ net1125 vssd1 vssd1 vccd1 vccd1 top.CPU.control_unit.instruction\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_161_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11537__A1 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08938__C1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11201__S net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08402__A1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_755 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07618__C top.CPU.control_unit.instruction\[29\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12380__X _06918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08982_ net783 _04619_ _04620_ net737 vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__o211a_1
XFILLER_142_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_143_Right_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07933_ net683 _03570_ _03571_ net608 vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__a31o_1
XFILLER_130_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08166__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10979__C net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout198_A net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07634__B net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12032__S net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07864_ top.CPU.registers.data\[349\] net1289 net1007 top.CPU.registers.data\[381\]
+ net931 vssd1 vssd1 vccd1 vccd1 _03503_ sky130_fd_sc_hd__a221o_1
XFILLER_113_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09603_ top.CPU.registers.data\[416\] top.CPU.registers.data\[384\] net810 vssd1
+ vssd1 vccd1 vccd1 _05242_ sky130_fd_sc_hd__mux2_1
XANTENNA__11156__B net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07795_ top.CPU.registers.data\[254\] net1384 net996 top.CPU.registers.data\[222\]
+ net920 vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__a221o_1
X_09534_ net757 _05169_ _05172_ net710 vssd1 vssd1 vccd1 vccd1 _05173_ sky130_fd_sc_hd__a211o_1
XFILLER_37_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11068__A3 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09666__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08746__A net1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10487__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09465_ net695 _05102_ _05103_ vssd1 vssd1 vccd1 vccd1 _05104_ sky130_fd_sc_hd__or3_1
XFILLER_58_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout153_X net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout532_A net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1274_A net1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08416_ _03988_ _04054_ vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__nand2_1
X_14063__233 clknet_leaf_191_clk vssd1 vssd1 vccd1 vccd1 net1702 sky130_fd_sc_hd__inv_2
XANTENNA__12017__A2 net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09396_ net708 _05033_ _05034_ vssd1 vssd1 vccd1 vccd1 _05035_ sky130_fd_sc_hd__or3_1
XANTENNA__10059__Y _05697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11225__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08347_ top.CPU.control_unit.instruction\[19\] _03160_ _03985_ vssd1 vssd1 vccd1
+ vccd1 _03986_ sky130_fd_sc_hd__o21a_2
XFILLER_11_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout320_X net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout418_X net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08752__Y _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11900__A net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08278_ _03915_ _03916_ net455 vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__mux2_1
X_14104__274 clknet_leaf_167_clk vssd1 vssd1 vccd1 vccd1 net1743 sky130_fd_sc_hd__inv_2
XANTENNA__12715__B _04728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout999_A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10516__A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1327_X net1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10240_ _05617_ _05872_ _05874_ _05868_ vssd1 vssd1 vccd1 vccd1 _05875_ sky130_fd_sc_hd__a211o_1
XFILLER_145_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout787_X net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10171_ net603 _05806_ _05807_ vssd1 vssd1 vccd1 vccd1 _05808_ sky130_fd_sc_hd__a21o_4
XANTENNA__08944__A2 net1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12731__A top.CPU.alu.program_counter\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_110_Right_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1105 net1109 vssd1 vssd1 vccd1 vccd1 net1105 sky130_fd_sc_hd__clkbuf_4
XFILLER_152_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1116 net1118 vssd1 vssd1 vccd1 vccd1 net1116 sky130_fd_sc_hd__clkbuf_2
Xfanout1127 net1147 vssd1 vssd1 vccd1 vccd1 net1127 sky130_fd_sc_hd__clkbuf_2
XFILLER_154_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1138 net1140 vssd1 vssd1 vccd1 vccd1 net1138 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout954_X net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout140 _06126_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__buf_1
Xfanout1149 net1151 vssd1 vssd1 vccd1 vccd1 net1149 sky130_fd_sc_hd__clkbuf_2
Xfanout151 _06780_ vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__buf_6
XANTENNA__13038__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09354__C1 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout162 _06760_ vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__clkbuf_8
X_14761__931 clknet_leaf_158_clk vssd1 vssd1 vccd1 vccd1 net2400 sky130_fd_sc_hd__inv_2
XANTENNA__10889__C _06471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout173 _06825_ vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__buf_2
Xfanout184 net187 vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__clkbuf_8
Xfanout195 _06759_ vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__buf_4
XANTENNA__10503__A2 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_190_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08927__Y _04566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09106__C1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15600_ net1934 _01810_ net1108 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[400\]
+ sky130_fd_sc_hd__dfrtp_1
X_12812_ top.CPU.alu.program_counter\[17\] _04123_ vssd1 vssd1 vccd1 vccd1 _07265_
+ sky130_fd_sc_hd__or2_1
X_13792_ net21 net1050 net885 net2772 vssd1 vssd1 vccd1 vccd1 _02673_ sky130_fd_sc_hd__o22a_1
XANTENNA__13453__A1 net1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14802__972 clknet_leaf_193_clk vssd1 vssd1 vccd1 vccd1 net2441 sky130_fd_sc_hd__inv_2
XANTENNA__11059__A3 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13968__138 clknet_leaf_200_clk vssd1 vssd1 vccd1 vccd1 net1607 sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_70_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15531_ net1865 _01741_ net1058 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[331\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11464__A0 _06311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12743_ top.CPU.control_unit.instruction\[7\] _07201_ _03251_ vssd1 vssd1 vccd1 vccd1
+ _07202_ sky130_fd_sc_hd__mux2_1
XANTENNA__10397__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15462_ net1796 _01672_ net1074 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[262\]
+ sky130_fd_sc_hd__dfrtp_1
X_12674_ _07132_ _07133_ _07130_ vssd1 vssd1 vccd1 vccd1 _07140_ sky130_fd_sc_hd__a21bo_1
XANTENNA__12008__A2 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10019__A1 _05332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11625_ _06428_ net3511 net212 vssd1 vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__mux2_1
XFILLER_168_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09758__Y _05397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15393_ net1727 _01603_ net1230 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[193\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11232__D net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_85_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11767__A1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11556_ net494 net476 _06669_ net248 net2646 vssd1 vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_94_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10507_ _05752_ _05937_ _05643_ vssd1 vssd1 vccd1 vccd1 _06131_ sky130_fd_sc_hd__o21a_1
X_11487_ net565 net488 _06617_ net256 net3530 vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__a32o_1
XANTENNA__10990__A2 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16014_ net2348 _02224_ net1107 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[814\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_155_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13226_ _02776_ net3368 _02796_ vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__mux2_1
XFILLER_136_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10438_ _04053_ _06064_ vssd1 vssd1 vccd1 vccd1 _06065_ sky130_fd_sc_hd__nand2_1
XFILLER_6_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08396__B1 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14881__1051 clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 net2520 sky130_fd_sc_hd__inv_2
X_13157_ _02744_ _02745_ _02746_ vssd1 vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__nor3_1
X_10369_ _05886_ _05998_ net389 vssd1 vssd1 vccd1 vccd1 _05999_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_143_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12108_ net565 net362 _06638_ net178 top.CPU.registers.data\[98\] vssd1 vssd1 vccd1
+ vccd1 _06822_ sky130_fd_sc_hd__a32o_1
XFILLER_97_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13088_ top.CPU.data_out\[23\] net2847 net558 vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_23_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12039_ net145 net3455 net150 vssd1 vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__mux2_1
XFILLER_19_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_69_Left_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09360__A2 net1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12787__S net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_158_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08794__S1 net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_1_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_1_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_92_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07580_ top.CPU.registers.data\[895\] net1334 net865 top.CPU.registers.data\[863\]
+ net802 vssd1 vssd1 vccd1 vccd1 _03219_ sky130_fd_sc_hd__o221a_1
XFILLER_129_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_38_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14047__217 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 net1686 sky130_fd_sc_hd__inv_2
XANTENNA__07470__A top.CPU.control_unit.instruction\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15729_ net2063 _01939_ net1195 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[529\]
+ sky130_fd_sc_hd__dfrtp_1
X_09250_ net764 _04875_ _04887_ _04888_ vssd1 vssd1 vccd1 vccd1 _04889_ sky130_fd_sc_hd__a22o_4
XTAP_TAPCELL_ROW_66_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08201_ top.CPU.registers.data\[983\] net1295 net1014 top.CPU.registers.data\[1015\]
+ net912 vssd1 vssd1 vccd1 vccd1 _03840_ sky130_fd_sc_hd__a221o_1
X_09181_ top.CPU.registers.data\[838\] net1316 net847 top.CPU.registers.data\[870\]
+ net742 vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_32_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08132_ top.CPU.registers.data\[981\] net1299 net1020 top.CPU.registers.data\[1013\]
+ net917 vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_78_Left_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09820__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12535__B _05367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16291__Q top.CPU.data_out\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08063_ top.CPU.registers.data\[980\] net1288 net1008 top.CPU.registers.data\[1012\]
+ net905 vssd1 vssd1 vccd1 vccd1 _03702_ sky130_fd_sc_hd__a221o_1
XANTENNA__07831__C1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09179__A2 net1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10055__B _03180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13380__A0 top.CPU.control_unit.instruction\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11866__S net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12551__A top.CPU.done vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1022_A net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14745__915 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 net2384 sky130_fd_sc_hd__inv_2
XFILLER_130_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08965_ top.CPU.registers.data\[553\] top.CPU.registers.data\[521\] net805 vssd1
+ vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__mux2_1
XANTENNA__08240__S net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout482_A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08139__B1 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09336__C1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_87_Left_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07916_ top.CPU.registers.data\[572\] top.CPU.registers.data\[540\] net996 vssd1
+ vssd1 vccd1 vccd1 _03555_ sky130_fd_sc_hd__mux2_1
XFILLER_57_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08896_ _04534_ vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_162_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10502__C net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11694__B1 net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07898__C1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07847_ top.CPU.registers.data\[765\] net1379 net979 top.CPU.registers.data\[733\]
+ net906 vssd1 vssd1 vccd1 vccd1 _03486_ sky130_fd_sc_hd__a221o_1
XFILLER_112_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout270_X net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1391_A net1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout747_A net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout368_X net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13435__A1 _03200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12238__A2 _06796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07778_ top.CPU.registers.data\[542\] net997 vssd1 vssd1 vccd1 vccd1 _03417_ sky130_fd_sc_hd__and2_1
X_09517_ net1407 _03150_ _04953_ _05155_ vssd1 vssd1 vccd1 vccd1 _05156_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_140_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15796__RESET_B net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout535_X net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout914_A net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1277_X net1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09859__X _05498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10010__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09448_ top.CPU.control_unit.instruction\[9\] net1048 _04953_ _05086_ vssd1 vssd1
+ vccd1 vccd1 _05087_ sky130_fd_sc_hd__a22o_2
XANTENNA__08862__A1 net1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11901__Y _06771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_96_Left_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09379_ _05009_ _05012_ _05017_ net630 vssd1 vssd1 vccd1 vccd1 _05018_ sky130_fd_sc_hd__a22o_4
XANTENNA_fanout702_X net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11749__A1 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11410_ _06542_ net280 net269 net3466 vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__a22o_1
X_12390_ top.CPU.addressnew\[7\] top.CPU.addressnew\[13\] top.CPU.addressnew\[12\]
+ top.CPU.addressnew\[4\] vssd1 vssd1 vccd1 vccd1 _06928_ sky130_fd_sc_hd__or4bb_1
XFILLER_165_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08614__A1 _03116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11213__A3 _06648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10517__Y _06141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10421__A1 _05733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11341_ net3443 net288 net281 _06036_ vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_169_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08090__A2 net1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10972__A2 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11272_ net483 net459 _06693_ net294 net2650 vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__a32o_1
XFILLER_134_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13011_ top.SPI.paroutput\[6\] _07429_ _07431_ net3050 vssd1 vssd1 vccd1 vccd1 _01212_
+ sky130_fd_sc_hd__a22o_1
X_10223_ _03544_ _05399_ net374 vssd1 vssd1 vccd1 vccd1 _05858_ sky130_fd_sc_hd__mux2_1
XANTENNA__08917__A2 net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14191__361 clknet_leaf_179_clk vssd1 vssd1 vccd1 vccd1 net1830 sky130_fd_sc_hd__inv_2
XFILLER_161_691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14488__658 clknet_leaf_160_clk vssd1 vssd1 vccd1 vccd1 net2127 sky130_fd_sc_hd__inv_2
X_10154_ net390 _05785_ _05759_ vssd1 vssd1 vccd1 vccd1 _05791_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11077__A net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14962_ clknet_leaf_94_clk net2670 net1267 vssd1 vssd1 vccd1 vccd1 top.SPI.paroutput\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10085_ _04020_ _04093_ net378 vssd1 vssd1 vccd1 vccd1 _05723_ sky130_fd_sc_hd__mux2_1
Xhold7 top.CPU.registers.data_out_r2_prev\[13\] vssd1 vssd1 vccd1 vccd1 net2564 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09342__A2 net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11685__B1 net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14529__699 clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 net2168 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_18_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13426__A1 _02849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12229__A2 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13775_ net3 net1051 net886 net3918 vssd1 vssd1 vccd1 vccd1 _02656_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_48_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10987_ net527 _06546_ vssd1 vssd1 vccd1 vccd1 _06547_ sky130_fd_sc_hd__nor2_2
XANTENNA__08302__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12726_ _07178_ _07180_ _07176_ vssd1 vssd1 vccd1 vccd1 _07187_ sky130_fd_sc_hd__o21ai_1
X_15514_ net1848 _01724_ net1250 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[314\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_149_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16494_ clknet_leaf_41_clk _02656_ net1116 vssd1 vssd1 vccd1 vccd1 top.mmio.mem_data_i\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15445_ net1779 _01655_ net1215 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[245\]
+ sky130_fd_sc_hd__dfrtp_1
X_12657_ top.CPU.alu.program_counter\[1\] _05156_ vssd1 vssd1 vccd1 vccd1 _07125_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__12636__A top.I2C.output_state\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11608_ net132 net3226 net214 vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__mux2_1
XANTENNA__08066__C1 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15376_ net1710 _01586_ net1156 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[176\]
+ sky130_fd_sc_hd__dfrtp_1
X_12588_ top.CPU.handler.readout top.wm.curr_state\[0\] _07054_ _03131_ top.wm.curr_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00075_ sky130_fd_sc_hd__a32o_1
XANTENNA__11204__A3 _06648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11539_ net3767 net252 _06737_ net491 vssd1 vssd1 vccd1 vccd1 _01993_ sky130_fd_sc_hd__a22o_1
XANTENNA__07813__C1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10156__A net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold407 top.CPU.registers.data\[688\] vssd1 vssd1 vccd1 vccd1 net2964 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold418 top.CPU.registers.data\[352\] vssd1 vssd1 vccd1 vccd1 net2975 sky130_fd_sc_hd__dlygate4sd3_1
X_14432__602 clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 net2071 sky130_fd_sc_hd__inv_2
Xhold429 top.CPU.registers.data\[445\] vssd1 vssd1 vccd1 vccd1 net2986 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13209_ top.I2C.within_byte_counter_reading\[2\] top.I2C.within_byte_counter_reading\[0\]
+ top.I2C.within_byte_counter_reading\[1\] vssd1 vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__or3b_2
XANTENNA__09566__C1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09664__B net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08464__S0 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout909 net910 vssd1 vssd1 vccd1 vccd1 net909 sky130_fd_sc_hd__clkbuf_4
XFILLER_140_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13913__83 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 net1552 sky130_fd_sc_hd__inv_2
XANTENNA__07592__A1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08750_ _04386_ _04388_ _03342_ vssd1 vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__o21ai_1
Xhold1107 top.CPU.registers.data\[626\] vssd1 vssd1 vccd1 vccd1 net3664 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08995__S net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1118 top.CPU.registers.data\[493\] vssd1 vssd1 vccd1 vccd1 net3675 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1129 top.I2C.data_out\[24\] vssd1 vssd1 vccd1 vccd1 net3686 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_144_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12468__A2 _03783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07701_ top.CPU.control_unit.instruction\[23\] net686 vssd1 vssd1 vccd1 vccd1 _03340_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__10479__B2 top.CPU.handler.toreg\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08681_ net1285 _04318_ _04319_ vssd1 vssd1 vccd1 vccd1 _04320_ sky130_fd_sc_hd__or3_1
XANTENNA__11676__B1 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07632_ _03161_ _03254_ _03255_ _03261_ _03269_ vssd1 vssd1 vccd1 vccd1 _03271_ sky130_fd_sc_hd__a311o_2
XTAP_TAPCELL_ROW_68_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07471__Y _03111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13417__A1 net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11428__B1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07563_ top.CPU.control_unit.instruction\[19\] net873 vssd1 vssd1 vccd1 vccd1 _03202_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09302_ net918 _04940_ vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__or2_1
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11153__C net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07494_ top.mmio.s1 vssd1 vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__inv_2
XANTENNA__08844__A1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09233_ top.CPU.registers.data\[165\] net1386 net806 top.CPU.registers.data\[133\]
+ net702 vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__a221o_1
XFILLER_10_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout230_A _06772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout328_A net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09164_ top.CPU.registers.data\[454\] net1316 net848 top.CPU.registers.data\[486\]
+ net767 vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__a221o_1
XFILLER_148_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08115_ _03739_ _03753_ vssd1 vssd1 vccd1 vccd1 _03754_ sky130_fd_sc_hd__nor2_4
XANTENNA__10403__B2 top.CPU.handler.toreg\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09095_ top.CPU.registers.data\[295\] top.CPU.registers.data\[263\] net832 vssd1
+ vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__mux2_1
XFILLER_119_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10954__A2 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08046_ net1380 net1045 net899 vssd1 vssd1 vccd1 vccd1 _03685_ sky130_fd_sc_hd__o21a_2
X_14175__345 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 net1814 sky130_fd_sc_hd__inv_2
Xhold930 top.CPU.registers.data\[750\] vssd1 vssd1 vccd1 vccd1 net3487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold941 top.CPU.registers.data\[728\] vssd1 vssd1 vccd1 vccd1 net3498 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout697_A net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold952 top.CPU.registers.data\[212\] vssd1 vssd1 vccd1 vccd1 net3509 sky130_fd_sc_hd__dlygate4sd3_1
Xhold963 top.CPU.registers.data\[771\] vssd1 vssd1 vccd1 vccd1 net3520 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09021__A1 top.CPU.control_unit.instruction\[29\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_115_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_164_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10167__B1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1404_A top.CPU.control_unit.instruction\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold974 top.CPU.registers.data\[218\] vssd1 vssd1 vccd1 vccd1 net3531 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold985 top.mmio.mem_data_i\[7\] vssd1 vssd1 vccd1 vccd1 net3542 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1025_X net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09066__S net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold996 top.CPU.registers.data\[54\] vssd1 vssd1 vccd1 vccd1 net3553 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09997_ _05633_ _05635_ net383 vssd1 vssd1 vccd1 vccd1 _05636_ sky130_fd_sc_hd__mux2_1
XFILLER_103_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout485_X net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07583__A1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14216__386 clknet_leaf_126_clk vssd1 vssd1 vccd1 vccd1 net1855 sky130_fd_sc_hd__inv_2
XANTENNA_fanout864_A net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08780__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08948_ top.CPU.registers.data\[938\] top.CPU.registers.data\[906\] net971 vssd1
+ vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09324__A2 net1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08879_ top.CPU.registers.data\[331\] net1311 net842 top.CPU.registers.data\[363\]
+ net762 vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout652_X net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1394_X net1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11131__A2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10910_ _05694_ _06498_ vssd1 vssd1 vccd1 vccd1 _06500_ sky130_fd_sc_hd__nor2_2
X_11890_ _06710_ net240 net190 net3378 vssd1 vssd1 vccd1 vccd1 _01673_ sky130_fd_sc_hd__a22o_1
XANTENNA__11682__A3 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11419__B1 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10841_ net3716 net227 net319 _06449_ vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__a22o_1
XFILLER_44_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout917_X net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13560_ net3976 net578 _03002_ vssd1 vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__a21o_1
X_10772_ _05754_ _05817_ vssd1 vssd1 vccd1 vccd1 _06384_ sky130_fd_sc_hd__nor2_1
XFILLER_12_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08296__C1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14880__1050 clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 net2519 sky130_fd_sc_hd__inv_2
XFILLER_52_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12511_ _04222_ _04255_ vssd1 vssd1 vccd1 vccd1 _07020_ sky130_fd_sc_hd__or2_1
XFILLER_13_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13491_ net4027 _04918_ net588 vssd1 vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__mux2_1
XFILLER_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15230_ net1564 _01440_ net1237 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_12442_ net1054 _06957_ vssd1 vssd1 vccd1 vccd1 _00051_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_43_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08145__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11198__A2 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08599__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15161_ clknet_leaf_42_clk _01371_ net1117 vssd1 vssd1 vccd1 vccd1 top.I2C.data_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12373_ _06912_ vssd1 vssd1 vccd1 vccd1 _06913_ sky130_fd_sc_hd__inv_2
XFILLER_154_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10945__A2 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07837__X _03476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11324_ net3520 net291 net359 net148 vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__a22o_1
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15092_ net1474 _01305_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r2_prev\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07810__A2 net1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09548__C1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13287__A top.CPU.handler.readout vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07556__Y _03195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11255_ net515 _06232_ net541 vssd1 vssd1 vccd1 vccd1 _06683_ sky130_fd_sc_hd__or3_1
XFILLER_79_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10206_ net224 _05830_ _05832_ _05836_ _05841_ vssd1 vssd1 vccd1 vccd1 _05842_ sky130_fd_sc_hd__o2111a_1
XANTENNA__09563__A2 net1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11186_ net660 net141 net429 vssd1 vssd1 vccd1 vccd1 _06652_ sky130_fd_sc_hd__and3_1
XFILLER_122_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11370__A2 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13574__X _03011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08771__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10137_ _03579_ _05509_ _05513_ net371 vssd1 vssd1 vccd1 vccd1 _05774_ sky130_fd_sc_hd__a31o_1
XFILLER_39_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11238__C net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15994_ net2328 _02204_ net1250 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[794\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11658__B1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14945_ clknet_leaf_65_clk _01191_ net1166 vssd1 vssd1 vccd1 vccd1 top.CPU.alu.program_counter\[28\]
+ sky130_fd_sc_hd__dfrtp_4
X_10068_ _04891_ net373 vssd1 vssd1 vccd1 vccd1 _05706_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07877__A2 net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16615_ net1346 vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__clkbuf_1
X_13827_ net2770 net334 net327 top.CPU.data_out\[29\] vssd1 vssd1 vccd1 vccd1 _02707_
+ sky130_fd_sc_hd__a22o_1
XFILLER_51_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16546_ clknet_leaf_85_clk _02708_ net1263 vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__dfrtp_1
X_13758_ _03091_ _03089_ top.I2C.which_data_address\[0\] vssd1 vssd1 vccd1 vccd1 _02643_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12083__B1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12709_ _07166_ _07171_ net125 vssd1 vssd1 vccd1 vccd1 _07172_ sky130_fd_sc_hd__mux2_1
X_13689_ net2673 net332 vssd1 vssd1 vccd1 vccd1 _02617_ sky130_fd_sc_hd__and2_1
X_16477_ clknet_leaf_89_clk _02639_ net1274 vssd1 vssd1 vccd1 vccd1 top.SPI.timem\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12366__A top.I2C.output_state\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08039__C1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15428_ net1762 _01638_ net1212 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[228\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_129_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11189__A2 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14159__329 clknet_leaf_179_clk vssd1 vssd1 vccd1 vccd1 net1798 sky130_fd_sc_hd__inv_2
X_15359_ net1693 _01569_ net1199 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[159\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_172_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold204 top.CPU.registers.data\[907\] vssd1 vssd1 vccd1 vccd1 net2761 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold215 top.mmio.mem_data_i\[27\] vssd1 vssd1 vccd1 vccd1 net2772 sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 top.CPU.registers.data\[435\] vssd1 vssd1 vccd1 vccd1 net2783 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13335__A0 top.CPU.control_unit.instruction\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold237 top.CPU.registers.data\[444\] vssd1 vssd1 vccd1 vccd1 net2794 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12813__B _04123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13197__A top.I2C.output_state\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09920_ _05543_ _05556_ _05558_ vssd1 vssd1 vccd1 vccd1 _05559_ sky130_fd_sc_hd__a21o_1
XANTENNA__09539__C1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold248 top.CPU.registers.data\[180\] vssd1 vssd1 vccd1 vccd1 net2805 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold259 top.I2C.data_out\[30\] vssd1 vssd1 vccd1 vccd1 net2816 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12532__C _07040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout706 _03212_ vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__buf_4
XANTENNA__08211__C1 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout717 net736 vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__buf_2
X_09851_ top.CPU.registers.data\[410\] net1000 _05489_ vssd1 vssd1 vccd1 vccd1 _05490_
+ sky130_fd_sc_hd__a21o_1
Xfanout728 net735 vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__clkbuf_2
XFILLER_98_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout739 net747 vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__clkbuf_2
X_08802_ top.CPU.registers.data\[76\] net1372 net968 top.CPU.registers.data\[108\]
+ net901 vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__o221a_1
XANTENNA__11361__A2 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_142_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ net613 _05414_ _05418_ net687 top.CPU.registers.data_out_r2_prev\[27\] vssd1
+ vssd1 vccd1 vccd1 _05421_ sky130_fd_sc_hd__o32a_1
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08733_ top.CPU.registers.data\[173\] top.CPU.registers.data\[141\] net969 vssd1
+ vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__mux2_1
XANTENNA__09306__A2 net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11649__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout180_A _06777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12310__A1 _03439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11113__A2 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout278_A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08664_ top.CPU.registers.data\[174\] top.CPU.registers.data\[142\] net981 vssd1
+ vssd1 vccd1 vccd1 _04303_ sky130_fd_sc_hd__mux2_1
XANTENNA__15388__RESET_B net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10321__B1 _05687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14560__730 clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 net2199 sky130_fd_sc_hd__inv_2
XANTENNA__12861__A2 _03756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11664__A3 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07615_ net1046 _03250_ _03253_ net882 _03147_ vssd1 vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__a32o_1
XANTENNA__11164__B net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08595_ top.CPU.registers.data\[175\] top.CPU.registers.data\[143\] net975 vssd1
+ vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1187_A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07546_ top.CPU.control_unit.instruction\[11\] net662 vssd1 vssd1 vccd1 vccd1 _03185_
+ sky130_fd_sc_hd__nand2_8
XANTENNA__12074__B1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14601__771 clknet_leaf_155_clk vssd1 vssd1 vccd1 vccd1 net2240 sky130_fd_sc_hd__inv_2
XANTENNA__10624__A1 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11821__A0 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10495__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10348__X _05979_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07477_ top.CPU.alu.program_counter\[17\] vssd1 vssd1 vccd1 vccd1 _03117_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout612_A net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout233_X net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09216_ net674 _04848_ _04854_ _04842_ vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__a31o_4
XFILLER_148_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13574__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09147_ top.CPU.registers.data\[903\] net1302 net1023 top.CPU.registers.data\[935\]
+ net919 vssd1 vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__a221o_1
XANTENNA__08045__A2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout400_X net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09242__A1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_45 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09078_ top.CPU.registers.data\[520\] net1004 vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__or2_1
XANTENNA__08450__C1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout981_A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08029_ top.CPU.registers.data\[756\] net1389 net816 top.CPU.registers.data\[724\]
+ net719 vssd1 vssd1 vccd1 vccd1 _03668_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_9_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold760 top.CPU.registers.data\[420\] vssd1 vssd1 vccd1 vccd1 net3317 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1407_X net1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold771 top.CPU.registers.data\[966\] vssd1 vssd1 vccd1 vccd1 net3328 sky130_fd_sc_hd__dlygate4sd3_1
Xhold782 top.CPU.registers.data\[487\] vssd1 vssd1 vccd1 vccd1 net3339 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11888__A0 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11040_ net3653 net367 _06579_ net324 vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__a22o_1
XFILLER_150_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold793 top.CPU.registers.data\[850\] vssd1 vssd1 vccd1 vccd1 net3350 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11352__A2 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13629__A1 top.CPU.alu.program_counter\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07833__A net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12991_ _07456_ _07420_ vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__nand2b_1
Xhold1460 top.CPU.handler.toreg\[2\] vssd1 vssd1 vccd1 vccd1 net4017 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08505__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07552__B net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11942_ _06485_ net345 net229 net3029 vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__a22o_1
XFILLER_18_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_24_Left_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11873_ _05960_ net189 _06768_ vssd1 vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_28_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16400_ clknet_leaf_64_clk _00023_ net1162 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13612_ net3726 net578 _03033_ _03034_ vssd1 vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__a22o_1
X_10824_ net370 _06432_ vssd1 vssd1 vccd1 vccd1 _06433_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_28_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13801__B2 top.CPU.data_out\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16331_ clknet_leaf_66_clk _02540_ net1166 vssd1 vssd1 vccd1 vccd1 top.CPU.addressnew\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10014__C_N _03407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13543_ _03439_ net585 net339 vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__a21o_1
XFILLER_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10258__X _05892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10755_ _04923_ net508 net503 _04921_ net443 vssd1 vssd1 vccd1 vccd1 _06368_ sky130_fd_sc_hd__o221a_1
XANTENNA__09481__A1 top.CPU.registers.data_out_r1_prev\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16262_ clknet_leaf_31_clk _02472_ net1126 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.toreg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_158_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13474_ net3962 _02958_ net124 vssd1 vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__mux2_1
X_10686_ net548 _04732_ vssd1 vssd1 vccd1 vccd1 _06302_ sky130_fd_sc_hd__nor2_1
X_15213_ net1547 _01423_ net1066 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_12425_ top.I2C.I2C_state\[21\] top.I2C.reader_state\[0\] _06949_ top.I2C.initiate_read_bit
+ vssd1 vssd1 vccd1 vccd1 _00068_ sky130_fd_sc_hd__a22o_1
XFILLER_139_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16193_ net2527 _02403_ net1224 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[993\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_166_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10379__B1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11240__D net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12914__A top.CPU.alu.program_counter\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10918__A2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15144_ clknet_leaf_46_clk _01354_ net1140 vssd1 vssd1 vccd1 vccd1 top.I2C.data_out\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_138_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12356_ net1340 top.I2C.output_state\[27\] top.I2C.output_state\[3\] vssd1 vssd1
+ vccd1 vccd1 _06900_ sky130_fd_sc_hd__a21o_1
XANTENNA__11040__B2 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12633__B top.I2C.output_state\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11307_ net2941 net290 net358 net141 vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__a22o_1
X_15075_ clknet_leaf_52_clk _00053_ net1132 vssd1 vssd1 vccd1 vccd1 top.I2C.output_state\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12287_ net2583 _03682_ net1121 vssd1 vssd1 vccd1 vccd1 _01395_ sky130_fd_sc_hd__mux2_1
XFILLER_107_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11879__A0 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11238_ _06539_ net460 net526 vssd1 vssd1 vccd1 vccd1 _06674_ sky130_fd_sc_hd__and3b_1
XFILLER_150_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11343__A2 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12540__B2 _03252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15828__RESET_B net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11169_ net1402 _05809_ net429 vssd1 vssd1 vccd1 vccd1 _06646_ sky130_fd_sc_hd__and3_1
XANTENNA__07743__A net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14544__714 clknet_leaf_196_clk vssd1 vssd1 vccd1 vccd1 net2183 sky130_fd_sc_hd__inv_2
X_15977_ net2311 _02187_ net1060 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[777\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08558__B net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14928_ clknet_leaf_61_clk _01174_ net1160 vssd1 vssd1 vccd1 vccd1 top.CPU.alu.program_counter\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10303__B1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12843__A2 _03986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12795__S net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07889__S net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08380_ top.CPU.registers.data_out_r1_prev\[18\] net877 net636 _04018_ _04004_ vssd1
+ vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__o221a_4
XANTENNA__12056__B1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10606__A1 _05643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16529_ clknet_leaf_100_clk _02691_ net1255 vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11803__B1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09472__A1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_clk_X clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11431__C net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08680__C1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13556__A0 top.CPU.alu.program_counter\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09001_ top.CPU.registers.data\[937\] top.CPU.registers.data\[905\] net965 vssd1
+ vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__mux2_1
XFILLER_118_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08658__S0 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11582__A2 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12471__A_N _04019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09903_ _04922_ _04923_ vssd1 vssd1 vccd1 vccd1 _05542_ sky130_fd_sc_hd__nor2_1
Xfanout503 net505 vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_4_9_0_clk_X clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout514 net523 vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__buf_4
Xfanout525 net533 vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__clkbuf_4
XFILLER_98_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout395_A net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11874__S net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout536 net537 vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__buf_4
XANTENNA__11334__A2 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout547 _03318_ vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__clkbuf_4
X_09834_ top.CPU.registers.data\[250\] net1385 net1002 top.CPU.registers.data\[218\]
+ net922 vssd1 vssd1 vccd1 vccd1 _05473_ sky130_fd_sc_hd__a221o_1
XANTENNA__10631__X _06250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout558 net561 vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__clkbuf_4
XANTENNA__15569__RESET_B net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10998__B _03170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout569 _03176_ vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09765_ top.CPU.registers.data\[347\] net1298 net1019 top.CPU.registers.data\[379\]
+ net942 vssd1 vssd1 vccd1 vccd1 _05404_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout562_A net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14287__457 clknet_leaf_192_clk vssd1 vssd1 vccd1 vccd1 net1926 sky130_fd_sc_hd__inv_2
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout183_X net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11175__A _05693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08716_ top.CPU.registers.data\[333\] net1311 net842 top.CPU.registers.data\[365\]
+ net762 vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__a221o_1
XFILLER_39_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08499__C1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09696_ top.CPU.registers.data\[825\] top.CPU.registers.data\[793\] net1001 vssd1
+ vssd1 vccd1 vccd1 _05335_ sky130_fd_sc_hd__mux2_1
XFILLER_66_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_159_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10845__A1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08647_ top.CPU.registers.data\[462\] net1320 net851 top.CPU.registers.data\[494\]
+ net770 vssd1 vssd1 vccd1 vccd1 _04286_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_159_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout350_X net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout827_A net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14328__498 clknet_leaf_168_clk vssd1 vssd1 vccd1 vccd1 net1967 sky130_fd_sc_hd__inv_2
XFILLER_109_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08578_ top.CPU.registers.data\[303\] top.CPU.registers.data\[271\] net811 vssd1
+ vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_25_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13795__B1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07529_ _03148_ net881 vssd1 vssd1 vccd1 vccd1 _03168_ sky130_fd_sc_hd__nand2_1
XFILLER_23_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09463__A1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08266__A2 net1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout615_X net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10540_ _06111_ _06162_ net310 vssd1 vssd1 vccd1 vccd1 _06163_ sky130_fd_sc_hd__mux2_1
XANTENNA__08671__C1 net1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11270__B2 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10471_ _05733_ _05890_ _05895_ _05753_ vssd1 vssd1 vccd1 vccd1 _06097_ sky130_fd_sc_hd__a22o_1
XANTENNA__09215__A1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08018__A2 net1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_157_Right_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12734__A top.CPU.alu.program_counter\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13011__A2 _07429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12210_ _06191_ net544 _06796_ net169 top.CPU.registers.data\[46\] vssd1 vssd1 vccd1
+ vccd1 _06872_ sky130_fd_sc_hd__a32o_1
X_13190_ _02764_ _02767_ _02769_ top.I2C.sda_out top.I2C.output_state\[2\] vssd1 vssd1
+ vccd1 vccd1 _02771_ sky130_fd_sc_hd__o32a_1
XANTENNA__11022__B2 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08423__C1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout984_X net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11573__A2 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10230__C1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08974__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12141_ net2965 net173 _06838_ vssd1 vssd1 vccd1 vccd1 _01492_ sky130_fd_sc_hd__a21o_1
XFILLER_68_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11069__B net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12072_ _06615_ net348 net178 net3296 vssd1 vssd1 vccd1 vccd1 _01527_ sky130_fd_sc_hd__a22o_1
X_14231__401 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 net1870 sky130_fd_sc_hd__inv_2
XFILLER_89_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold590 top.CPU.registers.data\[666\] vssd1 vssd1 vccd1 vccd1 net3147 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11325__A2 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11023_ net518 _06429_ net543 vssd1 vssd1 vccd1 vccd1 _06569_ sky130_fd_sc_hd__and3_1
X_15900_ net2234 _02110_ net1235 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[700\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10533__B1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09254__S net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07563__A top.CPU.control_unit.instruction\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15831_ net2165 _02041_ net1182 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[631\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_66_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_32_Left_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12974_ top.I2C.bit_timer_counter\[3\] _07407_ vssd1 vssd1 vccd1 vccd1 _07409_ sky130_fd_sc_hd__and2_1
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15762_ net2096 _01972_ net1102 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[562\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1290 top.CPU.registers.data\[332\] vssd1 vssd1 vccd1 vccd1 net3847 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10836__A1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11925_ net3302 net186 net350 _06336_ vssd1 vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__a22o_1
XFILLER_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15693_ net2027 _01903_ net1057 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[493\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_75_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12038__A0 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11856_ _06692_ net206 net155 net2652 vssd1 vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__a22o_1
XFILLER_159_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12589__A1 top.CPU.handler.readout vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13786__B1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10807_ net386 _06343_ _06415_ _06416_ net400 vssd1 vssd1 vccd1 vccd1 _06417_ sky130_fd_sc_hd__o221a_1
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11787_ net459 _06633_ net235 net161 net3276 vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__a32o_1
XANTENNA__10429__A net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16314_ clknet_leaf_84_clk _02523_ net1263 vssd1 vssd1 vccd1 vccd1 top.CPU.data_out\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13526_ top.CPU.data_out\[21\] net589 net339 _02983_ vssd1 vssd1 vccd1 vccd1 _02519_
+ sky130_fd_sc_hd__o22a_1
X_10738_ _06350_ _06351_ _06338_ _06349_ vssd1 vssd1 vccd1 vccd1 _06352_ sky130_fd_sc_hd__o211ai_4
XANTENNA__12576__D_N _07080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_41_Left_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13538__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13457_ net1399 net872 _02900_ net419 vssd1 vssd1 vccd1 vccd1 _02950_ sky130_fd_sc_hd__a31o_1
X_16245_ clknet_leaf_43_clk _02455_ net1117 vssd1 vssd1 vccd1 vccd1 top.CPU.control_unit.instruction\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10669_ _05279_ _05531_ _05564_ _05565_ net444 vssd1 vssd1 vccd1 vccd1 _06286_ sky130_fd_sc_hd__a221o_1
XFILLER_9_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_124_Right_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12408_ top.CPU.addressnew\[9\] top.CPU.addressnew\[10\] top.CPU.addressnew\[11\]
+ top.CPU.addressnew\[8\] vssd1 vssd1 vccd1 vccd1 _06934_ sky130_fd_sc_hd__or4bb_1
XTAP_TAPCELL_ROW_11_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09429__S net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12210__B1 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13388_ top.I2C.data_out\[22\] net555 _02859_ top.mmio.mem_data_i\[22\] vssd1 vssd1
+ vccd1 vccd1 _02909_ sky130_fd_sc_hd__a22o_1
X_16176_ net2510 _02386_ net1154 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[976\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 gpio_oeb[1] sky130_fd_sc_hd__buf_2
XFILLER_142_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07768__A1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput117 net117 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__buf_2
XANTENNA__11564__A2 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15127_ clknet_leaf_57_clk _01337_ net1146 vssd1 vssd1 vccd1 vccd1 top.I2C.within_byte_counter_writing\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_58_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12339_ net2585 _05154_ net1252 vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__mux2_1
XFILLER_49_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15058_ clknet_leaf_52_clk _00062_ net1132 vssd1 vssd1 vccd1 vccd1 top.I2C.output_state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09509__A2 net1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11316__A2 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07880_ top.CPU.registers.data\[604\] net1332 net863 top.CPU.registers.data\[636\]
+ net754 vssd1 vssd1 vccd1 vccd1 _03519_ sky130_fd_sc_hd__a221o_1
XANTENNA__10524__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_50_Left_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09017__X _04656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10611__B _06230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09550_ net711 _05178_ _05181_ _05187_ _05188_ vssd1 vssd1 vccd1 vccd1 _05189_ sky130_fd_sc_hd__o32a_2
X_14015__185 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 net1654 sky130_fd_sc_hd__inv_2
X_08501_ _04136_ _04139_ net639 vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__a21o_1
XANTENNA__10827__A1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09481_ top.CPU.registers.data_out_r1_prev\[2\] net875 _05105_ _05119_ vssd1 vssd1
+ vccd1 vccd1 _05120_ sky130_fd_sc_hd__o211ai_4
XANTENNA__09693__A1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08432_ net709 _04069_ _04070_ vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__or3_1
XANTENNA__10984__D net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08363_ _04000_ _04001_ net692 vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__a21o_1
XFILLER_23_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout143_A _06173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16450__RESET_B net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11252__A1 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11161__C net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08294_ top.CPU.registers.data\[467\] net1326 net857 top.CPU.registers.data\[499\]
+ net774 vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__a221o_1
X_14672__842 clknet_leaf_196_clk vssd1 vssd1 vccd1 vccd1 net2311 sky130_fd_sc_hd__inv_2
XANTENNA__11869__S net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout408_A _05023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13002__X _07429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09748__A2 net1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12201__B1 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08405__C1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14713__883 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 net2352 sky130_fd_sc_hd__inv_2
XANTENNA__11555__A2 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10763__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12487__A1_N _04566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1317_A net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout300 _06645_ vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__clkbuf_4
Xfanout311 net315 vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__buf_4
XANTENNA_fanout398_X net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1309 net1323 vssd1 vssd1 vccd1 vccd1 net1309 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout777_A net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11307__A2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout322 _03195_ vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__clkbuf_4
Xfanout333 net334 vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__buf_2
XANTENNA__10802__A net1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout344 net346 vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__buf_4
XFILLER_98_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08184__A1 top.CPU.control_unit.instruction\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout355 net356 vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1105_X net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout366 net369 vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__clkbuf_8
XFILLER_47_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout377 net380 vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__buf_2
X_09817_ net710 _05452_ _05453_ net642 vssd1 vssd1 vccd1 vccd1 _05456_ sky130_fd_sc_hd__a31o_1
Xfanout388 net393 vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__clkbuf_2
XFILLER_98_1006 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout399 net400 vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__buf_2
XANTENNA_fanout565_X net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout944_A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13874__44 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 net1513 sky130_fd_sc_hd__inv_2
X_09748_ top.CPU.registers.data\[859\] net1328 net862 top.CPU.registers.data\[891\]
+ net777 vssd1 vssd1 vccd1 vccd1 _05387_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout732_X net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09679_ top.CPU.registers.data\[857\] net1336 net869 top.CPU.registers.data\[889\]
+ net757 vssd1 vssd1 vccd1 vccd1 _05318_ sky130_fd_sc_hd__a221o_1
XANTENNA__11055__D net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11710_ _06545_ net206 net420 net3196 vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__a22o_1
XANTENNA__11491__A1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _07154_ _07151_ net125 vssd1 vssd1 vccd1 vccd1 _07155_ sky130_fd_sc_hd__mux2_1
X_11641_ _06058_ net201 net425 net3699 vssd1 vssd1 vccd1 vccd1 _01910_ sky130_fd_sc_hd__a22o_1
XANTENNA__08239__A2 net1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11572_ net570 _06683_ vssd1 vssd1 vccd1 vccd1 _06744_ sky130_fd_sc_hd__nor2_1
XANTENNA__11243__B2 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13311_ top.CPU.control_unit.instruction\[1\] _02852_ net667 vssd1 vssd1 vccd1 vccd1
+ _02435_ sky130_fd_sc_hd__mux2_1
Xinput19 DAT_I[25] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__buf_1
XFILLER_168_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10523_ net511 _06060_ _06130_ _06146_ _06129_ vssd1 vssd1 vccd1 vccd1 _06147_ sky130_fd_sc_hd__a311o_2
X_13242_ _02803_ _02804_ _02805_ net3614 vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__a22o_1
XFILLER_109_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16030_ net2364 _02240_ net1237 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[830\]
+ sky130_fd_sc_hd__dfrtp_1
X_10454_ net224 _06080_ _06078_ _06073_ vssd1 vssd1 vccd1 vccd1 _06081_ sky130_fd_sc_hd__o211a_2
XANTENNA__09739__A2 net1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08153__S net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08006__X _03645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12183__B net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11546__A2 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13173_ top.I2C.byte_manager_state\[2\] top.I2C.output_state\[14\] _06916_ vssd1
+ vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__and3_1
X_10385_ _05752_ _05778_ vssd1 vssd1 vccd1 vccd1 _06014_ sky130_fd_sc_hd__or2_1
XFILLER_123_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_107_Left_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12124_ top.CPU.registers.data\[90\] net655 _06749_ vssd1 vssd1 vccd1 vccd1 _06830_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_92_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10134__D net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12055_ net567 _06606_ net242 net179 net3184 vssd1 vssd1 vccd1 vccd1 _01536_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_53_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_53_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11849__A3 net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09372__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11006_ net2987 net216 _06558_ net311 vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__a22o_1
X_15814_ net2148 _02024_ net1075 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[614\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09712__S net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10809__A1 _05672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10809__B2 _05665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15745_ net2079 _01955_ net1250 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[545\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_92_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12957_ _07394_ _07395_ vssd1 vssd1 vccd1 vccd1 _07396_ sky130_fd_sc_hd__nor2_1
XANTENNA__13471__A2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_116_Left_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11482__A1 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11908_ net3564 net184 net346 _05963_ vssd1 vssd1 vccd1 vccd1 _01658_ sky130_fd_sc_hd__a22o_1
XANTENNA__08883__C1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15676_ net2010 _01886_ net1194 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[476\]
+ sky130_fd_sc_hd__dfrtp_1
X_12888_ top.CPU.alu.program_counter\[24\] _07322_ vssd1 vssd1 vccd1 vccd1 _07334_
+ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_16_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09427__A1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11839_ _06670_ net200 net153 net2843 vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__a22o_1
X_14656__826 clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 net2295 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_99_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07989__A1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11785__A2 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13509_ top.CPU.data_out\[13\] net587 _02969_ _02974_ vssd1 vssd1 vccd1 vccd1 _02511_
+ sky130_fd_sc_hd__o22a_1
X_14400__570 clknet_leaf_112_clk vssd1 vssd1 vccd1 vccd1 net2039 sky130_fd_sc_hd__inv_2
XANTENNA__12374__A top.I2C.output_state\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16228_ clknet_leaf_29_clk _02438_ net1151 vssd1 vssd1 vccd1 vccd1 top.CPU.control_unit.instruction\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_127_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09286__S0 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11537__A2 _06311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16159_ net2493 _02369_ net1219 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[959\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07618__D net1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08981_ top.CPU.registers.data\[457\] net1309 net840 top.CPU.registers.data\[489\]
+ net761 vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__a221o_1
XANTENNA__13409__S net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07932_ top.CPU.registers.data\[476\] net1303 net1023 top.CPU.registers.data\[508\]
+ net920 vssd1 vssd1 vccd1 vccd1 _03571_ sky130_fd_sc_hd__a221o_1
XANTENNA__16289__Q top.CPU.data_out\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07863_ top.CPU.registers.data\[285\] net980 _03501_ vssd1 vssd1 vccd1 vccd1 _03502_
+ sky130_fd_sc_hd__a21o_1
XFILLER_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10979__D net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07913__A1 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09602_ top.CPU.registers.data\[224\] net1387 net810 top.CPU.registers.data\[192\]
+ net765 vssd1 vssd1 vccd1 vccd1 _05241_ sky130_fd_sc_hd__a221o_1
XFILLER_113_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07794_ top.CPU.registers.data\[94\] net1303 net1025 top.CPU.registers.data\[126\]
+ net944 vssd1 vssd1 vccd1 vccd1 _03433_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_108_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09533_ net803 _05170_ _05171_ net732 vssd1 vssd1 vccd1 vccd1 _05172_ sky130_fd_sc_hd__o211a_1
XFILLER_71_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10768__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout260_A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout358_A net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12670__A0 top.CPU.alu.program_counter\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09464_ net795 _05097_ _05098_ net748 vssd1 vssd1 vccd1 vccd1 _05103_ sky130_fd_sc_hd__o211a_1
XANTENNA__08874__C1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08238__S net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08415_ _03989_ _04053_ vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__nand2_1
X_09395_ net797 _05029_ _05030_ net751 vssd1 vssd1 vccd1 vccd1 _05034_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout525_A net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14399__569 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 net2038 sky130_fd_sc_hd__inv_2
XANTENNA_fanout146_X net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1267_A net1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08346_ net899 _03159_ vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__nand2b_2
XANTENNA__11225__A1 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09858__A net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08626__C1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11776__A2 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11599__S net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08277_ net1365 net1045 net899 vssd1 vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__o21a_2
XFILLER_20_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08641__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout313_X net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10516__B _06139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout894_A net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11528__A2 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10008__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09051__C1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10170_ top.CPU.fetch.current_ra\[29\] net1043 net882 top.CPU.handler.toreg\[29\]
+ vssd1 vssd1 vccd1 vccd1 _05807_ sky130_fd_sc_hd__a22o_1
XFILLER_121_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_167_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12731__B top.CPU.alu.program_counter\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout682_X net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13319__S net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11628__A net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1106 net1108 vssd1 vssd1 vccd1 vccd1 net1106 sky130_fd_sc_hd__clkbuf_4
XFILLER_154_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1117 net1118 vssd1 vssd1 vccd1 vccd1 net1117 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12489__B1 _04633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout130 _06464_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__buf_2
Xfanout1128 net1136 vssd1 vssd1 vccd1 vccd1 net1128 sky130_fd_sc_hd__clkbuf_4
Xfanout1139 net1140 vssd1 vssd1 vccd1 vccd1 net1139 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13150__A1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout141 _06105_ vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__buf_2
XANTENNA__09354__B1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout152 net153 vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__buf_4
XANTENNA__13150__B2 top.CPU.alu.program_counter\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout163 _06760_ vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__clkbuf_4
Xfanout174 _06825_ vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__buf_4
XFILLER_87_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout185 net187 vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout947_X net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11700__A2 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout196 net197 vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__buf_4
X_12811_ top.CPU.alu.program_counter\[17\] _04123_ vssd1 vssd1 vccd1 vccd1 _07264_
+ sky130_fd_sc_hd__nor2_1
X_13791_ net20 net1052 net887 net3875 vssd1 vssd1 vccd1 vccd1 _02672_ sky130_fd_sc_hd__a22o_1
XFILLER_170_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13453__A2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14343__513 clknet_leaf_185_clk vssd1 vssd1 vccd1 vccd1 net1982 sky130_fd_sc_hd__inv_2
XANTENNA__11363__A net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07560__B _03154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12661__A0 _03100_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15530_ net1864 _01740_ net1088 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[330\]
+ sky130_fd_sc_hd__dfrtp_1
X_12742_ net1379 net1363 _03159_ vssd1 vssd1 vccd1 vccd1 _07201_ sky130_fd_sc_hd__mux2_1
XANTENNA__08865__C1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12178__B net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12673_ _07137_ _07138_ vssd1 vssd1 vccd1 vccd1 _07139_ sky130_fd_sc_hd__and2_1
X_15461_ net1795 _01671_ net1063 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[261\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09409__A1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_190_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_190_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_13_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11624_ net148 net3220 net214 vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__mux2_1
XFILLER_8_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15392_ net1726 _01602_ net1092 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[192\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07559__Y _03198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11555_ _06668_ net262 net248 net2995 vssd1 vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__a22o_1
XANTENNA__09290__C1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08632__A2 net1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10506_ _04193_ _05575_ vssd1 vssd1 vccd1 vccd1 _06130_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_94_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11486_ net484 net473 _06616_ net255 net3340 vssd1 vssd1 vccd1 vccd1 _02038_ sky130_fd_sc_hd__a32o_1
XFILLER_155_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11519__A2 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13225_ _02780_ _02792_ vssd1 vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__nand2_1
XFILLER_137_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16013_ net2347 _02223_ net1076 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[813\]
+ sky130_fd_sc_hd__dfrtp_1
X_10437_ net370 _05964_ vssd1 vssd1 vccd1 vccd1 _06064_ sky130_fd_sc_hd__nor2_1
XFILLER_170_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10727__B1 _06139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12192__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13156_ top.I2C.output_state\[6\] top.I2C.output_state\[22\] top.I2C.output_state\[19\]
+ top.I2C.output_state\[23\] vssd1 vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__or4_1
X_10368_ _05941_ _05997_ net310 vssd1 vssd1 vccd1 vccd1 _05998_ sky130_fd_sc_hd__mux2_1
XFILLER_98_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12107_ net3961 net178 _06821_ _06730_ vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__a22o_1
XFILLER_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13087_ top.CPU.data_out\[22\] net3243 net559 vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__mux2_1
X_10299_ top.CPU.fetch.current_ra\[25\] net1043 net882 top.CPU.handler.toreg\[25\]
+ vssd1 vssd1 vccd1 vccd1 _05932_ sky130_fd_sc_hd__a22o_1
XFILLER_111_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09790__X _05429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13141__A1 top.CPU.data_out\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12038_ net142 net3150 net150 vssd1 vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__mux2_1
XANTENNA__08699__A2 net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13951__121 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 net1590 sky130_fd_sc_hd__inv_2
XANTENNA__11152__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11273__A net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14086__256 clknet_leaf_122_clk vssd1 vssd1 vccd1 vccd1 net1725 sky130_fd_sc_hd__inv_2
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15728_ net2062 _01938_ net1156 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[528\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08320__A1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_103_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15659_ net1993 _01869_ net1059 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[459\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08871__A2 net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_181_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_181_clk
+ sky130_fd_sc_hd__clkbuf_8
X_08200_ top.CPU.registers.data\[855\] net1295 net1014 top.CPU.registers.data\[887\]
+ net937 vssd1 vssd1 vccd1 vccd1 _03839_ sky130_fd_sc_hd__a221o_1
XANTENNA__11207__B2 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14127__297 clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 net1766 sky130_fd_sc_hd__inv_2
X_09180_ top.CPU.registers.data\[742\] net1386 net814 top.CPU.registers.data\[710\]
+ net718 vssd1 vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_32_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11758__A2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08131_ net957 _03763_ _03769_ vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__and3_1
XANTENNA__07469__Y _03109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08623__A2 net1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08062_ top.CPU.registers.data\[852\] net1288 net1008 top.CPU.registers.data\[884\]
+ net931 vssd1 vssd1 vccd1 vccd1 _03701_ sky130_fd_sc_hd__a221o_1
XFILLER_128_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09033__C1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10718__B1 _06332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08387__A1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08521__S net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11391__B1 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13139__S _07418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14784__954 clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 net2423 sky130_fd_sc_hd__inv_2
XFILLER_170_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11930__A2 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08964_ _04600_ _04602_ vssd1 vssd1 vccd1 vccd1 _04603_ sky130_fd_sc_hd__or2_2
XANTENNA_fanout1015_A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09336__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07915_ top.CPU.registers.data\[604\] net1302 net1023 top.CPU.registers.data\[636\]
+ net943 vssd1 vssd1 vccd1 vccd1 _03554_ sky130_fd_sc_hd__a221o_1
X_08895_ _04501_ _04532_ vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__and2_1
XFILLER_130_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_162_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11882__S net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout475_A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14030__200 clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 net1669 sky130_fd_sc_hd__inv_2
XANTENNA__10502__D net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14825__995 clknet_leaf_155_clk vssd1 vssd1 vccd1 vccd1 net2464 sky130_fd_sc_hd__inv_2
XFILLER_29_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07846_ net952 _03479_ _03481_ _03484_ vssd1 vssd1 vccd1 vccd1 _03485_ sky130_fd_sc_hd__a31o_1
XANTENNA__12891__B1 top.CPU.alu.program_counter\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13844__14 clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 net1483 sky130_fd_sc_hd__inv_2
X_07777_ _03411_ _03415_ vssd1 vssd1 vccd1 vccd1 _03416_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_123_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout263_X net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout642_A net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1384_A net1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09516_ net1041 net1039 net1285 vssd1 vssd1 vccd1 vccd1 _05155_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_140_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09447_ net1365 _04595_ vssd1 vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__or2_1
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11997__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout430_X net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_172_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_172_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_12_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout528_X net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout907_A net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09588__A _05226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09378_ net607 _05013_ _05014_ _05015_ _05016_ vssd1 vssd1 vccd1 vccd1 _05017_ sky130_fd_sc_hd__o32a_1
XFILLER_40_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11749__A2 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08329_ top.CPU.registers.data\[179\] net1383 net988 top.CPU.registers.data\[147\]
+ net678 vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__a221o_1
XFILLER_165_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08075__B1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09811__A1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10527__A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11340_ net3469 net288 net282 _06011_ vssd1 vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_169_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11271_ net515 _06562_ vssd1 vssd1 vccd1 vccd1 _06693_ sky130_fd_sc_hd__nor2_1
XFILLER_134_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13010_ top.SPI.paroutput\[5\] _07429_ _07431_ net3221 vssd1 vssd1 vccd1 vccd1 _01211_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08378__A1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10222_ _05429_ net507 _05680_ _05433_ _05856_ vssd1 vssd1 vccd1 vccd1 _05857_ sky130_fd_sc_hd__a221o_1
XFILLER_152_158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12174__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07836__A _03474_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11629__Y _06756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12461__B _05498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11382__B1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11921__A2 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10153_ _05788_ _05789_ net389 vssd1 vssd1 vccd1 vccd1 _05790_ sky130_fd_sc_hd__mux2_1
X_13935__105 clknet_leaf_192_clk vssd1 vssd1 vccd1 vccd1 net1574 sky130_fd_sc_hd__inv_2
XFILLER_0_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11077__B _06373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input36_A gpio_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14961_ clknet_leaf_93_clk net2719 net1268 vssd1 vssd1 vccd1 vccd1 top.SPI.paroutput\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10084_ _05711_ _05721_ net399 vssd1 vssd1 vccd1 vccd1 _05722_ sky130_fd_sc_hd__mux2_1
Xhold8 top.I2C.I2C_state\[18\] vssd1 vssd1 vccd1 vccd1 net2565 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13573__A top.CPU.alu.program_counter\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11685__A1 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08550__A1 top.CPU.control_unit.instruction\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11093__A net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11437__B2 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13774_ net33 net1049 net884 net3747 vssd1 vssd1 vccd1 vccd1 _02655_ sky130_fd_sc_hd__o22a_1
XANTENNA__08954__X _04593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10986_ net1405 _03170_ net146 vssd1 vssd1 vccd1 vccd1 _06546_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_48_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15513_ net1847 _01723_ net1244 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[313\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11988__A2 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12725_ _07183_ _07184_ vssd1 vssd1 vccd1 vccd1 _07186_ sky130_fd_sc_hd__nand2_1
X_16493_ clknet_leaf_41_clk _02655_ net1115 vssd1 vssd1 vccd1 vccd1 top.mmio.mem_data_i\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_163_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_163_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08853__A2 net1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15444_ net1778 _01654_ net1073 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[244\]
+ sky130_fd_sc_hd__dfrtp_1
X_12656_ top.CPU.alu.program_counter\[1\] _05156_ vssd1 vssd1 vccd1 vccd1 _07124_
+ sky130_fd_sc_hd__nand2_1
X_11607_ _06056_ net3216 net213 vssd1 vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__mux2_1
X_12587_ net3841 _03131_ top.wm.curr_state\[0\] _07090_ vssd1 vssd1 vccd1 vccd1 _00076_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09263__C1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15375_ net1709 _01585_ net1088 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[175\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10437__A net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07813__B1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11538_ _03182_ net474 _06510_ vssd1 vssd1 vccd1 vccd1 _06737_ sky130_fd_sc_hd__and3_1
XFILLER_144_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14471__641 clknet_leaf_187_clk vssd1 vssd1 vccd1 vccd1 net2110 sky130_fd_sc_hd__inv_2
Xhold408 top.CPU.registers.data\[82\] vssd1 vssd1 vccd1 vccd1 net2965 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold419 top.CPU.registers.data\[368\] vssd1 vssd1 vccd1 vccd1 net2976 sky130_fd_sc_hd__dlygate4sd3_1
X_11469_ net148 net3297 net265 vssd1 vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__mux2_1
XFILLER_7_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14768__938 clknet_leaf_198_clk vssd1 vssd1 vccd1 vccd1 net2407 sky130_fd_sc_hd__inv_2
XANTENNA__09566__B1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12165__A2 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13208_ net3760 _02779_ _02784_ _02773_ vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__a22o_1
XFILLER_48_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09030__A2 net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11373__B1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08464__S1 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07577__C1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11912__A2 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13139_ top.SPI.command\[1\] top.CPU.data_out\[1\] _07418_ vssd1 vssd1 vccd1 vccd1
+ _01290_ sky130_fd_sc_hd__mux2_1
X_14512__682 clknet_leaf_199_clk vssd1 vssd1 vccd1 vccd1 net2151 sky130_fd_sc_hd__inv_2
XFILLER_31_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10172__A net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09318__A0 _04951_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14809__979 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 net2448 sky130_fd_sc_hd__inv_2
Xhold1108 top.CPU.registers.data\[645\] vssd1 vssd1 vccd1 vccd1 net3665 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1119 top.CPU.registers.data\[1022\] vssd1 vssd1 vccd1 vccd1 net3676 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11125__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07700_ _03116_ _03331_ vssd1 vssd1 vccd1 vccd1 _03339_ sky130_fd_sc_hd__nor2_1
XFILLER_66_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08680_ top.CPU.registers.data\[590\] net1378 net981 top.CPU.registers.data\[622\]
+ net908 vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__o221a_1
XANTENNA__11676__A1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07631_ _03161_ _03254_ _03255_ _03261_ _03269_ vssd1 vssd1 vccd1 vccd1 _03270_ sky130_fd_sc_hd__a311oi_4
XTAP_TAPCELL_ROW_68_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07562_ net1048 _03164_ net1039 vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__or3_1
XFILLER_0_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09301_ top.CPU.registers.data\[676\] top.CPU.registers.data\[644\] net992 vssd1
+ vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__mux2_1
XANTENNA__11979__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07493_ top.SPI.busy vssd1 vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_154_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_154_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_22_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08583__Y _04222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09232_ _04869_ _04870_ net640 vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__a21o_1
XFILLER_167_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10651__A2 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09163_ top.CPU.registers.data\[422\] top.CPU.registers.data\[390\] net814 vssd1
+ vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__mux2_1
XFILLER_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12038__S net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10347__A net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout223_A _06469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08114_ net643 _03749_ _03752_ net709 _03746_ vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__o311a_1
X_09094_ top.CPU.alu.program_counter\[7\] net1034 vssd1 vssd1 vccd1 vccd1 _04733_
+ sky130_fd_sc_hd__nor2_1
XFILLER_163_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11877__S net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08045_ net880 net451 _03651_ vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__o21ai_2
XANTENNA__09006__C1 _03342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10634__X _06253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold920 top.CPU.registers.data\[132\] vssd1 vssd1 vccd1 vccd1 net3477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold931 top.CPU.registers.data\[497\] vssd1 vssd1 vccd1 vccd1 net3488 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12156__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold942 top.CPU.registers.data\[796\] vssd1 vssd1 vccd1 vccd1 net3499 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08251__S net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold953 top.CPU.registers.data\[799\] vssd1 vssd1 vccd1 vccd1 net3510 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold964 top.CPU.registers.data\[859\] vssd1 vssd1 vccd1 vccd1 net3521 sky130_fd_sc_hd__dlygate4sd3_1
Xhold975 top.CPU.data_out\[7\] vssd1 vssd1 vccd1 vccd1 net3532 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_164_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold986 top.I2C.output_state\[17\] vssd1 vssd1 vccd1 vccd1 net3543 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_164_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11903__A2 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold997 top.CPU.registers.data\[1010\] vssd1 vssd1 vccd1 vccd1 net3554 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09996_ _04634_ net377 _05634_ vssd1 vssd1 vccd1 vccd1 _05635_ sky130_fd_sc_hd__o21ba_1
XFILLER_89_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1018_X net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09309__B1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09871__A _03476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout380_X net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08947_ net626 _04582_ _04585_ vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__or3_1
XFILLER_28_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout478_X net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout857_A net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_84_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_13 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08878_ top.CPU.registers.data\[299\] top.CPU.registers.data\[267\] net807 vssd1
+ vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__mux2_1
XFILLER_85_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07829_ net791 _03463_ _03464_ net743 vssd1 vssd1 vccd1 vccd1 _03468_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout645_X net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1387_X net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10840_ net531 _06448_ vssd1 vssd1 vccd1 vccd1 _06449_ sky130_fd_sc_hd__nor2_1
XANTENNA__09088__A2 _04726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10627__C1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_99_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10771_ _06382_ _06051_ net416 _06381_ vssd1 vssd1 vccd1 vccd1 _06383_ sky130_fd_sc_hd__o2bb2a_1
Xclkbuf_leaf_145_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_145_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_44_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout812_X net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12510_ _04291_ _04324_ _04362_ _04391_ vssd1 vssd1 vccd1 vccd1 _07019_ sky130_fd_sc_hd__o22a_1
XANTENNA_clkbuf_leaf_142_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13490_ top.CPU.data_out\[4\] _04951_ net587 vssd1 vssd1 vccd1 vccd1 _02502_ sky130_fd_sc_hd__mux2_1
XFILLER_13_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08426__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12441_ net1341 top.I2C.output_state\[4\] top.I2C.output_state\[19\] vssd1 vssd1
+ vccd1 vccd1 _06957_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_22_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09245__C1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14455__625 clknet_leaf_76_clk vssd1 vssd1 vccd1 vccd1 net2094 sky130_fd_sc_hd__inv_2
X_12372_ _03124_ _06911_ vssd1 vssd1 vccd1 vccd1 _06912_ sky130_fd_sc_hd__nor2_1
X_15160_ clknet_leaf_42_clk _01370_ net1117 vssd1 vssd1 vccd1 vccd1 top.I2C.data_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_166_784 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09260__A2 net1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_157_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11323_ net3004 net291 net359 net147 vssd1 vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__a22o_1
XFILLER_125_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15091_ net1473 _01304_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r2_prev\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_4_0_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_0_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_5_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12472__A _03955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12147__A2 _06749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11254_ net2904 net293 _06682_ net311 vssd1 vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_37_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13287__B _03126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11355__B1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10205_ _05741_ _05828_ _05840_ _05733_ vssd1 vssd1 vccd1 vccd1 _05841_ sky130_fd_sc_hd__a22oi_1
XFILLER_140_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11185_ net1402 net488 _06651_ net299 net2888 vssd1 vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__a32o_1
XANTENNA__08771__A1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10136_ _03579_ _05509_ _05513_ vssd1 vssd1 vccd1 vccd1 _05773_ sky130_fd_sc_hd__a21oi_1
XFILLER_67_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11107__B1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15993_ net2327 _02203_ net1244 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[793\]
+ sky130_fd_sc_hd__dfrtp_1
X_14944_ clknet_leaf_66_clk _01190_ net1165 vssd1 vssd1 vccd1 vccd1 top.CPU.alu.program_counter\[27\]
+ sky130_fd_sc_hd__dfrtp_4
X_10067_ _04829_ net377 vssd1 vssd1 vccd1 vccd1 _05705_ sky130_fd_sc_hd__nor2_1
XFILLER_48_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10720__A net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09720__B1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload1_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16614_ net1346 vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_1
XFILLER_47_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13826_ net88 net338 net329 net3772 vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__a22o_1
XFILLER_62_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09079__A2 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16545_ clknet_leaf_99_clk _02707_ net1256 vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__dfrtp_1
X_13757_ _03089_ _03090_ vssd1 vssd1 vccd1 vccd1 _03091_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_136_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_136_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_100_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10969_ net518 net440 net133 net546 vssd1 vssd1 vccd1 vccd1 _06536_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_63_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11551__A net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12708_ _07169_ _07170_ vssd1 vssd1 vccd1 vccd1 _07171_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16476_ clknet_leaf_88_clk _02638_ net1274 vssd1 vssd1 vccd1 vccd1 top.SPI.timem\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08336__S net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13688_ net2706 net336 vssd1 vssd1 vccd1 vccd1 _02616_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_80_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15427_ net1761 _01637_ net1207 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[227\]
+ sky130_fd_sc_hd__dfrtp_1
X_12639_ top.I2C.output_state\[26\] net2632 vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__and2_1
XFILLER_79_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09956__A _03650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14198__368 clknet_leaf_180_clk vssd1 vssd1 vccd1 vccd1 net1837 sky130_fd_sc_hd__inv_2
XFILLER_156_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15358_ net1692 _01568_ net1239 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[158\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_145_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold205 top.SPI.paroutput\[9\] vssd1 vssd1 vccd1 vccd1 net2762 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10454__X _06081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12382__A top.CPU.handler.readout vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15289_ net1623 _01499_ net1223 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[89\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold216 top.CPU.registers.data\[568\] vssd1 vssd1 vccd1 vccd1 net2773 sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 top.CPU.registers.data\[170\] vssd1 vssd1 vccd1 vccd1 net2784 sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 net39 vssd1 vssd1 vccd1 vccd1 net2795 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12138__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09167__S net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07476__A top.CPU.control_unit.instruction\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold249 top.CPU.registers.data\[895\] vssd1 vssd1 vccd1 vccd1 net2806 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11346__B1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09962__Y _05601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09850_ top.CPU.registers.data\[442\] net1027 net921 vssd1 vssd1 vccd1 vccd1 _05489_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__08211__B1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout707 net709 vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__buf_4
Xfanout718 net722 vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__clkbuf_4
Xfanout729 net734 vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08762__A1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08801_ _04438_ _04439_ net935 vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__mux2_1
XANTENNA__16404__RESET_B net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09781_ net956 _05411_ _05410_ net939 vssd1 vssd1 vccd1 vccd1 _05420_ sky130_fd_sc_hd__o211a_1
XFILLER_58_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08732_ top.CPU.registers.data\[45\] top.CPU.registers.data\[13\] net969 vssd1 vssd1
+ vccd1 vccd1 _04371_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08514__A1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16297__Q top.CPU.data_out\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08663_ top.CPU.registers.data\[46\] top.CPU.registers.data\[14\] net981 vssd1 vssd1
+ vccd1 vccd1 _04302_ sky130_fd_sc_hd__mux2_1
XFILLER_82_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10321__A1 _05643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout173_A _06825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07614_ top.CPU.control_unit.instruction\[14\] _03252_ vssd1 vssd1 vccd1 vccd1 _03253_
+ sky130_fd_sc_hd__nand2_1
XFILLER_81_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08594_ top.CPU.registers.data\[47\] top.CPU.registers.data\[15\] net975 vssd1 vssd1
+ vccd1 vccd1 _04233_ sky130_fd_sc_hd__mux2_1
XFILLER_54_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08278__A0 _03915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07545_ net563 _03183_ vssd1 vssd1 vccd1 vccd1 _03184_ sky130_fd_sc_hd__nand2_2
XANTENNA__12074__A1 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_138_Right_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_127_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_127_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09475__C1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10085__A0 _04020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_5_0_clk_X clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1082_A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout438_A net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14142__312 clknet_leaf_152_clk vssd1 vssd1 vccd1 vccd1 net1781 sky130_fd_sc_hd__inv_2
X_07476_ top.CPU.control_unit.instruction\[23\] vssd1 vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_157_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08246__S net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14439__609 clknet_leaf_183_clk vssd1 vssd1 vccd1 vccd1 net2078 sky130_fd_sc_hd__inv_2
XFILLER_167_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09215_ net618 _04849_ _04850_ _04853_ vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__a31o_1
XFILLER_148_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10077__A _04765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout226_X net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout605_A _03349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1347_A net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09866__A _05367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13574__A1 _03137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09146_ net944 _04784_ vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__or2_1
XFILLER_148_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11585__B1 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07789__C1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09077_ top.CPU.registers.data\[936\] top.CPU.registers.data\[904\] top.CPU.registers.data\[808\]
+ top.CPU.registers.data\[776\] net975 net1281 vssd1 vssd1 vccd1 vccd1 _04716_ sky130_fd_sc_hd__mux4_1
XFILLER_163_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12129__A2 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08028_ top.CPU.registers.data\[596\] net1318 net849 top.CPU.registers.data\[628\]
+ net743 vssd1 vssd1 vccd1 vccd1 _03667_ sky130_fd_sc_hd__a221o_1
XFILLER_162_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold750 top.CPU.registers.data\[959\] vssd1 vssd1 vccd1 vccd1 net3307 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout974_A net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11337__B1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold761 top.CPU.registers.data\[473\] vssd1 vssd1 vccd1 vccd1 net3318 sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 top.CPU.registers.data\[528\] vssd1 vssd1 vccd1 vccd1 net3329 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold783 top.CPU.registers.data\[628\] vssd1 vssd1 vccd1 vccd1 net3340 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1302_X net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold794 top.CPU.registers.data\[125\] vssd1 vssd1 vccd1 vccd1 net3351 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14921__RESET_B net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09979_ net410 _05616_ vssd1 vssd1 vccd1 vccd1 _05618_ sky130_fd_sc_hd__or2_1
XANTENNA__10560__A1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout762_X net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12990_ top.SPI.register\[2\] net1354 net2610 _07419_ vssd1 vssd1 vccd1 vccd1 _07420_
+ sky130_fd_sc_hd__or4_1
Xhold1450 top.CPU.handler.state\[2\] vssd1 vssd1 vccd1 vccd1 net4007 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1461 top.CPU.control_unit.instruction\[2\] vssd1 vssd1 vccd1 vccd1 net4018 sky130_fd_sc_hd__dlygate4sd3_1
X_11941_ _06484_ net352 net232 net3255 vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__a22o_1
XANTENNA__08010__A _03613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07713__C1 net1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11872_ net3067 net189 vssd1 vssd1 vccd1 vccd1 _06768_ sky130_fd_sc_hd__nand2_1
XFILLER_44_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09540__S net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13611_ top.CPU.alu.program_counter\[24\] net1350 net582 vssd1 vssd1 vccd1 vccd1
+ _03034_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_28_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10823_ _05195_ _05267_ vssd1 vssd1 vccd1 vccd1 _06432_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_28_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_105_Right_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_118_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_118_clk
+ sky130_fd_sc_hd__clkbuf_8
X_16330_ clknet_leaf_67_clk _02539_ net1168 vssd1 vssd1 vccd1 vccd1 top.CPU.addressnew\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13542_ top.CPU.data_out\[29\] net589 net339 _02991_ vssd1 vssd1 vccd1 vccd1 _02527_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11812__A1 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10754_ net413 _06025_ _06366_ _06365_ _06014_ vssd1 vssd1 vccd1 vccd1 _06367_ sky130_fd_sc_hd__a32o_1
XFILLER_111_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09481__A2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11090__B net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16261_ clknet_leaf_33_clk _02471_ net1125 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.toreg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_13473_ net1397 net873 _02921_ net418 vssd1 vssd1 vccd1 vccd1 _02958_ sky130_fd_sc_hd__a31o_1
X_10685_ net410 _06201_ _06300_ _06299_ _05940_ vssd1 vssd1 vccd1 vccd1 _06301_ sky130_fd_sc_hd__o32a_1
XANTENNA__13565__A1 _03005_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15212_ net1546 _01422_ net1078 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_12424_ top.I2C.output_state\[20\] _06948_ vssd1 vssd1 vccd1 vccd1 _06949_ sky130_fd_sc_hd__nand2_1
X_16192_ net2526 _02402_ net1092 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[992\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09233__A2 net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12914__B _05429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10379__B2 top.CPU.handler.toreg\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11576__B1 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15143_ clknet_leaf_47_clk _01353_ net1131 vssd1 vssd1 vccd1 vccd1 top.I2C.data_out\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_127_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12355_ _06894_ _06899_ vssd1 vssd1 vccd1 vccd1 _00062_ sky130_fd_sc_hd__nor2_1
XANTENNA__08441__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11040__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07795__A2 net1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11306_ net3419 net291 _06704_ _06084_ vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__a22o_1
X_15074_ clknet_leaf_50_clk _00017_ net1130 vssd1 vssd1 vccd1 vccd1 top.I2C.output_state\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_12286_ _03754_ _06887_ _06889_ vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11328__B1 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11237_ net3086 net295 _06673_ net317 vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__a22o_1
XFILLER_68_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output67_A net1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11168_ net137 net3548 net299 vssd1 vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__mux2_1
XFILLER_95_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13237__S _06948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07952__C1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10119_ net417 net407 vssd1 vssd1 vccd1 vccd1 _05757_ sky130_fd_sc_hd__nand2_1
XFILLER_49_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14583__753 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 net2222 sky130_fd_sc_hd__inv_2
X_15976_ net2310 _02186_ net1088 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[776\]
+ sky130_fd_sc_hd__dfrtp_1
X_11099_ net3816 net302 _06607_ net484 vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__a22o_1
X_14927_ clknet_leaf_45_clk _01173_ net1160 vssd1 vssd1 vccd1 vccd1 top.CPU.alu.program_counter\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11500__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08855__A net1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14624__794 clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 net2263 sky130_fd_sc_hd__inv_2
XANTENNA__09450__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13809_ net3811 net333 net326 top.CPU.data_out\[11\] vssd1 vssd1 vccd1 vccd1 _02689_
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_109_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_109_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09457__C1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11281__A net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10606__A2 _05824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16528_ clknet_leaf_99_clk _02690_ net1257 vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__dfrtp_1
XANTENNA__15450__RESET_B net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12096__B net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16459_ clknet_leaf_87_clk _02621_ net1271 vssd1 vssd1 vccd1 vccd1 top.SPI.timem\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13005__B1 _07431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08680__B1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09000_ net950 _04635_ _04638_ net624 vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__a211o_1
XANTENNA__13556__A1 _06410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08590__A net1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08658__S1 net1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11567__B1 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07786__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10790__B2 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09902_ _04796_ _04798_ vssd1 vssd1 vccd1 vccd1 _05541_ sky130_fd_sc_hd__nand2_2
XFILLER_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout504 net505 vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_130_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout515 net523 vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08196__C1 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout526 net533 vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__clkbuf_4
XFILLER_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout537 _06574_ vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__buf_2
X_09833_ top.CPU.registers.data\[90\] net1305 net1028 top.CPU.registers.data\[122\]
+ net945 vssd1 vssd1 vccd1 vccd1 _05472_ sky130_fd_sc_hd__a221o_1
Xfanout548 net550 vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__clkbuf_4
Xfanout559 net561 vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout290_A net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout388_A net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07653__B _03262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09764_ top.CPU.registers.data\[411\] net1298 net1019 top.CPU.registers.data\[443\]
+ net916 vssd1 vssd1 vccd1 vccd1 _05403_ sky130_fd_sc_hd__a221o_1
XANTENNA__10360__A net1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08715_ top.CPU.registers.data\[301\] top.CPU.registers.data\[269\] net807 vssd1
+ vssd1 vccd1 vccd1 _04354_ sky130_fd_sc_hd__mux2_1
XANTENNA__13492__A0 top.CPU.data_out\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09695_ top.CPU.registers.data\[409\] net1306 net1029 top.CPU.registers.data\[441\]
+ net922 vssd1 vssd1 vccd1 vccd1 _05334_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout555_A net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout176_X net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1297_A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10845__A2 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08646_ net792 _04283_ _04284_ net720 vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_159_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08577_ top.CPU.registers.data\[335\] net1315 net846 top.CPU.registers.data\[367\]
+ net740 vssd1 vssd1 vccd1 vccd1 _04216_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout343_X net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout722_A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09999__A0 _04363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07528_ _03148_ net881 vssd1 vssd1 vccd1 vccd1 _03167_ sky130_fd_sc_hd__and2_4
XANTENNA__10519__B net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout510_X net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07459_ top.CPU.registers.data_out_r2_prev\[12\] vssd1 vssd1 vccd1 vccd1 _03099_
+ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_172_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08671__B1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11270__A2 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1252_X net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout608_X net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10470_ _06094_ _06095_ vssd1 vssd1 vccd1 vccd1 _06096_ sky130_fd_sc_hd__nand2_1
XFILLER_108_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12734__B _04598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11022__A2 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08423__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09129_ net678 _04766_ _04767_ vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__and3_1
XFILLER_136_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09620__C1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12140_ net563 _06652_ net236 vssd1 vssd1 vccd1 vccd1 _06838_ sky130_fd_sc_hd__and3_1
XFILLER_123_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08005__A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout977_X net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12071_ _06614_ net352 net178 net3485 vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__a22o_1
X_14270__440 clknet_leaf_150_clk vssd1 vssd1 vccd1 vccd1 net1909 sky130_fd_sc_hd__inv_2
XFILLER_151_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12750__A top.CPU.alu.program_counter\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold580 top.CPU.fetch.current_ra\[1\] vssd1 vssd1 vccd1 vccd1 net3137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold591 top.CPU.registers.data\[938\] vssd1 vssd1 vccd1 vccd1 net3148 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_110_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11022_ net3612 net218 _06568_ net317 vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_38_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14567__737 clknet_leaf_185_clk vssd1 vssd1 vccd1 vccd1 net2206 sky130_fd_sc_hd__inv_2
XFILLER_173_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11730__B1 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13057__S net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15830_ net2164 _02040_ net1222 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[630\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07563__B net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08011__Y _03650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14311__481 clknet_leaf_186_clk vssd1 vssd1 vccd1 vccd1 net1950 sky130_fd_sc_hd__inv_2
XFILLER_66_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11085__B net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14608__778 clknet_leaf_199_clk vssd1 vssd1 vccd1 vccd1 net2247 sky130_fd_sc_hd__inv_2
XANTENNA__12286__A1 _03754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15761_ net2095 _01971_ net1195 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[561\]
+ sky130_fd_sc_hd__dfrtp_1
X_12973_ top.I2C.bit_timer_counter\[3\] _07407_ vssd1 vssd1 vccd1 vccd1 _07408_ sky130_fd_sc_hd__or2_1
XANTENNA__09687__C1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1280 top.I2C.data_out\[14\] vssd1 vssd1 vccd1 vccd1 net3837 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09151__A1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1291 top.CPU.registers.data\[922\] vssd1 vssd1 vccd1 vccd1 net3848 sky130_fd_sc_hd__dlygate4sd3_1
X_11924_ net3517 net184 net341 _06314_ vssd1 vssd1 vccd1 vccd1 _01642_ sky130_fd_sc_hd__a22o_1
XANTENNA__15279__RESET_B net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15692_ net2026 _01902_ net1070 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[492\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_75_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11813__B net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09439__C1 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11855_ _06691_ net233 net152 net2906 vssd1 vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__a22o_1
XFILLER_26_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10806_ net305 _06414_ net394 vssd1 vssd1 vccd1 vccd1 _06416_ sky130_fd_sc_hd__a21o_1
XFILLER_159_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11786_ net468 _06632_ net238 net162 net3122 vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__a32o_1
XANTENNA__10429__B _06056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16313_ clknet_leaf_83_clk _02522_ net1261 vssd1 vssd1 vccd1 vccd1 top.CPU.data_out\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_13525_ _03783_ net584 vssd1 vssd1 vccd1 vccd1 _02983_ sky130_fd_sc_hd__and2_1
X_10737_ _05275_ net446 vssd1 vssd1 vccd1 vccd1 _06351_ sky130_fd_sc_hd__nand2_1
XFILLER_9_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16244_ clknet_leaf_44_clk _02454_ net1124 vssd1 vssd1 vccd1 vccd1 top.CPU.control_unit.instruction\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13456_ top.CPU.handler.toreg\[17\] _02949_ net123 vssd1 vssd1 vccd1 vccd1 _02483_
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10668_ _04732_ _05564_ _05531_ _05279_ vssd1 vssd1 vccd1 vccd1 _06285_ sky130_fd_sc_hd__a211oi_1
XFILLER_12_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09206__A2 net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11549__B1 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12407_ top.SPI.register\[2\] _06932_ net2610 vssd1 vssd1 vccd1 vccd1 _00070_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_11_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16175_ net2509 _02385_ net1097 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[975\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10445__A net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10599_ _06135_ _06218_ net387 vssd1 vssd1 vccd1 vccd1 _06219_ sky130_fd_sc_hd__mux2_1
X_13387_ net1368 _02908_ net667 vssd1 vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__mux2_1
XFILLER_12_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07768__A2 _03405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
X_15126_ clknet_leaf_53_clk top.I2C.sda_oeb_n net1135 vssd1 vssd1 vccd1 vccd1 top.I2C.sda_oeb
+ sky130_fd_sc_hd__dfrtp_1
Xoutput118 net118 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_58_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12338_ net2598 _05084_ net1174 vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15057_ clknet_leaf_51_clk _00061_ net1132 vssd1 vssd1 vccd1 vccd1 top.I2C.output_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_75_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12269_ net3254 _06428_ net432 vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__mux2_1
XFILLER_101_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10524__B2 top.CPU.handler.toreg\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11721__B1 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07925__C1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08193__A2 net1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13762__Y _03093_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15959_ net2293 _02169_ net1182 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[759\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09678__C1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09142__A1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08500_ net694 _04137_ _04138_ vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__or3_1
X_09480_ net795 _05111_ _05118_ _03110_ net643 vssd1 vssd1 vccd1 vccd1 _05119_ sky130_fd_sc_hd__a221o_1
XANTENNA__09693__A2 _05330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12029__A1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08431_ net796 _04065_ _04066_ net750 vssd1 vssd1 vccd1 vccd1 _04070_ sky130_fd_sc_hd__o211a_1
X_08362_ top.CPU.registers.data\[850\] net1317 net848 top.CPU.registers.data\[882\]
+ net742 vssd1 vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__a221o_1
XFILLER_51_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11788__B1 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08102__C1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08293_ top.CPU.registers.data\[435\] top.CPU.registers.data\[403\] net826 vssd1
+ vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__mux2_1
XANTENNA__11252__A2 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout136_A _05879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10058__C _03185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10460__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08405__B1 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09602__C1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12046__S net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout303_A _06604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14254__424 clknet_leaf_165_clk vssd1 vssd1 vccd1 vccd1 net1893 sky130_fd_sc_hd__inv_2
XFILLER_133_746 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11960__B1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11885__S net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1212_A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08169__C1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout301 _06604_ vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07664__A _03262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09355__S net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout312 net315 vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__buf_4
Xfanout323 net324 vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__buf_4
XANTENNA__16399__D net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout334 net335 vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__buf_2
XFILLER_87_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout293_X net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout672_A net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10802__B net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11712__B1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout345 net346 vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__buf_4
XFILLER_113_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout356 _06732_ vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11186__A net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09816_ top.CPU.registers.data\[762\] net1394 net838 top.CPU.registers.data\[730\]
+ net733 vssd1 vssd1 vccd1 vccd1 _05455_ sky130_fd_sc_hd__a221o_1
Xfanout367 net369 vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__buf_4
Xfanout378 net380 vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1000_X net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout389 net392 vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__clkbuf_4
XFILLER_143_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07931__A2 net1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09747_ top.CPU.registers.data\[827\] top.CPU.registers.data\[795\] net827 vssd1
+ vssd1 vccd1 vccd1 _05386_ sky130_fd_sc_hd__mux2_1
XFILLER_100_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13465__B1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout460_X net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09669__C1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout937_A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11473__X _06728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09678_ top.CPU.registers.data\[985\] net1336 net869 top.CPU.registers.data\[1017\]
+ net732 vssd1 vssd1 vccd1 vccd1 _05317_ sky130_fd_sc_hd__a221o_1
XANTENNA__09684__A2 net1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07603__S net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09090__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08629_ net792 _04267_ _04266_ net720 vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__o211a_1
XFILLER_15_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11491__A2 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08892__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11640_ _06036_ net203 net426 net3590 vssd1 vssd1 vccd1 vccd1 _01911_ sky130_fd_sc_hd__a22o_1
XFILLER_30_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11779__B1 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11571_ _06682_ net259 net246 net2712 vssd1 vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__a22o_1
XANTENNA__11243__A2 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12745__A top.CPU.alu.program_counter\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09841__C1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13310_ _02830_ _02851_ vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__nor2_1
XFILLER_7_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07998__A2 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10522_ _06142_ _06144_ _06145_ vssd1 vssd1 vccd1 vccd1 _06146_ sky130_fd_sc_hd__or3b_1
XFILLER_109_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10453_ net413 _06079_ vssd1 vssd1 vccd1 vccd1 _06080_ sky130_fd_sc_hd__nor2_1
X_13241_ top.I2C.output_state\[28\] _02803_ vssd1 vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__nand2_2
XFILLER_170_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13172_ _06916_ _03120_ top.I2C.byte_manager_state\[2\] vssd1 vssd1 vccd1 vccd1 _02756_
+ sky130_fd_sc_hd__mux2_1
X_10384_ _03719_ _03789_ _05965_ _06012_ net370 vssd1 vssd1 vccd1 vccd1 _06013_ sky130_fd_sc_hd__a311o_1
XANTENNA__10754__A1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11951__B1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12123_ net3965 net653 _06829_ vssd1 vssd1 vccd1 vccd1 _01501_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_92_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12054_ _06601_ _06731_ vssd1 vssd1 vccd1 vccd1 _06796_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_53_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11703__B1 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09372__A1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11096__A net1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11005_ net524 _06557_ vssd1 vssd1 vccd1 vccd1 _06558_ sky130_fd_sc_hd__nor2_1
XANTENNA__10204__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08580__C1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout890 _02829_ vssd1 vssd1 vccd1 vccd1 net890 sky130_fd_sc_hd__buf_2
X_15813_ net2147 _02023_ net1083 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[613\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07922__A2 net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13456__A0 top.CPU.handler.toreg\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12259__A1 _06230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_13_0_clk_X clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15744_ net2078 _01954_ net1094 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[544\]
+ sky130_fd_sc_hd__dfrtp_1
X_12956_ net1363 top.CPU.alu.program_counter\[31\] vssd1 vssd1 vccd1 vccd1 _07395_
+ sky130_fd_sc_hd__and2b_1
XFILLER_80_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08332__C1 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11907_ net3291 net186 net352 _05935_ vssd1 vssd1 vccd1 vccd1 _01659_ sky130_fd_sc_hd__a22o_1
X_15675_ net2009 _01885_ net1213 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[475\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11482__A2 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12887_ _07331_ _07332_ net127 vssd1 vssd1 vccd1 vccd1 _07333_ sky130_fd_sc_hd__o21ai_1
XFILLER_33_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13759__A1 _02803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11838_ _06669_ net209 net155 net2685 vssd1 vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__a22o_1
X_14695__865 clknet_leaf_183_clk vssd1 vssd1 vccd1 vccd1 net2334 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_99_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12655__A _03100_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11769_ _06612_ net202 net161 net3394 vssd1 vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_40_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_174_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10442__A0 _03684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13508_ _04390_ _02966_ vssd1 vssd1 vccd1 vccd1 _02974_ sky130_fd_sc_hd__nor2_1
XFILLER_146_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10993__B2 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16227_ clknet_leaf_30_clk _02437_ net1152 vssd1 vssd1 vccd1 vccd1 top.CPU.control_unit.instruction\[3\]
+ sky130_fd_sc_hd__dfrtp_2
X_14238__408 clknet_leaf_150_clk vssd1 vssd1 vccd1 vccd1 net1877 sky130_fd_sc_hd__inv_2
X_13439_ _02875_ _02937_ _02939_ vssd1 vssd1 vccd1 vccd1 _02941_ sky130_fd_sc_hd__a21o_1
XFILLER_61_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09286__S1 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12195__B1 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08399__C1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11537__A3 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16158_ net2492 _02368_ net1239 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[958\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_115_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11942__B1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15109_ net1491 _01322_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r2_prev\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11558__X _06741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08980_ top.CPU.registers.data\[425\] top.CPU.registers.data\[393\] net805 vssd1
+ vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__mux2_1
X_16089_ net2423 _02299_ net1245 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[889\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10903__A net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09175__S net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07931_ top.CPU.registers.data\[348\] net1303 net1023 top.CPU.registers.data\[380\]
+ net943 vssd1 vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__a221o_1
XANTENNA__08166__A2 net1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07862_ top.CPU.registers.data\[317\] net1007 net931 vssd1 vssd1 vccd1 vccd1 _03501_
+ sky130_fd_sc_hd__a21o_1
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09601_ top.CPU.registers.data\[160\] top.CPU.registers.data\[128\] net810 vssd1
+ vssd1 vccd1 vccd1 _05240_ sky130_fd_sc_hd__mux2_1
XANTENNA__08571__C1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11170__B2 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07793_ net621 _03429_ _03430_ _03431_ vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__a31o_1
XANTENNA__08586__Y _04225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09115__A1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09532_ top.CPU.registers.data\[577\] net1335 net868 top.CPU.registers.data\[609\]
+ net780 vssd1 vssd1 vccd1 vccd1 _05171_ sky130_fd_sc_hd__a221o_1
XFILLER_58_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08323__C1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09463_ net795 _05091_ _05092_ net723 vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout253_A _06733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08414_ _04020_ _04051_ vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__nand2_1
X_09394_ net797 _05027_ _05028_ net727 vssd1 vssd1 vccd1 vccd1 _05033_ sky130_fd_sc_hd__o211a_1
XANTENNA__11225__A2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08345_ net627 _03982_ _03983_ _03979_ vssd1 vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__a31o_4
XANTENNA__08626__B1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12565__A _06371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout420_A net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1162_A net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_31_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout518_A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout139_X net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08276_ net629 _03902_ _03904_ _03912_ _03914_ vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__a32o_4
XFILLER_149_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12186__B1 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13396__A net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1107 net1108 vssd1 vssd1 vccd1 vccd1 net1107 sky130_fd_sc_hd__clkbuf_4
Xfanout1118 net1147 vssd1 vssd1 vccd1 vccd1 net1118 sky130_fd_sc_hd__clkbuf_2
Xfanout120 net122 vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__clkbuf_4
Xfanout1129 net1136 vssd1 vssd1 vccd1 vccd1 net1129 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_98_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_98_clk sky130_fd_sc_hd__clkbuf_8
Xfanout131 _06464_ vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout675_X net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout142 _06253_ vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__buf_2
Xfanout153 net155 vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__clkbuf_8
XFILLER_102_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout164 _06757_ vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__buf_6
XFILLER_101_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout175 _06825_ vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08562__C1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout186 net187 vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__buf_4
XFILLER_87_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout197 net202 vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__clkbuf_4
XFILLER_101_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout842_X net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09106__A1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12810_ top.CPU.alu.program_counter\[16\] _07263_ net1361 vssd1 vssd1 vccd1 vccd1
+ _01179_ sky130_fd_sc_hd__mux2_1
XFILLER_16_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13790_ net19 net1050 net885 net2955 vssd1 vssd1 vccd1 vccd1 _02671_ sky130_fd_sc_hd__o22a_1
X_14382__552 clknet_leaf_165_clk vssd1 vssd1 vccd1 vccd1 net2021 sky130_fd_sc_hd__inv_2
XANTENNA__12110__B1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12741_ top.CPU.alu.program_counter\[10\] _07200_ net1360 vssd1 vssd1 vccd1 vccd1
+ _01173_ sky130_fd_sc_hd__mux2_1
X_14679__849 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 net2318 sky130_fd_sc_hd__inv_2
XANTENNA__12178__C net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10672__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15460_ net1794 _01670_ net1219 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[260\]
+ sky130_fd_sc_hd__dfrtp_1
X_12672_ top.CPU.alu.program_counter\[4\] _04955_ vssd1 vssd1 vccd1 vccd1 _07138_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_13_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423__593 clknet_leaf_76_clk vssd1 vssd1 vccd1 vccd1 net2062 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ _06391_ net3336 net214 vssd1 vssd1 vccd1 vccd1 _01926_ sky130_fd_sc_hd__mux2_1
XANTENNA__10547__X _06170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15391_ net1725 _01601_ net1220 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[191\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_129_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12475__A _04090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09814__C1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_22_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__11767__A3 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11554_ _06667_ net261 net248 net2920 vssd1 vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__a22o_1
XANTENNA__09290__B1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10505_ _04193_ _05289_ _06128_ vssd1 vssd1 vccd1 vccd1 _06129_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_94_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11485_ net490 net474 _06615_ net256 net2845 vssd1 vssd1 vccd1 vccd1 _02039_ sky130_fd_sc_hd__a32o_1
X_16012_ net2346 _02222_ net1079 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[812\]
+ sky130_fd_sc_hd__dfrtp_1
X_13224_ _02776_ net3468 _02795_ vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__mux2_1
X_10436_ net512 _05585_ _06062_ _06059_ _05295_ vssd1 vssd1 vccd1 vccd1 _06063_ sky130_fd_sc_hd__a311oi_1
XANTENNA__09042__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10727__B2 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11924__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09593__A1 net1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08396__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13155_ top.I2C.output_state\[3\] top.I2C.output_state\[10\] top.I2C.output_state\[11\]
+ top.I2C.output_state\[16\] vssd1 vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__or4_1
X_10367_ _03822_ _03889_ net375 vssd1 vssd1 vccd1 vccd1 _05997_ sky130_fd_sc_hd__mux2_1
XFILLER_98_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_362 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12106_ top.CPU.registers.data\[99\] net653 _03185_ vssd1 vssd1 vccd1 vccd1 _06821_
+ sky130_fd_sc_hd__o21a_1
XFILLER_124_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11538__B net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10298_ net445 _05930_ _05929_ _05910_ vssd1 vssd1 vccd1 vccd1 _05931_ sky130_fd_sc_hd__o211ai_4
X_13086_ top.CPU.data_out\[21\] net2755 net558 vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__mux2_1
XANTENNA__13677__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_89_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_89_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09345__A1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12037_ _06230_ net3701 net150 vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__mux2_1
XANTENNA__11152__A1 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13990__160 clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 net1629 sky130_fd_sc_hd__inv_2
XFILLER_65_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08305__C1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15727_ net2061 _01937_ net1104 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[527\]
+ sky130_fd_sc_hd__dfrtp_1
X_12939_ top.CPU.alu.program_counter\[28\] _07362_ top.CPU.alu.program_counter\[29\]
+ vssd1 vssd1 vccd1 vccd1 _07380_ sky130_fd_sc_hd__a21oi_1
XFILLER_61_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08320__A2 _03955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15658_ net1992 _01868_ net1087 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[458\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11207__A2 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08608__B1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13601__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15589_ net1923 _01799_ net1062 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[389\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09805__C1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_13_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_32_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08130_ net627 _03768_ _03767_ net606 vssd1 vssd1 vccd1 vccd1 _03769_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_32_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09281__A0 _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09820__A2 net1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10966__B2 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08061_ top.CPU.registers.data_out_r2_prev\[20\] net685 net618 _03693_ _03699_ vssd1
+ vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__o2111a_1
XANTENNA__07831__A1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12168__B1 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09033__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10718__A1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11915__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10633__A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11391__A1 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07595__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08963_ _04567_ _04599_ vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__nor2_1
XANTENNA__13668__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08139__A2 net1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07914_ top.CPU.registers.data\[764\] net1384 net995 top.CPU.registers.data\[732\]
+ net919 vssd1 vssd1 vccd1 vccd1 _03553_ sky130_fd_sc_hd__a221o_1
XFILLER_97_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08894_ _04501_ _04532_ vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__nor2_1
XFILLER_111_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1008_A net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08544__C1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07898__A1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07845_ net674 _03482_ _03483_ net604 vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__a31o_1
XANTENNA__12891__A1 top.CPU.alu.program_counter\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout370_A net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14366__536 clknet_leaf_153_clk vssd1 vssd1 vccd1 vccd1 net2005 sky130_fd_sc_hd__inv_2
XANTENNA__11694__A2 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout468_A net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07776_ net944 _03414_ net608 vssd1 vssd1 vccd1 vccd1 _03415_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_123_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14110__280 clknet_leaf_151_clk vssd1 vssd1 vccd1 vccd1 net1749 sky130_fd_sc_hd__inv_2
X_09515_ _05133_ _05140_ _05152_ _05153_ vssd1 vssd1 vccd1 vccd1 _05154_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_140_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14407__577 clknet_leaf_186_clk vssd1 vssd1 vccd1 vccd1 net2046 sky130_fd_sc_hd__inv_2
XANTENNA_fanout256_X net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout635_A net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1377_A net1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09446_ _05084_ vssd1 vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__inv_2
X_09377_ net679 _04996_ _04997_ net613 vssd1 vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout423_X net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout802_A net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08328_ top.CPU.registers.data\[83\] net1296 net1016 top.CPU.registers.data\[115\]
+ net955 vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__a221o_1
XANTENNA__11749__A3 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08075__A1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09272__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_5 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10957__B2 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08259_ top.CPU.registers.data\[86\] net1307 net1030 top.CPU.registers.data\[118\]
+ net959 vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1332_X net1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07676__X _03315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11270_ net2989 net296 _06692_ net321 vssd1 vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__a22o_1
XANTENNA__10709__A1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout792_X net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11906__B1 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10221_ _05432_ net510 vssd1 vssd1 vccd1 vccd1 _05856_ sky130_fd_sc_hd__nor2_1
XFILLER_161_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11382__A1 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10152_ _05644_ _05648_ net306 vssd1 vssd1 vccd1 vccd1 _05789_ sky130_fd_sc_hd__mux2_1
X_13974__144 clknet_leaf_174_clk vssd1 vssd1 vccd1 vccd1 net1613 sky130_fd_sc_hd__inv_2
XFILLER_79_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14960_ clknet_leaf_89_clk _01205_ net1273 vssd1 vssd1 vccd1 vccd1 top.SPI.dcx sky130_fd_sc_hd__dfrtp_1
X_10083_ _05717_ _05720_ net388 vssd1 vssd1 vccd1 vccd1 _05721_ sky130_fd_sc_hd__mux2_1
XFILLER_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11077__C net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold9 _00028_ vssd1 vssd1 vccd1 vccd1 net2566 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_87_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13573__B top.CPU.handler.state\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input29_A DAT_I[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11093__B net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13773_ net32 net1051 net886 net4019 vssd1 vssd1 vccd1 vccd1 _02654_ sky130_fd_sc_hd__a22o_1
XANTENNA__11437__A2 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13831__B1 _03096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10985_ net3576 net217 _06545_ net321 vssd1 vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__a22o_1
XFILLER_16_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08302__A2 net1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15512_ net1846 _01722_ net1102 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[312\]
+ sky130_fd_sc_hd__dfrtp_1
X_12724_ _07184_ vssd1 vssd1 vccd1 vccd1 _07185_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16492_ clknet_leaf_41_clk _02654_ net1116 vssd1 vssd1 vccd1 vccd1 top.mmio.mem_data_i\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15443_ net1777 _01653_ net1187 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[243\]
+ sky130_fd_sc_hd__dfrtp_1
X_12655_ _03100_ _05087_ vssd1 vssd1 vccd1 vccd1 _07123_ sky130_fd_sc_hd__xnor2_1
XFILLER_90_52 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11606_ _06033_ net3327 net214 vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__mux2_1
XANTENNA__08066__A1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15374_ net1708 _01584_ net1190 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[174\]
+ sky130_fd_sc_hd__dfrtp_1
X_12586_ _06919_ _07054_ _07089_ vssd1 vssd1 vccd1 vccd1 _07090_ sky130_fd_sc_hd__and3_1
XFILLER_156_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09263__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09802__A2 net1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11537_ net483 _06311_ net355 net251 net3128 vssd1 vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__a32o_1
XFILLER_172_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold409 top.CPU.registers.data\[446\] vssd1 vssd1 vccd1 vccd1 net2966 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09015__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11468_ net147 net3688 net265 vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__mux2_1
XFILLER_99_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13207_ top.I2C.data_out\[20\] net892 _02755_ vssd1 vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__mux2_1
XANTENNA__14921__Q top.CPU.alu.program_counter\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13362__A2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10419_ _03685_ net506 net509 _03721_ vssd1 vssd1 vccd1 vccd1 _06047_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__10453__A net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15475__RESET_B net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11399_ _06527_ net283 net269 net3344 vssd1 vssd1 vccd1 vccd1 _02112_ sky130_fd_sc_hd__a22o_1
XFILLER_135_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08774__C1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13138_ net4024 top.CPU.data_out\[0\] _07418_ vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__mux2_1
XFILLER_112_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10172__B _05808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14053__223 clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 net1692 sky130_fd_sc_hd__inv_2
XANTENNA__09318__A1 _04955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13764__A net1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13114__A2 net1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13069_ top.CPU.data_out\[4\] net3438 net559 vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__mux2_1
XANTENNA__10740__X _06354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1109 top.CPU.data_out\[5\] vssd1 vssd1 vccd1 vccd1 net3666 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_24_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_2_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__11125__A1 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08526__C1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_119_Right_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12873__A1 top.CPU.alu.program_counter\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07630_ _03265_ _03267_ _03268_ _03262_ vssd1 vssd1 vccd1 vccd1 _03269_ sky130_fd_sc_hd__a31oi_2
XANTENNA__10884__B1 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07561_ net1047 _03163_ net1038 vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__and3_2
XANTENNA__11428__A2 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13822__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09300_ top.CPU.registers.data\[548\] top.CPU.registers.data\[516\] net992 vssd1
+ vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__mux2_1
XANTENNA__07727__S1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07492_ top.wm.curr_state\[0\] vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__inv_2
XFILLER_110_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09231_ top.CPU.registers.data\[645\] net1310 net840 top.CPU.registers.data\[677\]
+ net702 vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__a221o_1
XFILLER_22_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09162_ net789 _04799_ _04800_ net692 vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__o211a_1
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14751__921 clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 net2390 sky130_fd_sc_hd__inv_2
XANTENNA__10939__B2 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08113_ net798 _03750_ _03751_ net752 vssd1 vssd1 vccd1 vccd1 _03752_ sky130_fd_sc_hd__o211a_1
X_09093_ _04730_ _04731_ vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__nand2_2
XFILLER_174_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout216_A net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08044_ net880 net451 _03651_ vssd1 vssd1 vccd1 vccd1 _03683_ sky130_fd_sc_hd__o21a_2
XANTENNA__08532__S net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold910 top.SPI.state\[1\] vssd1 vssd1 vccd1 vccd1 net3467 sky130_fd_sc_hd__dlygate4sd3_1
Xhold921 top.CPU.registers.data\[837\] vssd1 vssd1 vccd1 vccd1 net3478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold932 top.CPU.registers.data\[272\] vssd1 vssd1 vccd1 vccd1 net3489 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold943 top.CPU.registers.data\[50\] vssd1 vssd1 vccd1 vccd1 net3500 sky130_fd_sc_hd__dlygate4sd3_1
X_13958__128 clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 net1597 sky130_fd_sc_hd__inv_2
Xhold954 top.CPU.registers.data\[514\] vssd1 vssd1 vccd1 vccd1 net3511 sky130_fd_sc_hd__dlygate4sd3_1
Xhold965 top.CPU.registers.data\[259\] vssd1 vssd1 vccd1 vccd1 net3522 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08765__C1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold976 top.CPU.registers.data\[222\] vssd1 vssd1 vccd1 vccd1 net3533 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_164_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_1_0_clk_X clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold987 top.CPU.registers.data\[656\] vssd1 vssd1 vccd1 vccd1 net3544 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_164_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold998 top.CPU.registers.data\[982\] vssd1 vssd1 vccd1 vccd1 net3555 sky130_fd_sc_hd__dlygate4sd3_1
X_09995_ _04698_ net372 vssd1 vssd1 vccd1 vccd1 _05634_ sky130_fd_sc_hd__nor2_1
X_13904__74 clknet_leaf_194_clk vssd1 vssd1 vccd1 vccd1 net1543 sky130_fd_sc_hd__inv_2
XANTENNA_fanout585_A net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_134_Left_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09309__A1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11893__S net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08780__A2 net1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08946_ _04583_ _04584_ net673 vssd1 vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__o21a_1
XFILLER_9_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09216__X _04855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08877_ net784 _04514_ _04515_ net738 vssd1 vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__o211a_1
XFILLER_151_25 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout373_X net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout752_A net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11194__A _06213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07828_ net791 _03461_ _03462_ net719 vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__o211a_1
XANTENNA__11419__A2 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout540_X net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07759_ top.CPU.registers.data\[318\] top.CPU.registers.data\[286\] net833 vssd1
+ vssd1 vccd1 vccd1 _03398_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1282_X net1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout638_X net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08296__A1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10770_ _05671_ _06045_ _06140_ vssd1 vssd1 vccd1 vccd1 _06382_ sky130_fd_sc_hd__o21a_1
XANTENNA__12092__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10809__Y _06419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_143_Left_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09429_ top.CPU.registers.data\[226\] top.CPU.registers.data\[194\] net986 vssd1
+ vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout805_X net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12440_ net898 _06956_ vssd1 vssd1 vccd1 vccd1 _00053_ sky130_fd_sc_hd__nor2_1
XANTENNA__09245__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14494__664 clknet_leaf_150_clk vssd1 vssd1 vccd1 vccd1 net2133 sky130_fd_sc_hd__inv_2
X_12371_ top.I2C.within_byte_counter_writing\[0\] top.I2C.within_byte_counter_writing\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06911_ sky130_fd_sc_hd__nand2_1
XANTENNA__13592__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13201__X _02780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11322_ net3640 net289 net357 _06373_ vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__a22o_1
XANTENNA__09538__S net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13568__B _06309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15090_ net1472 _01303_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r2_prev\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_119_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12472__B _03984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09548__A1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11253_ net524 _06213_ net542 vssd1 vssd1 vccd1 vccd1 _06682_ sky130_fd_sc_hd__and3_1
X_14037__207 clknet_leaf_168_clk vssd1 vssd1 vccd1 vccd1 net1676 sky130_fd_sc_hd__inv_2
XANTENNA__10273__A net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_152_Left_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10204_ _05837_ _05839_ net392 vssd1 vssd1 vccd1 vccd1 _05840_ sky130_fd_sc_hd__mux2_1
XANTENNA__12899__S net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11184_ net132 net430 vssd1 vssd1 vccd1 vccd1 _06651_ sky130_fd_sc_hd__and2_1
XFILLER_121_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07574__A3 net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10135_ net3676 net227 net321 _05772_ vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_89_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15992_ net2326 _02202_ net1150 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[792\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11107__A1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14943_ clknet_leaf_68_clk _01189_ net1165 vssd1 vssd1 vccd1 vccd1 top.CPU.alu.program_counter\[26\]
+ sky130_fd_sc_hd__dfrtp_4
X_10066_ net305 _05703_ _05702_ vssd1 vssd1 vccd1 vccd1 _05704_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11658__A2 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10720__B _06333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09181__C1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09720__A1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16613_ net1346 vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__clkbuf_1
X_13825_ net2810 net338 net329 top.CPU.data_out\[27\] vssd1 vssd1 vccd1 vccd1 _02705_
+ sky130_fd_sc_hd__a22o_1
XFILLER_91_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08684__Y _04323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_161_Left_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16544_ clknet_leaf_84_clk net3773 net1263 vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__dfrtp_1
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13756_ top.I2C.I2C_state\[0\] _03088_ vssd1 vssd1 vccd1 vccd1 _03090_ sky130_fd_sc_hd__nand2_1
XANTENNA__12083__A2 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10968_ net3682 net217 _06535_ net314 vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__a22o_1
XFILLER_44_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12707_ _07158_ _07159_ _07156_ vssd1 vssd1 vccd1 vccd1 _07170_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09302__A net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11551__B net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16475_ clknet_leaf_88_clk _02637_ net1273 vssd1 vssd1 vccd1 vccd1 top.SPI.timem\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_14735__905 clknet_leaf_178_clk vssd1 vssd1 vccd1 vccd1 net2374 sky130_fd_sc_hd__inv_2
X_13687_ net2644 net336 vssd1 vssd1 vccd1 vccd1 _02615_ sky130_fd_sc_hd__and2_1
X_10899_ net662 _06105_ net436 vssd1 vssd1 vccd1 vccd1 _06493_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_80_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15426_ net1760 _01636_ net1171 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[226\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08039__A1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12638_ top.I2C.output_state\[14\] net3923 vssd1 vssd1 vccd1 vccd1 _00009_ sky130_fd_sc_hd__and2_1
XFILLER_129_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15357_ net1691 _01567_ net1119 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[157\]
+ sky130_fd_sc_hd__dfrtp_1
X_12569_ _06124_ _06210_ _07073_ vssd1 vssd1 vccd1 vccd1 _07074_ sky130_fd_sc_hd__or3_1
XANTENNA__12663__A top.CPU.alu.program_counter\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07798__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold206 top.SPI.percount\[2\] vssd1 vssd1 vccd1 vccd1 net2763 sky130_fd_sc_hd__dlygate4sd3_1
X_15288_ net1622 _01498_ net1103 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[88\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12382__B _03126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold217 top.CPU.registers.data\[160\] vssd1 vssd1 vccd1 vccd1 net2774 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold228 top.SPI.parameters\[28\] vssd1 vssd1 vccd1 vccd1 net2785 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_170_Left_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11279__A net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09539__A1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold239 _02595_ vssd1 vssd1 vccd1 vccd1 net2796 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_125_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08747__C1 _03116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout708 net709 vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout719 net722 vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__clkbuf_4
XFILLER_140_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08800_ top.CPU.registers.data\[172\] top.CPU.registers.data\[140\] net969 vssd1
+ vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__mux2_1
XANTENNA__07565__A3 net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09780_ net679 _05408_ _05409_ net916 vssd1 vssd1 vccd1 vccd1 _05419_ sky130_fd_sc_hd__o211a_1
XFILLER_100_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10911__A net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07970__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08731_ net1366 _04366_ _04369_ vssd1 vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11649__A2 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09172__C1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1290 net1291 vssd1 vssd1 vccd1 vccd1 net1290 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16444__RESET_B net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08662_ net1367 _04297_ _04300_ vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__o21a_1
XFILLER_27_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07613_ _03108_ net1279 _03158_ vssd1 vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__and3_2
X_08593_ net1284 _04230_ _04231_ _04229_ vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__o31a_1
XFILLER_35_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout166_A _06757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10609__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08278__A1 _03916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07544_ _03180_ _03181_ vssd1 vssd1 vccd1 vccd1 _03183_ sky130_fd_sc_hd__nor2_1
XANTENNA__09475__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13271__B2 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14181__351 clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 net1820 sky130_fd_sc_hd__inv_2
XFILLER_14_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07475_ net1365 vssd1 vssd1 vccd1 vccd1 _03115_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_157_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14478__648 clknet_leaf_165_clk vssd1 vssd1 vccd1 vccd1 net2117 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_157_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1075_A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09214_ net625 _04851_ _04852_ net604 vssd1 vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__a31o_1
XFILLER_167_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10077__B net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11888__S net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11034__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09145_ top.CPU.registers.data\[807\] top.CPU.registers.data\[775\] net995 vssd1
+ vssd1 vccd1 vccd1 _04784_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14222__392 clknet_leaf_166_clk vssd1 vssd1 vccd1 vccd1 net1861 sky130_fd_sc_hd__inv_2
XANTENNA_fanout1242_A net1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout219_X net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07789__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14519__689 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 net2158 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_135_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09076_ net1284 _04713_ _04714_ vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__or3_1
XANTENNA__08450__A1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08027_ _03662_ _03665_ net636 vssd1 vssd1 vccd1 vccd1 _03666_ sky130_fd_sc_hd__a21oi_1
XFILLER_150_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold740 top.CPU.registers.data\[643\] vssd1 vssd1 vccd1 vccd1 net3297 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1030_X net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold751 top.CPU.registers.data\[193\] vssd1 vssd1 vccd1 vccd1 net3308 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold762 top.CPU.registers.data\[227\] vssd1 vssd1 vccd1 vccd1 net3319 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold773 top.CPU.registers.data\[504\] vssd1 vssd1 vccd1 vccd1 net3330 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold784 top.CPU.registers.data\[485\] vssd1 vssd1 vccd1 vccd1 net3341 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout490_X net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold795 top.CPU.registers.data\[722\] vssd1 vssd1 vccd1 vccd1 net3352 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout967_A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10380__X _06010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09978_ net410 _05616_ vssd1 vssd1 vccd1 vccd1 _05617_ sky130_fd_sc_hd__nor2_1
X_08929_ top.CPU.registers.data\[426\] top.CPU.registers.data\[394\] top.CPU.registers.data\[298\]
+ top.CPU.registers.data\[266\] net972 net1281 vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__mux4_1
XFILLER_76_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout755_X net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1440 top.CPU.handler.toreg\[20\] vssd1 vssd1 vccd1 vccd1 net3997 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1451 top.CPU.handler.toreg\[8\] vssd1 vssd1 vccd1 vccd1 net4008 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08505__A2 net1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11940_ _06481_ net352 net232 net3531 vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__a22o_1
Xhold1462 top.mmio.mem_data_i\[8\] vssd1 vssd1 vccd1 vccd1 net4019 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08910__C1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16114__RESET_B net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout922_X net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11871_ _06707_ net241 net191 net3005 vssd1 vssd1 vccd1 vccd1 _01691_ sky130_fd_sc_hd__a22o_1
X_13610_ net1350 _05958_ vssd1 vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__nand2_1
X_10822_ _05672_ _06114_ _06120_ _05665_ vssd1 vssd1 vccd1 vccd1 _06431_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_28_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12065__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09466__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13541_ _03508_ net584 vssd1 vssd1 vccd1 vccd1 _02991_ sky130_fd_sc_hd__and2_1
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10753_ _05672_ _06026_ vssd1 vssd1 vccd1 vccd1 _06366_ sky130_fd_sc_hd__nand2_1
XFILLER_13_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09218__A0 _04855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16260_ clknet_leaf_34_clk _02470_ net1121 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.toreg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_158_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13472_ net3986 _02957_ net123 vssd1 vssd1 vccd1 vccd1 _02491_ sky130_fd_sc_hd__mux2_1
X_10684_ _05945_ _06139_ vssd1 vssd1 vccd1 vccd1 _06300_ sky130_fd_sc_hd__nor2_1
XANTENNA__08961__A _04567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15211_ net1545 _01421_ net1065 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11798__S net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12423_ top.I2C.within_byte_counter_reading\[2\] top.I2C.within_byte_counter_reading\[1\]
+ top.I2C.within_byte_counter_reading\[0\] vssd1 vssd1 vccd1 vccd1 _06948_ sky130_fd_sc_hd__and3_2
X_16191_ net2525 _02401_ net1222 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[991\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12483__A _03819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15142_ clknet_leaf_46_clk _01352_ net1140 vssd1 vssd1 vccd1 vccd1 top.I2C.data_out\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08977__C1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12354_ net1341 top.I2C.output_state\[22\] net3208 vssd1 vssd1 vccd1 vccd1 _06899_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__08172__S net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11305_ net3120 net290 net358 _06056_ vssd1 vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__a22o_1
X_15073_ clknet_leaf_52_clk _00051_ net1132 vssd1 vssd1 vccd1 vccd1 top.I2C.output_state\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_141_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12285_ net2562 _06887_ vssd1 vssd1 vccd1 vccd1 _06889_ sky130_fd_sc_hd__nand2_1
XFILLER_84_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08729__C1 net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11236_ net529 _06035_ net546 vssd1 vssd1 vccd1 vccd1 _06673_ sky130_fd_sc_hd__and3_1
X_11167_ net491 _06473_ _06643_ net299 net3792 vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__a32o_1
XFILLER_122_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10118_ _05740_ _05742_ _05755_ _05736_ vssd1 vssd1 vccd1 vccd1 _05756_ sky130_fd_sc_hd__o211a_1
X_13895__65 clknet_leaf_182_clk vssd1 vssd1 vccd1 vccd1 net1534 sky130_fd_sc_hd__inv_2
XFILLER_95_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15975_ net2309 _02185_ net1203 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[775\]
+ sky130_fd_sc_hd__dfrtp_1
X_11098_ net460 net526 _05810_ vssd1 vssd1 vccd1 vccd1 _06607_ sky130_fd_sc_hd__and3_1
XFILLER_76_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10049_ _05519_ _05683_ _05615_ vssd1 vssd1 vccd1 vccd1 _05688_ sky130_fd_sc_hd__or3b_1
X_14926_ clknet_leaf_31_clk _01172_ net1152 vssd1 vssd1 vccd1 vccd1 top.CPU.alu.program_counter\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_76_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10303__A2 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14165__335 clknet_leaf_170_clk vssd1 vssd1 vccd1 vccd1 net1804 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_82_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13808_ net3770 net333 net326 top.CPU.data_out\[10\] vssd1 vssd1 vccd1 vccd1 _02688_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09457__B1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12056__A2 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11281__B _06570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13739_ top.SPI.timem\[17\] _03077_ net3874 vssd1 vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__a21oi_1
XFILLER_149_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16527_ clknet_leaf_100_clk _02689_ net1257 vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__dfrtp_1
XFILLER_91_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11803__A2 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14206__376 clknet_leaf_154_clk vssd1 vssd1 vccd1 vccd1 net1845 sky130_fd_sc_hd__inv_2
XFILLER_149_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16458_ clknet_leaf_87_clk _02620_ net1271 vssd1 vssd1 vccd1 vccd1 top.SPI.timem\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15409_ net1743 _01619_ net1191 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[209\]
+ sky130_fd_sc_hd__dfrtp_1
X_16389_ clknet_leaf_87_clk _00069_ net1264 vssd1 vssd1 vccd1 vccd1 top.SPI.register\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_117_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_83_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11567__A1 _06678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09178__S net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_152_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12543__D _06450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09901_ _05536_ _05537_ _05539_ vssd1 vssd1 vccd1 vccd1 _05540_ sky130_fd_sc_hd__a21bo_1
XFILLER_132_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13495__Y _02966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_98_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout505 _05679_ vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_130_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08196__B1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13428__S net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout516 net523 vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__clkbuf_4
XFILLER_141_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09832_ top.CPU.registers.data\[154\] net1000 _05470_ vssd1 vssd1 vccd1 vccd1 _05471_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__09393__C1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout527 net533 vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__buf_2
XFILLER_99_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_171_Right_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout538 net539 vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_141_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout549 net550 vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__clkbuf_2
XFILLER_112_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09763_ top.CPU.registers.data\[315\] top.CPU.registers.data\[283\] net991 vssd1
+ vssd1 vccd1 vccd1 _05402_ sky130_fd_sc_hd__mux2_1
XFILLER_101_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10360__B net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout283_A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_21_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08714_ top.CPU.registers.data\[77\] net1312 net843 top.CPU.registers.data\[109\]
+ net762 vssd1 vssd1 vccd1 vccd1 _04353_ sky130_fd_sc_hd__a221o_1
XFILLER_39_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08499__A1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13492__A1 _04855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09694_ top.CPU.registers.data\[313\] top.CPU.registers.data\[281\] net1001 vssd1
+ vssd1 vccd1 vccd1 _05333_ sky130_fd_sc_hd__mux2_1
XFILLER_55_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11175__C _06648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08645_ top.CPU.registers.data\[334\] net1322 net853 top.CPU.registers.data\[366\]
+ net770 vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_156_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12568__A _06147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10845__A3 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout548_A net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout169_X net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1192_A net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08576_ top.CPU.registers.data\[463\] net1315 net846 top.CPU.registers.data\[495\]
+ net717 vssd1 vssd1 vccd1 vccd1 _04215_ sky130_fd_sc_hd__a221o_1
XANTENNA__13244__B2 _02803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10359__Y _05990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_36_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13835__5 clknet_leaf_135_clk vssd1 vssd1 vccd1 vccd1 net1474 sky130_fd_sc_hd__inv_2
XANTENNA__09999__A1 _04430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07527_ _03152_ net1045 _03159_ _03163_ vssd1 vssd1 vccd1 vccd1 _03166_ sky130_fd_sc_hd__and4b_1
XANTENNA__13795__A2 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout715_A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07458_ top.CPU.registers.data_out_r2_prev\[31\] vssd1 vssd1 vccd1 vccd1 _03098_
+ sky130_fd_sc_hd__inv_2
XFILLER_23_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15507__RESET_B net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout503_X net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09128_ top.CPU.registers.data\[583\] net1296 net1016 top.CPU.registers.data\[615\]
+ net938 vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__a221o_1
XFILLER_157_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09059_ net1034 net449 _04667_ vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__a21oi_2
XANTENNA__08974__A2 net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12070_ net565 net362 _06613_ _06804_ _06803_ vssd1 vssd1 vccd1 vccd1 _01529_ sky130_fd_sc_hd__a41o_1
XFILLER_1_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout872_X net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold570 top.CPU.registers.data\[192\] vssd1 vssd1 vccd1 vccd1 net3127 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold581 top.CPU.registers.data\[690\] vssd1 vssd1 vccd1 vccd1 net3138 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08187__B1 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold592 top.CPU.registers.data\[474\] vssd1 vssd1 vccd1 vccd1 net3149 sky130_fd_sc_hd__dlygate4sd3_1
X_11021_ net528 _06567_ vssd1 vssd1 vccd1 vccd1 _06568_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_38_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_109_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12242__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10551__A net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11730__A1 _06577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09136__C1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15760_ net2094 _01970_ net1157 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[560\]
+ sky130_fd_sc_hd__dfrtp_1
X_12972_ _07407_ top.I2C.bit_timer_state\[0\] _07405_ vssd1 vssd1 vccd1 vccd1 _01197_
+ sky130_fd_sc_hd__and3b_1
XANTENNA__12286__A2 _06887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14149__319 clknet_leaf_112_clk vssd1 vssd1 vccd1 vccd1 net1788 sky130_fd_sc_hd__inv_2
Xhold1270 top.CPU.registers.data\[962\] vssd1 vssd1 vccd1 vccd1 net3827 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input11_A DAT_I[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1281 top.I2C.inter_received vssd1 vssd1 vccd1 vccd1 net3838 sky130_fd_sc_hd__dlygate4sd3_1
X_11923_ net3718 net184 net341 _06293_ vssd1 vssd1 vccd1 vccd1 _01643_ sky130_fd_sc_hd__a22o_1
XANTENNA__07698__C1 net1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15691_ net2025 _01901_ net1057 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[491\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11494__B1 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1292 top.CPU.registers.data\[48\] vssd1 vssd1 vccd1 vccd1 net3849 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09439__B1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11854_ _06689_ net234 net152 net2677 vssd1 vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__a22o_1
XFILLER_60_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_831 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10805_ net382 _06378_ vssd1 vssd1 vccd1 vccd1 _06415_ sky130_fd_sc_hd__and2_1
XANTENNA__13786__A2 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11785_ _06631_ net199 net160 net3076 vssd1 vssd1 vccd1 vccd1 _01770_ sky130_fd_sc_hd__a22o_1
XFILLER_159_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13524_ top.CPU.data_out\[20\] net589 net339 _02982_ vssd1 vssd1 vccd1 vccd1 _02518_
+ sky130_fd_sc_hd__o22a_1
X_16312_ clknet_leaf_96_clk _02521_ net1247 vssd1 vssd1 vccd1 vccd1 top.CPU.data_out\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09787__A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10736_ _04923_ _05274_ _04862_ vssd1 vssd1 vccd1 vccd1 _06350_ sky130_fd_sc_hd__o21a_1
XFILLER_13_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08662__A1 net1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12925__B _03576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16243_ clknet_leaf_33_clk _02453_ net1123 vssd1 vssd1 vccd1 vccd1 top.CPU.control_unit.instruction\[19\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_173_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13538__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13455_ net1399 net872 _02897_ net419 vssd1 vssd1 vccd1 vccd1 _02949_ sky130_fd_sc_hd__a31o_1
X_10667_ _06282_ _06283_ _06277_ vssd1 vssd1 vccd1 vccd1 _06284_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_97_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12406_ _03120_ top.I2C.I2C_state\[10\] net2602 vssd1 vssd1 vccd1 vccd1 _00027_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_97_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16174_ net2508 _02384_ net1107 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[974\]
+ sky130_fd_sc_hd__dfrtp_1
X_13386_ _02830_ _02907_ vssd1 vssd1 vccd1 vccd1 _02908_ sky130_fd_sc_hd__nor2_1
XANTENNA__09611__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12210__A2 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10598_ _06177_ _06217_ net306 vssd1 vssd1 vccd1 vccd1 _06218_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15125_ clknet_leaf_57_clk net2560 net1144 vssd1 vssd1 vccd1 vccd1 top.CPU.done sky130_fd_sc_hd__dfstp_2
XFILLER_154_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14550__720 clknet_leaf_175_clk vssd1 vssd1 vccd1 vccd1 net2189 sky130_fd_sc_hd__inv_2
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__buf_2
X_12337_ net2597 _05018_ net1208 vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__mux2_1
Xoutput119 net119 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_58_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15056_ clknet_leaf_59_clk _00060_ net1134 vssd1 vssd1 vccd1 vccd1 top.I2C.output_state\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_75_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12268_ net2936 net149 net433 vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__mux2_1
XANTENNA__10509__C1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08178__B1 net1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09375__C1 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11219_ net493 net468 _06664_ net295 net2846 vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__a32o_1
X_12199_ net361 _06742_ _06866_ net169 net3774 vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__a32o_1
XANTENNA__10524__A2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput90 net90 vssd1 vssd1 vccd1 vccd1 DAT_O[2] sky130_fd_sc_hd__buf_2
XANTENNA__09027__A _04634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09127__C1 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15958_ net2292 _02168_ net1227 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[758\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_83_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11485__B1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15889_ net2223 _02099_ net1192 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[689\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11292__A net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08430_ net796 _04063_ _04064_ net725 vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__o211a_1
XFILLER_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08361_ top.CPU.registers.data\[978\] net1317 net848 top.CPU.registers.data\[1010\]
+ net718 vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__a221o_1
XANTENNA__08102__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07769__X _03408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08292_ top.CPU.registers.data\[243\] net1393 net826 top.CPU.registers.data\[211\]
+ net774 vssd1 vssd1 vccd1 vccd1 _03931_ sky130_fd_sc_hd__a221o_1
XANTENNA__09850__B1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15600__RESET_B net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10636__A net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09602__B1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12201__A2 _06796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14293__463 clknet_leaf_172_clk vssd1 vssd1 vccd1 vccd1 net1932 sky130_fd_sc_hd__inv_2
XFILLER_160_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10763__A2 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08540__S net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08169__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09366__C1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout498_A net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout302 _06604_ vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout313 net314 vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__buf_4
XANTENNA__10371__A net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout324 net325 vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__clkbuf_8
Xfanout335 _03047_ vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1205_A net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10802__C net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout346 _06771_ vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input3_A DAT_I[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout357 net359 vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__buf_8
XFILLER_59_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09815_ top.CPU.registers.data\[602\] net1337 net867 top.CPU.registers.data\[634\]
+ net758 vssd1 vssd1 vccd1 vccd1 _05454_ sky130_fd_sc_hd__a221o_1
XANTENNA__11186__B net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout368 net369 vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__buf_8
Xfanout379 net380 vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout665_A net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09118__C1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout286_X net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09746_ net797 _05383_ _05384_ net727 vssd1 vssd1 vccd1 vccd1 _05385_ sky130_fd_sc_hd__o211a_1
XANTENNA__13465__A1 net1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09677_ top.CPU.registers.data_out_r1_prev\[25\] net876 _05311_ _05315_ net780 vssd1
+ vssd1 vccd1 vccd1 _05316_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout453_X net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout832_A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08628_ top.CPU.registers.data\[814\] top.CPU.registers.data\[782\] net819 vssd1
+ vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__mux2_1
XANTENNA__07695__A2 _03154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08559_ top.CPU.registers.data\[47\] top.CPU.registers.data\[15\] net811 vssd1 vssd1
+ vccd1 vccd1 _04198_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout620_X net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1362_X net1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12585__X _07089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11779__A1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout718_X net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11570_ _06681_ net262 net247 net2881 vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__a22o_1
XANTENNA__08715__S net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10521_ _04191_ _05669_ _06131_ _06133_ vssd1 vssd1 vccd1 vccd1 _06145_ sky130_fd_sc_hd__o22a_1
XANTENNA__07852__C1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14534__704 clknet_leaf_126_clk vssd1 vssd1 vccd1 vccd1 net2173 sky130_fd_sc_hd__inv_2
XFILLER_109_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13240_ net892 top.I2C.data_out\[15\] _02789_ vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__mux2_1
X_10452_ _05860_ _06044_ _06071_ net406 vssd1 vssd1 vccd1 vccd1 _06079_ sky130_fd_sc_hd__o22a_1
XFILLER_155_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10203__A1 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13171_ top.I2C.within_byte_counter_reading\[2\] _02754_ _02755_ _02752_ vssd1 vssd1
+ vccd1 vccd1 _01336_ sky130_fd_sc_hd__a22o_1
XANTENNA__11400__B1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10383_ _03719_ _05965_ _03789_ vssd1 vssd1 vccd1 vccd1 _06012_ sky130_fd_sc_hd__a21oi_1
XFILLER_124_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12122_ net136 net363 net356 net174 top.CPU.registers.data\[91\] vssd1 vssd1 vccd1
+ vccd1 _06829_ sky130_fd_sc_hd__a32o_1
XANTENNA__09546__S net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13576__B _06251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09357__C1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12053_ _06605_ net351 net179 net3728 vssd1 vssd1 vccd1 vccd1 _01537_ sky130_fd_sc_hd__a22o_1
XANTENNA__10281__A net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12900__A0 top.CPU.alu.program_counter\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11004_ _06291_ net540 vssd1 vssd1 vccd1 vccd1 _06557_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_53_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11096__B net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout880 _03198_ vssd1 vssd1 vccd1 vccd1 net880 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout891 net893 vssd1 vssd1 vccd1 vccd1 net891 sky130_fd_sc_hd__buf_2
X_15812_ net2146 _02022_ net1186 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[612\]
+ sky130_fd_sc_hd__dfrtp_1
X_13865__35 clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 net1504 sky130_fd_sc_hd__inv_2
XFILLER_19_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09281__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11467__B1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09124__A2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12955_ top.CPU.alu.program_counter\[31\] net1363 vssd1 vssd1 vccd1 vccd1 _07394_
+ sky130_fd_sc_hd__and2b_1
X_15743_ net2077 _01953_ net1224 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[543\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08332__B1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11906_ net3673 net186 net352 _05908_ vssd1 vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__a22o_1
XFILLER_18_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12886_ _07328_ _07330_ vssd1 vssd1 vccd1 vccd1 _07332_ sky130_fd_sc_hd__nor2_1
XANTENNA__08883__A1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15674_ net2008 _01884_ net1252 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[474\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11219__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11837_ net470 _06668_ net242 net154 net3054 vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_16_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10518__A1_N net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11768_ net470 _06611_ net241 net163 net3068 vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__a32o_1
XFILLER_13_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12655__B _05087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14924__Q top.CPU.alu.program_counter\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13507_ top.CPU.data_out\[12\] net587 _02969_ _02973_ vssd1 vssd1 vccd1 vccd1 _02510_
+ sky130_fd_sc_hd__o22a_1
XFILLER_9_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10719_ _06333_ vssd1 vssd1 vccd1 vccd1 _06334_ sky130_fd_sc_hd__inv_2
XFILLER_147_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07843__C1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11699_ _06530_ net207 net421 net2794 vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__a22o_1
XANTENNA__10993__A2 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14277__447 clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 net1916 sky130_fd_sc_hd__inv_2
X_13438_ net4008 _02940_ net121 vssd1 vssd1 vccd1 vccd1 _02474_ sky130_fd_sc_hd__mux2_1
X_16226_ clknet_leaf_29_clk _02436_ net1153 vssd1 vssd1 vccd1 vccd1 top.CPU.control_unit.instruction\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_77_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12195__A1 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08399__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08938__A2 net1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16157_ net2491 _02367_ net1119 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[957\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_142_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13369_ top.CPU.control_unit.instruction\[16\] _02895_ net671 vssd1 vssd1 vccd1 vccd1
+ _02450_ sky130_fd_sc_hd__mux2_1
XANTENNA__12671__A top.CPU.alu.program_counter\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14021__191 clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 net1660 sky130_fd_sc_hd__inv_2
XFILLER_142_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09456__S net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15108_ net1490 _01321_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r2_prev\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_14318__488 clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 net1957 sky130_fd_sc_hd__inv_2
X_16088_ net2422 _02298_ net1148 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[888\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_138_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10903__B net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11287__A net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15039_ clknet_leaf_91_clk _01284_ net1269 vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__dfrtp_1
X_07930_ top.CPU.registers.data\[284\] net996 _03568_ vssd1 vssd1 vccd1 vccd1 _03569_
+ sky130_fd_sc_hd__a21o_1
XFILLER_123_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08020__C1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07861_ top.CPU.registers.data\[413\] net980 _03499_ vssd1 vssd1 vccd1 vccd1 _03500_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_147_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09600_ top.CPU.registers.data\[64\] net1313 net846 top.CPU.registers.data\[96\]
+ net766 vssd1 vssd1 vccd1 vccd1 _05239_ sky130_fd_sc_hd__a221o_1
XANTENNA__08571__B1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11170__A2 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07792_ net628 _03427_ _03428_ net614 vssd1 vssd1 vccd1 vccd1 _03431_ sky130_fd_sc_hd__a31o_1
XANTENNA__09191__S net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09531_ top.CPU.registers.data\[545\] top.CPU.registers.data\[513\] net837 vssd1
+ vssd1 vccd1 vccd1 _05170_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_108_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08323__B1 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09462_ net707 _05099_ _05100_ vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__or3_1
XFILLER_36_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08413_ _04020_ _04051_ vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__and2_1
X_09393_ top.CPU.registers.data\[451\] net1328 net859 top.CPU.registers.data\[483\]
+ net775 vssd1 vssd1 vccd1 vccd1 _05032_ sky130_fd_sc_hd__a221o_1
XFILLER_40_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout246_A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08344_ net955 _03961_ _03980_ net606 vssd1 vssd1 vccd1 vccd1 _03983_ sky130_fd_sc_hd__a211o_1
XANTENNA__08087__C1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09823__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09220__A _04829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07659__B _03252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11630__B1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08275_ net947 _03899_ _03900_ _03913_ net608 vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__a311o_1
XANTENNA_fanout413_A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13383__A0 net1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12186__A1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout201_X net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1322_A net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08270__S net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_167_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11197__A net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1108 net1109 vssd1 vssd1 vccd1 vccd1 net1108 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1110_X net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout121 net122 vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_35_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1119 net1122 vssd1 vssd1 vccd1 vccd1 net1119 sky130_fd_sc_hd__clkbuf_4
XFILLER_87_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout132 _06085_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__buf_2
XFILLER_102_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09354__A2 net1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout143 _06173_ vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__buf_2
XANTENNA__11697__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout154 net155 vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__buf_6
XANTENNA_fanout570_X net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout165 _06757_ vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout176 _06795_ vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__clkbuf_8
Xfanout187 _06769_ vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__clkbuf_8
Xfanout198 net202 vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__clkbuf_4
XFILLER_75_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09729_ top.CPU.registers.data\[571\] top.CPU.registers.data\[539\] net828 vssd1
+ vssd1 vccd1 vccd1 _05368_ sky130_fd_sc_hd__mux2_1
XFILLER_28_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout835_X net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08314__B1 net1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09511__C1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12740_ _07193_ _07199_ net127 vssd1 vssd1 vccd1 vccd1 _07200_ sky130_fd_sc_hd__mux2_1
XFILLER_28_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10121__B1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12671_ top.CPU.alu.program_counter\[4\] _04955_ vssd1 vssd1 vccd1 vccd1 _07137_
+ sky130_fd_sc_hd__nand2_1
XFILLER_70_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12756__A top.CPU.alu.program_counter\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13204__X _02782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11622_ _06373_ net3020 net212 vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__mux2_1
XANTENNA__08617__A1 net1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15390_ net1724 _01600_ net1239 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[190\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12475__B _04122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10424__A1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11621__A0 _06354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11553_ net567 net493 _06666_ net249 net2662 vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__a32o_1
XANTENNA__07825__C1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10504_ _05290_ net446 vssd1 vssd1 vccd1 vccd1 _06128_ sky130_fd_sc_hd__and2_1
XFILLER_11_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14005__175 clknet_leaf_176_clk vssd1 vssd1 vccd1 vccd1 net1644 sky130_fd_sc_hd__inv_2
X_11484_ net496 net475 _06614_ net256 net3151 vssd1 vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_94_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07840__A2 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16011_ net2345 _02221_ net1064 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[811\]
+ sky130_fd_sc_hd__dfrtp_1
X_13223_ _02774_ _02792_ vssd1 vssd1 vccd1 vccd1 _02795_ sky130_fd_sc_hd__nand2_1
Xwire599 _06931_ vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__clkbuf_2
XFILLER_143_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10435_ _05584_ _06061_ _05297_ vssd1 vssd1 vccd1 vccd1 _06062_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12491__A _04763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13154_ _06895_ _06907_ _02743_ _06891_ vssd1 vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__o22a_1
XFILLER_128_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09593__A2 net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10366_ _03921_ net509 net504 _03919_ _05995_ vssd1 vssd1 vccd1 vccd1 _05996_ sky130_fd_sc_hd__o221a_1
XFILLER_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_29_Left_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12105_ net3987 net653 _06820_ vssd1 vssd1 vccd1 vccd1 _01510_ sky130_fd_sc_hd__o21a_1
XFILLER_111_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13085_ top.CPU.data_out\[20\] net3215 net559 vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__mux2_1
X_10297_ _05367_ _05596_ vssd1 vssd1 vccd1 vccd1 _05930_ sky130_fd_sc_hd__xnor2_1
X_12036_ _06589_ _06779_ _06781_ net3030 vssd1 vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__a22o_1
XANTENNA__08002__C1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11688__B1 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11152__A2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14662__832 clknet_leaf_123_clk vssd1 vssd1 vccd1 vccd1 net2301 sky130_fd_sc_hd__inv_2
XFILLER_77_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13429__A1 _02858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12453__A2_N _03439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08305__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09502__C1 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10112__A0 _03544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15726_ net2060 _01936_ net1193 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[526\]
+ sky130_fd_sc_hd__dfrtp_1
X_12938_ _07377_ _07378_ vssd1 vssd1 vccd1 vccd1 _07379_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11273__C net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08856__A1 net1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14703__873 clknet_leaf_179_clk vssd1 vssd1 vccd1 vccd1 net2342 sky130_fd_sc_hd__inv_2
XFILLER_61_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_38_Left_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11860__B1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15657_ net1991 _01867_ net1056 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[457\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ top.CPU.alu.program_counter\[22\] _07316_ net1359 vssd1 vssd1 vccd1 vccd1
+ _01185_ sky130_fd_sc_hd__mux2_1
XFILLER_33_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08355__S net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09805__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15588_ net1922 _01798_ net1221 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[388\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10457__Y _06084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10415__A1 _03242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11612__A0 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09281__A1 _04919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10966__A2 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08060_ net674 _03694_ _03695_ _03698_ net610 vssd1 vssd1 vccd1 vccd1 _03699_ sky130_fd_sc_hd__a311o_1
XFILLER_135_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13365__A0 net1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09569__C1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13497__A _04726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16209_ net2543 _02419_ net1176 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[1009\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07766__Y _03405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Left_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08241__C1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10633__B _06251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11391__A2 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08962_ _04600_ vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__inv_2
XANTENNA__09336__A2 net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07913_ net961 _03546_ _03548_ _03551_ vssd1 vssd1 vccd1 vccd1 _03552_ sky130_fd_sc_hd__a31o_1
XFILLER_25_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11679__B1 net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08893_ top.CPU.alu.program_counter\[11\] _04531_ net1033 vssd1 vssd1 vccd1 vccd1
+ _04532_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_127_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12340__A1 _05226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout196_A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07844_ top.CPU.registers.data\[253\] net1379 net979 top.CPU.registers.data\[221\]
+ net905 vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_162_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12891__A2 _07322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07775_ _03412_ _03413_ net621 vssd1 vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout363_A net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_56_Left_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09514_ _05145_ _05146_ net681 vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_140_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09445_ _05070_ _05071_ _05076_ _05083_ vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__a22o_2
XANTENNA__11851__B1 net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout151_X net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout530_A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1272_A net1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout628_A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout249_X net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09376_ net939 _04994_ _04995_ net956 vssd1 vssd1 vccd1 vccd1 _05015_ sky130_fd_sc_hd__o211a_1
X_08327_ top.CPU.registers.data\[51\] top.CPU.registers.data\[19\] net988 vssd1 vssd1
+ vccd1 vccd1 _03966_ sky130_fd_sc_hd__mux2_1
XFILLER_166_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07807__C1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09272__A1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout416_X net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10957__A2 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08258_ top.CPU.registers.data\[54\] top.CPU.registers.data\[22\] net1002 vssd1 vssd1
+ vccd1 vccd1 _03897_ sky130_fd_sc_hd__mux2_1
XANTENNA__08480__C1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout997_A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_65_Left_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09024__A1 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10824__A net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08189_ top.CPU.registers.data\[87\] net1295 net1014 top.CPU.registers.data\[119\]
+ net937 vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1325_X net1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10220_ net445 _05599_ _05854_ vssd1 vssd1 vccd1 vccd1 _05855_ sky130_fd_sc_hd__o21bai_1
XFILLER_106_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10151_ _05637_ _05645_ net306 vssd1 vssd1 vccd1 vccd1 _05788_ sky130_fd_sc_hd__mux2_1
XANTENNA__10590__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07692__X _03331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14646__816 clknet_leaf_181_clk vssd1 vssd1 vccd1 vccd1 net2285 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_50_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10082_ _05718_ _05719_ net383 vssd1 vssd1 vccd1 vccd1 _05720_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout952_X net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12250__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11685__A3 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09125__A _04763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13772_ net31 net1049 net884 net3542 vssd1 vssd1 vccd1 vccd1 _02653_ sky130_fd_sc_hd__o22a_1
XANTENNA__12095__B1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11093__C net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10984_ net519 net442 net140 net545 vssd1 vssd1 vccd1 vccd1 _06545_ sky130_fd_sc_hd__and4_1
X_15511_ net1845 _01721_ net1181 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[311\]
+ sky130_fd_sc_hd__dfrtp_1
X_12723_ top.CPU.alu.program_counter\[9\] _04660_ vssd1 vssd1 vccd1 vccd1 _07184_
+ sky130_fd_sc_hd__or2_1
XANTENNA__11842__B1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16491_ clknet_leaf_40_clk _02653_ net1115 vssd1 vssd1 vccd1 vccd1 top.mmio.mem_data_i\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12654_ top.CPU.alu.program_counter\[2\] _05087_ vssd1 vssd1 vccd1 vccd1 _07122_
+ sky130_fd_sc_hd__and2_1
X_15442_ net1776 _01652_ net1101 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[242\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08175__S net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11605_ _06487_ net428 net208 net215 net2918 vssd1 vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__a32o_1
XFILLER_169_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14899__1069 clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 net2538 sky130_fd_sc_hd__inv_2
X_12585_ _03130_ net598 vssd1 vssd1 vccd1 vccd1 _07089_ sky130_fd_sc_hd__and2_2
X_15373_ net1707 _01583_ net1067 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[173\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09795__A _05399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11536_ net478 _06290_ net354 net250 net3230 vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_61_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11070__B2 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07813__A2 net1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11467_ net3665 net264 net259 _06594_ vssd1 vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__a22o_1
XFILLER_171_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13206_ net3824 _02779_ _02783_ _02773_ vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__a22o_1
X_10418_ net411 _06045_ net224 vssd1 vssd1 vccd1 vccd1 _06046_ sky130_fd_sc_hd__a21o_1
XANTENNA__09566__A2 net1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11398_ _06526_ net282 net269 net2668 vssd1 vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__a22o_1
XANTENNA__07577__A1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11373__A2 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08774__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13137_ net2763 _02737_ _02734_ vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__mux2_1
XFILLER_125_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10349_ _03858_ _05670_ net506 _03823_ vssd1 vssd1 vccd1 vccd1 _05980_ sky130_fd_sc_hd__a22o_1
XFILLER_124_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14092__262 clknet_leaf_188_clk vssd1 vssd1 vccd1 vccd1 net1731 sky130_fd_sc_hd__inv_2
XFILLER_140_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13764__B net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13068_ top.CPU.data_out\[3\] net2683 net558 vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__mux2_1
X_14389__559 clknet_leaf_173_clk vssd1 vssd1 vccd1 vccd1 net2028 sky130_fd_sc_hd__inv_2
XANTENNA__11125__A2 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12322__A1 _04048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12019_ _05960_ net150 _06786_ vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__o21ai_1
XFILLER_94_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12873__A2 _03916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11676__A3 net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10884__A1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07560_ net1408 _03154_ _03155_ vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_85_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15709_ net2043 _01919_ net1113 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[509\]
+ sky130_fd_sc_hd__dfrtp_1
X_07491_ net1 vssd1 vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__inv_2
XANTENNA__11833__B1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_1028 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09230_ top.CPU.registers.data\[901\] net1310 net841 top.CPU.registers.data\[933\]
+ net690 vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__a221o_1
XFILLER_167_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09161_ top.CPU.registers.data\[230\] net1389 net814 top.CPU.registers.data\[198\]
+ net767 vssd1 vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__a221o_1
X_14790__960 clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 net2429 sky130_fd_sc_hd__inv_2
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10939__A2 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08112_ top.CPU.registers.data\[981\] net1329 net860 top.CPU.registers.data\[1013\]
+ net776 vssd1 vssd1 vccd1 vccd1 _03751_ sky130_fd_sc_hd__a221o_1
XFILLER_174_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09092_ _04698_ _04729_ vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__or2_1
XANTENNA__11061__B2 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08462__C1 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08043_ _03679_ _03680_ _03681_ _03666_ vssd1 vssd1 vccd1 vccd1 _03682_ sky130_fd_sc_hd__a211oi_2
XFILLER_147_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09006__A1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold900 top.CPU.registers.data\[24\] vssd1 vssd1 vccd1 vccd1 net3457 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_174_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold911 top.I2C.data_out\[25\] vssd1 vssd1 vccd1 vccd1 net3468 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12562__C _06124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold922 top.CPU.registers.data\[671\] vssd1 vssd1 vccd1 vccd1 net3479 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout209_A net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14333__503 clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 net1972 sky130_fd_sc_hd__inv_2
X_13997__167 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 net1636 sky130_fd_sc_hd__inv_2
XANTENNA__12010__A0 _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold933 top.CPU.registers.data\[1011\] vssd1 vssd1 vccd1 vccd1 net3490 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold944 top.CPU.registers.data\[680\] vssd1 vssd1 vccd1 vccd1 net3501 sky130_fd_sc_hd__dlygate4sd3_1
Xhold955 top.CPU.registers.data\[953\] vssd1 vssd1 vccd1 vccd1 net3512 sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 top.CPU.registers.data\[741\] vssd1 vssd1 vccd1 vccd1 net3523 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold977 top.CPU.registers.data\[848\] vssd1 vssd1 vccd1 vccd1 net3534 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_164_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09994_ _04532_ _04567_ net378 vssd1 vssd1 vccd1 vccd1 _05633_ sky130_fd_sc_hd__mux2_1
Xhold988 top.mmio.mem_data_i\[6\] vssd1 vssd1 vccd1 vccd1 net3545 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1020_A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold999 net76 vssd1 vssd1 vccd1 vccd1 net3556 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10572__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1118_A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08945_ top.CPU.registers.data\[714\] net1374 net971 top.CPU.registers.data\[746\]
+ net928 vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout480_A net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12313__A1 _05428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout578_A net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout199_X net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09714__C1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08876_ top.CPU.registers.data\[459\] net1311 net842 top.CPU.registers.data\[491\]
+ net762 vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__a221o_1
XANTENNA__09190__A0 top.CPU.alu.program_counter\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11194__B net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07827_ top.CPU.registers.data\[477\] net1318 net849 top.CPU.registers.data\[509\]
+ net768 vssd1 vssd1 vccd1 vccd1 _03466_ sky130_fd_sc_hd__a221o_1
XANTENNA__10875__B2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout366_X net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout745_A net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07758_ top.CPU.registers.data\[94\] net1333 net864 top.CPU.registers.data\[126\]
+ net781 vssd1 vssd1 vccd1 vccd1 _03397_ sky130_fd_sc_hd__a221o_1
XFILLER_37_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07689_ _03285_ net632 _03306_ _03326_ _03327_ vssd1 vssd1 vccd1 vccd1 _03328_ sky130_fd_sc_hd__a311o_1
XANTENNA__10378__X _06008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout912_A net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout533_X net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1275_X net1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10819__A net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09428_ top.CPU.registers.data\[162\] net1383 net986 top.CPU.registers.data\[130\]
+ net677 vssd1 vssd1 vccd1 vccd1 _05067_ sky130_fd_sc_hd__a221o_1
XFILLER_44_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09359_ top.CPU.registers.data\[323\] net1297 net1018 top.CPU.registers.data\[355\]
+ net939 vssd1 vssd1 vccd1 vccd1 _04998_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout700_X net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08048__A2 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13941__111 clknet_leaf_174_clk vssd1 vssd1 vccd1 vccd1 net1580 sky130_fd_sc_hd__inv_2
X_12370_ _06905_ _06908_ _06909_ _06907_ vssd1 vssd1 vccd1 vccd1 _00042_ sky130_fd_sc_hd__a31o_1
XANTENNA__11052__B2 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11321_ net3207 net290 net358 _06354_ vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__a22o_1
XFILLER_5_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12245__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08205__C1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11252_ net486 net461 _06681_ net293 net2658 vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__a32o_1
XANTENNA__12001__B1 net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14076__246 clknet_leaf_140_clk vssd1 vssd1 vccd1 vccd1 net1715 sky130_fd_sc_hd__inv_2
XANTENNA__10273__B _05906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12552__A1 top.CPU.done vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10203_ net385 _05730_ _05838_ vssd1 vssd1 vccd1 vccd1 _05839_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11355__A2 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11183_ _06057_ net3730 net298 vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__mux2_1
XFILLER_79_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10134_ net1407 net576 net522 net137 vssd1 vssd1 vccd1 vccd1 _05772_ sky130_fd_sc_hd__and4_1
XFILLER_122_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15991_ net2325 _02201_ net1173 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[791\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12304__A1 _04986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14117__287 clknet_leaf_112_clk vssd1 vssd1 vccd1 vccd1 net1756 sky130_fd_sc_hd__inv_2
XANTENNA__11107__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08508__B1 net1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10195__A2_N net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13076__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14942_ clknet_leaf_66_clk _01188_ net1165 vssd1 vssd1 vccd1 vccd1 top.CPU.alu.program_counter\[25\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09126__Y _04765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10065_ net372 _05266_ vssd1 vssd1 vccd1 vccd1 _05703_ sky130_fd_sc_hd__nand2_1
XFILLER_76_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09181__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16612_ net1347 vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_1
X_13824_ net3110 net337 net329 top.CPU.data_out\[26\] vssd1 vssd1 vccd1 vccd1 _02704_
+ sky130_fd_sc_hd__a22o_1
XFILLER_165_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13804__B2 top.CPU.data_out\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11815__A0 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16543_ clknet_leaf_91_clk net2811 net1270 vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__dfrtp_1
XFILLER_141_92 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10618__B2 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13755_ top.I2C.I2C_state\[16\] _03088_ vssd1 vssd1 vccd1 vccd1 _03089_ sky130_fd_sc_hd__nand2_1
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10967_ net516 _05962_ net544 vssd1 vssd1 vccd1 vccd1 _06535_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_63_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12706_ _07167_ _07168_ vssd1 vssd1 vccd1 vccd1 _07169_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_63_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16474_ clknet_leaf_88_clk _02636_ net1274 vssd1 vssd1 vccd1 vccd1 top.SPI.timem\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_14774__944 clknet_leaf_180_clk vssd1 vssd1 vccd1 vccd1 net2413 sky130_fd_sc_hd__inv_2
X_13686_ net2638 net336 vssd1 vssd1 vccd1 vccd1 _02614_ sky130_fd_sc_hd__and2_1
X_10898_ net488 net464 _06492_ net222 net3021 vssd1 vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_80_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15425_ net1759 _01635_ net1230 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[225\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12637_ top.I2C.output_state\[14\] net3698 vssd1 vssd1 vccd1 vccd1 _00010_ sky130_fd_sc_hd__and2_1
XANTENNA__09236__A1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12944__A top.CPU.alu.program_counter\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09729__S net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12568_ _06147_ _06228_ _06251_ _07072_ vssd1 vssd1 vccd1 vccd1 _07073_ sky130_fd_sc_hd__or4_1
XANTENNA__08444__C1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15356_ net1690 _01566_ net1236 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[156\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11043__B2 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14815__985 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 net2454 sky130_fd_sc_hd__inv_2
XANTENNA__08995__A0 top.CPU.alu.program_counter\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12663__B _05021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07798__A1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_152_Right_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11519_ net3525 net253 _06734_ _06483_ vssd1 vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__a22o_1
XFILLER_145_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12499_ _05019_ _05054_ _05085_ _05121_ _07002_ vssd1 vssd1 vccd1 vccd1 _07008_ sky130_fd_sc_hd__o221a_1
X_15287_ net1621 _01497_ net1185 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[87\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold207 top.CPU.registers.data\[163\] vssd1 vssd1 vccd1 vccd1 net2764 sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 top.SPI.parameters\[8\] vssd1 vssd1 vccd1 vccd1 net2775 sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 _01270_ vssd1 vssd1 vccd1 vccd1 net2786 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_160_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15696__RESET_B net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11346__A2 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08211__A2 net1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout709 _03212_ vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__buf_2
XFILLER_124_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13494__B _03200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10911__B net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08730_ net1283 _04367_ _04368_ vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__or3_1
XANTENNA__12846__A2 _03986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1280 net1282 vssd1 vssd1 vccd1 vccd1 net1280 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09172__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08661_ net1283 _04298_ _04299_ vssd1 vssd1 vccd1 vccd1 _04300_ sky130_fd_sc_hd__or3_1
Xfanout1291 net1292 vssd1 vssd1 vccd1 vccd1 net1291 sky130_fd_sc_hd__clkbuf_4
XFILLER_22_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07722__A1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07612_ net1279 _03158_ vssd1 vssd1 vccd1 vccd1 _03251_ sky130_fd_sc_hd__nand2_2
X_08592_ top.CPU.registers.data\[463\] net1375 net974 top.CPU.registers.data\[495\]
+ net1365 vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__o221a_1
XFILLER_54_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07543_ net1404 net661 vssd1 vssd1 vccd1 vccd1 _03182_ sky130_fd_sc_hd__nand2_1
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11282__B2 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07474_ net1368 vssd1 vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__inv_2
XANTENNA__08683__C1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13559__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09213_ top.CPU.registers.data\[454\] net1287 net1006 top.CPU.registers.data\[486\]
+ net904 vssd1 vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_157_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1068_A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09144_ top.CPU.registers.data\[455\] net1302 net1024 top.CPU.registers.data\[487\]
+ net920 vssd1 vssd1 vccd1 vccd1 _04783_ sky130_fd_sc_hd__a221o_1
XANTENNA__11034__A1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12231__B1 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11585__A2 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09075_ top.CPU.registers.data\[840\] net1376 net975 top.CPU.registers.data\[872\]
+ net1281 vssd1 vssd1 vccd1 vccd1 _04714_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_135_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10793__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08115__Y _03754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1235_A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08026_ net693 _03663_ _03664_ vssd1 vssd1 vccd1 vccd1 _03665_ sky130_fd_sc_hd__or3_1
Xhold730 top.CPU.registers.data\[457\] vssd1 vssd1 vccd1 vccd1 net3287 sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 top.CPU.registers.data\[723\] vssd1 vssd1 vccd1 vccd1 net3298 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout695_A net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08738__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11337__A2 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold752 top.CPU.registers.data\[364\] vssd1 vssd1 vccd1 vccd1 net3309 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold763 top.CPU.registers.data\[488\] vssd1 vssd1 vccd1 vccd1 net3320 sky130_fd_sc_hd__dlygate4sd3_1
Xhold774 top.CPU.registers.data\[727\] vssd1 vssd1 vccd1 vccd1 net3331 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10545__B1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold785 top.CPU.registers.data\[499\] vssd1 vssd1 vccd1 vccd1 net3342 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1023_X net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold796 top.CPU.registers.data\[145\] vssd1 vssd1 vccd1 vccd1 net3353 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09977_ _03285_ _03310_ net547 _03324_ vssd1 vssd1 vccd1 vccd1 _05616_ sky130_fd_sc_hd__a31oi_4
XANTENNA_fanout862_A _03203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout483_X net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08928_ net1034 _04566_ _04536_ vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__a21oi_4
X_14898__1068 clknet_leaf_201_clk vssd1 vssd1 vccd1 vccd1 net2537 sky130_fd_sc_hd__inv_2
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1430 top.CPU.registers.data\[100\] vssd1 vssd1 vccd1 vccd1 net3987 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1441 top.CPU.handler.state\[6\] vssd1 vssd1 vccd1 vccd1 net3998 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1452 top.CPU.registers.data\[68\] vssd1 vssd1 vccd1 vccd1 net4009 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout650_X net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08859_ top.CPU.registers.data_out_r2_prev\[11\] net688 vssd1 vssd1 vccd1 vccd1 _04498_
+ sky130_fd_sc_hd__nor2_1
Xhold1463 top.CPU.registers.data\[111\] vssd1 vssd1 vccd1 vccd1 net4020 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout748_X net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1392_X net1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11933__A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11870_ _06706_ net242 net191 net3901 vssd1 vssd1 vccd1 vccd1 _01692_ sky130_fd_sc_hd__a22o_1
X_14461__631 clknet_leaf_130_clk vssd1 vssd1 vccd1 vccd1 net2100 sky130_fd_sc_hd__inv_2
XFILLER_45_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_979 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09403__A net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10821_ net3693 net226 net316 _06430_ vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__a22o_1
X_14758__928 clknet_leaf_133_clk vssd1 vssd1 vccd1 vccd1 net2397 sky130_fd_sc_hd__inv_2
XANTENNA_fanout915_X net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10752_ net411 _06363_ _06364_ _06139_ vssd1 vssd1 vccd1 vccd1 _06365_ sky130_fd_sc_hd__a31o_1
X_13540_ net3772 net591 net340 _02990_ vssd1 vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__o22a_1
X_14502__672 clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 net2141 sky130_fd_sc_hd__inv_2
X_13471_ net1399 net872 _02918_ net418 vssd1 vssd1 vccd1 vccd1 _02957_ sky130_fd_sc_hd__a31o_1
XANTENNA__10836__X _06445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10683_ _06297_ _06298_ _06139_ vssd1 vssd1 vccd1 vccd1 _06299_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09218__A1 _04856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12422_ top.I2C.within_byte_counter_reading\[1\] top.I2C.within_byte_counter_reading\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06947_ sky130_fd_sc_hd__nand2_1
X_15210_ net1544 _01420_ net1094 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13579__B _06228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16190_ net2524 _02400_ net1204 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[990\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_154_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12483__B _03854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11576__A2 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15141_ clknet_leaf_47_clk _01351_ net1131 vssd1 vssd1 vccd1 vccd1 top.I2C.data_out\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_12353_ net898 _06898_ vssd1 vssd1 vccd1 vccd1 _00063_ sky130_fd_sc_hd__nor2_1
XFILLER_139_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08441__A2 net1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11304_ net3045 net291 net359 _06033_ vssd1 vssd1 vccd1 vccd1 _02199_ sky130_fd_sc_hd__a22o_1
X_15072_ clknet_leaf_52_clk _00050_ net1132 vssd1 vssd1 vccd1 vccd1 top.I2C.output_state\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_107_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12284_ net2589 _03888_ net1222 vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__mux2_1
XANTENNA__09077__S0 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12525__A1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11328__A2 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12525__B2 _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11235_ net2962 net295 _06672_ net318 vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__a22o_1
XFILLER_122_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08689__A _04294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11166_ _03189_ _06644_ vssd1 vssd1 vccd1 vccd1 _06645_ sky130_fd_sc_hd__or2_4
XANTENNA__07952__A1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10117_ net396 _05747_ _05751_ _05754_ vssd1 vssd1 vccd1 vccd1 _05755_ sky130_fd_sc_hd__a211o_1
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12004__A net1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15974_ net2308 _02184_ net1080 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[774\]
+ sky130_fd_sc_hd__dfrtp_1
X_11097_ net492 net468 _06606_ net304 net3290 vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__a32o_1
XFILLER_95_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10048_ _03321_ _05686_ net413 vssd1 vssd1 vccd1 vccd1 _05687_ sky130_fd_sc_hd__a21o_1
X_14925_ clknet_leaf_31_clk _01171_ net1152 vssd1 vssd1 vccd1 vccd1 top.CPU.alu.program_counter\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_64_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11500__A2 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold90 top.CPU.registers.data\[828\] vssd1 vssd1 vccd1 vccd1 net2647 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_35_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12658__B _05232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13789__B1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14927__Q top.CPU.alu.program_counter\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13807_ net3624 net333 net326 top.CPU.data_out\[9\] vssd1 vssd1 vccd1 vccd1 _02687_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_82_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11562__B _06731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10459__A net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11999_ _06568_ net348 net182 net2764 vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__a22o_1
XFILLER_17_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_11_Left_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16526_ clknet_leaf_100_clk _02688_ net1255 vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__dfrtp_1
X_13738_ net3996 _03077_ _03078_ vssd1 vssd1 vccd1 vccd1 _02636_ sky130_fd_sc_hd__o21a_1
XFILLER_31_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16457_ clknet_leaf_87_clk _02619_ net1271 vssd1 vssd1 vccd1 vccd1 top.SPI.timem\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09209__A1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13669_ net2837 net331 net330 top.CPU.addressnew\[2\] vssd1 vssd1 vccd1 vccd1 _02597_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13005__A2 _07429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08680__A2 net1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15408_ net1742 _01618_ net1156 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[208\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11016__B2 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16388_ clknet_leaf_87_clk _00073_ net1271 vssd1 vssd1 vccd1 vccd1 top.SPI.state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_157_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11567__A2 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15339_ net1673 _01549_ net1066 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[139\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10194__A net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09900_ _04364_ _04393_ _04396_ _05538_ vssd1 vssd1 vccd1 vccd1 _05539_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_113_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_20_Left_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout506 _05676_ vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_130_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire451_X net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09194__S net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09393__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09831_ top.CPU.registers.data\[186\] net1027 net921 vssd1 vssd1 vccd1 vccd1 _05470_
+ sky130_fd_sc_hd__a21o_1
Xfanout517 net518 vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__clkbuf_4
Xfanout528 net533 vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__buf_4
XANTENNA_clkload13_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout539 _06574_ vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__buf_4
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09762_ top.CPU.registers.data\[923\] net1298 net1018 top.CPU.registers.data\[955\]
+ net915 vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__a221o_1
XFILLER_6_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10360__C net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08713_ top.CPU.registers.data\[45\] top.CPU.registers.data\[13\] net808 vssd1 vssd1
+ vccd1 vccd1 _04352_ sky130_fd_sc_hd__mux2_1
X_09693_ net1036 _05330_ _05301_ vssd1 vssd1 vccd1 vccd1 _05332_ sky130_fd_sc_hd__a21oi_4
XFILLER_55_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14445__615 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 net2084 sky130_fd_sc_hd__inv_2
XANTENNA_fanout276_A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08644_ top.CPU.registers.data\[302\] top.CPU.registers.data\[270\] net819 vssd1
+ vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__mux2_1
XFILLER_55_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12568__B _06228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08575_ net788 _04209_ _04210_ _04213_ net641 vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__a311o_1
XANTENNA__09448__A1 top.CPU.control_unit.instruction\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_81_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07526_ top.CPU.control_unit.instruction\[0\] top.CPU.control_unit.instruction\[1\]
+ _03157_ vssd1 vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__and3_1
XANTENNA__10998__C_N _06253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07457_ top.CPU.registers.data_out_r1_prev\[31\] vssd1 vssd1 vccd1 vccd1 _03097_
+ sky130_fd_sc_hd__inv_2
XANTENNA_fanout231_X net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout610_A net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08671__A2 net1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout329_X net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout708_A net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09127_ top.CPU.registers.data\[743\] net1383 net988 top.CPU.registers.data\[711\]
+ net913 vssd1 vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__a221o_1
XFILLER_148_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09620__A1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09081__C1 net1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08423__A2 net1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09058_ _04696_ vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__inv_2
XFILLER_68_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08009_ _03613_ _03647_ vssd1 vssd1 vccd1 vccd1 _03648_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout698_X net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold560 top.I2C.output_state\[27\] vssd1 vssd1 vccd1 vccd1 net3117 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10518__B1 _06141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1405_X net1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09384__A0 _05018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold571 top.CPU.registers.data\[584\] vssd1 vssd1 vccd1 vccd1 net3128 sky130_fd_sc_hd__dlygate4sd3_1
X_11020_ net1406 _03170_ net148 vssd1 vssd1 vccd1 vccd1 _06567_ sky130_fd_sc_hd__or3b_1
Xhold582 top.CPU.registers.data\[496\] vssd1 vssd1 vccd1 vccd1 net3139 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_173_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold593 top.CPU.registers.data\[139\] vssd1 vssd1 vccd1 vccd1 net3150 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10551__B _06173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout865_X net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07934__A1 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11730__A2 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_902 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12971_ net1411 _07406_ vssd1 vssd1 vccd1 vccd1 _07407_ sky130_fd_sc_hd__and2b_1
XANTENNA__13483__A2 net1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14188__358 clknet_leaf_194_clk vssd1 vssd1 vccd1 vccd1 net1827 sky130_fd_sc_hd__inv_2
XANTENNA__13354__S net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1260 top.CPU.registers.data\[414\] vssd1 vssd1 vccd1 vccd1 net3817 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1271 top.CPU.registers.data\[49\] vssd1 vssd1 vccd1 vccd1 net3828 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1282 _00026_ vssd1 vssd1 vccd1 vccd1 net3839 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12691__A0 top.CPU.alu.program_counter\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11922_ net3782 net184 net342 _06272_ vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__a22o_1
Xhold1293 top.mmio.mem_data_i\[13\] vssd1 vssd1 vccd1 vccd1 net3850 sky130_fd_sc_hd__dlygate4sd3_1
X_15690_ net2024 _01900_ net1087 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[490\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11853_ net457 _06687_ net233 net152 net2661 vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__a32o_1
X_14229__399 clknet_leaf_173_clk vssd1 vssd1 vccd1 vccd1 net1868 sky130_fd_sc_hd__inv_2
XFILLER_72_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10804_ _05700_ _05709_ vssd1 vssd1 vccd1 vccd1 _06414_ sky130_fd_sc_hd__nor2_1
X_11784_ _06629_ net197 net160 net3610 vssd1 vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__a22o_1
XFILLER_14_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08647__C1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16311_ clknet_leaf_96_clk _02520_ net1247 vssd1 vssd1 vccd1 vccd1 top.CPU.data_out\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13523_ _03716_ net584 vssd1 vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__and2_1
X_10735_ net548 _04862_ _06347_ _06348_ vssd1 vssd1 vccd1 vccd1 _06349_ sky130_fd_sc_hd__o211a_1
XANTENNA__07870__A0 _03508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16242_ clknet_leaf_44_clk _02452_ net1124 vssd1 vssd1 vccd1 vccd1 top.CPU.control_unit.instruction\[18\]
+ sky130_fd_sc_hd__dfrtp_4
X_10666_ _05671_ _05914_ _05923_ _06203_ vssd1 vssd1 vccd1 vccd1 _06283_ sky130_fd_sc_hd__o211ai_2
X_13454_ top.CPU.handler.toreg\[16\] _02948_ net123 vssd1 vssd1 vccd1 vccd1 _02482_
+ sky130_fd_sc_hd__mux2_1
XFILLER_173_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10726__B _06139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_201_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11549__A2 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12405_ _03120_ top.I2C.I2C_state\[9\] net2615 vssd1 vssd1 vccd1 vccd1 _00039_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_97_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13385_ top.I2C.data_out\[21\] net556 _02906_ vssd1 vssd1 vccd1 vccd1 _02907_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09072__C1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16173_ net2507 _02383_ net1069 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[973\]
+ sky130_fd_sc_hd__dfrtp_1
X_10597_ _04363_ _04430_ net373 vssd1 vssd1 vccd1 vccd1 _06217_ sky130_fd_sc_hd__mux2_1
XFILLER_12_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10757__B1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12210__A3 _06796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15124_ clknet_leaf_47_clk _01336_ net1131 vssd1 vssd1 vccd1 vccd1 top.I2C.within_byte_counter_reading\[2\]
+ sky130_fd_sc_hd__dfrtp_2
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__buf_2
XFILLER_127_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12336_ net2618 _04951_ net1219 vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15217__RESET_B net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15055_ clknet_leaf_50_clk _00052_ net1129 vssd1 vssd1 vccd1 vccd1 top.I2C.output_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12267_ net2807 _06391_ net433 vssd1 vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__mux2_1
XANTENNA__10742__A net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11218_ net532 net442 _05771_ net545 vssd1 vssd1 vccd1 vccd1 _06664_ sky130_fd_sc_hd__and4_1
X_14132__302 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 net1771 sky130_fd_sc_hd__inv_2
X_12198_ top.CPU.registers.data\[52\] net649 vssd1 vssd1 vccd1 vccd1 _06866_ sky130_fd_sc_hd__or2_1
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 DAT_O[20] sky130_fd_sc_hd__buf_2
XANTENNA__12005__Y _06780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput91 net91 vssd1 vssd1 vccd1 vccd1 DAT_O[30] sky130_fd_sc_hd__buf_2
XFILLER_150_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07925__A1 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11721__A2 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11149_ net572 net524 _06374_ vssd1 vssd1 vccd1 vccd1 _06634_ sky130_fd_sc_hd__and3_1
XANTENNA__09127__B1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15957_ net2291 _02167_ net1215 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[757\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11485__A1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08886__C1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15888_ net2222 _02098_ net1154 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[688\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_52_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09978__A net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08360_ _03997_ _03998_ net704 vssd1 vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__a21o_1
XANTENNA__11237__B2 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08638__C1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16509_ clknet_leaf_59_clk _02671_ net1137 vssd1 vssd1 vccd1 vccd1 top.mmio.mem_data_i\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11788__A2 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08291_ top.CPU.registers.data\[179\] top.CPU.registers.data\[147\] net825 vssd1
+ vssd1 vccd1 vccd1 _03930_ sky130_fd_sc_hd__mux2_1
XANTENNA__10917__A net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10460__A2 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14897__1067 clknet_leaf_188_clk vssd1 vssd1 vccd1 vccd1 net2536 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_115_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09063__C1 net1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08405__A2 net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08821__S net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11960__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09366__B1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout303 _06604_ vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__clkbuf_8
Xfanout314 net315 vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__buf_4
Xfanout325 _03190_ vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__buf_8
Xfanout336 net338 vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11712__A2 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10802__D net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout347 net349 vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__clkbuf_4
X_09814_ top.CPU.registers.data\[858\] net1335 net867 top.CPU.registers.data\[890\]
+ net758 vssd1 vssd1 vccd1 vccd1 _05453_ sky130_fd_sc_hd__a221o_1
XANTENNA__11186__C net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout358 net359 vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__buf_2
Xfanout369 _06576_ vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1100_A net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10920__B1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09745_ top.CPU.registers.data\[347\] net1331 net862 top.CPU.registers.data\[379\]
+ net775 vssd1 vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__a221o_1
XFILLER_28_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout560_A net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout181_X net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09669__A1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13465__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout279_X net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09676_ net710 _05314_ net638 vssd1 vssd1 vccd1 vccd1 _05315_ sky130_fd_sc_hd__a21o_1
XANTENNA__08877__C1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08627_ top.CPU.registers.data\[846\] net1320 net851 top.CPU.registers.data\[878\]
+ net769 vssd1 vssd1 vccd1 vccd1 _04266_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout446_X net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08892__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout825_A net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1188_X net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08558_ top.CPU.registers.data\[175\] net1387 vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__and2_1
XANTENNA__08629__C1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07509_ _03105_ net1279 vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__nand2_2
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout613_X net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08489_ top.CPU.registers.data\[48\] top.CPU.registers.data\[16\] net821 vssd1 vssd1
+ vccd1 vccd1 _04128_ sky130_fd_sc_hd__mux2_1
XFILLER_168_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09841__A1 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1355_X net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10520_ _03315_ _04193_ net506 _04189_ _06143_ vssd1 vssd1 vccd1 vccd1 _06144_ sky130_fd_sc_hd__a221o_1
XFILLER_52_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09099__S net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14573__743 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 net2212 sky130_fd_sc_hd__inv_2
XFILLER_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10451_ _06075_ _06077_ vssd1 vssd1 vccd1 vccd1 _06078_ sky130_fd_sc_hd__nor2_1
XANTENNA__09054__C1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10739__B1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13170_ top.I2C.within_byte_counter_reading\[2\] _06947_ vssd1 vssd1 vccd1 vccd1
+ _02755_ sky130_fd_sc_hd__nor2_2
X_10382_ net3642 net227 net318 _06011_ vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout982_X net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14614__784 clknet_leaf_175_clk vssd1 vssd1 vccd1 vccd1 net2253 sky130_fd_sc_hd__inv_2
X_12121_ net3945 net175 _06828_ _06647_ vssd1 vssd1 vccd1 vccd1 _01502_ sky130_fd_sc_hd__a22o_1
XANTENNA__11951__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12253__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09357__B1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12052_ net551 _03181_ net457 _06751_ vssd1 vssd1 vccd1 vccd1 _06795_ sky130_fd_sc_hd__or4_4
Xhold390 top.CPU.registers.data\[613\] vssd1 vssd1 vccd1 vccd1 net2947 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11003_ net3148 net216 _06556_ net312 vssd1 vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__a22o_1
XANTENNA__11703__A2 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11096__C net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08580__A1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09109__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout870 _03203_ vssd1 vssd1 vccd1 vccd1 net870 sky130_fd_sc_hd__buf_4
X_15811_ net2145 _02021_ net1212 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[611\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09415__X _05054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout881 net883 vssd1 vssd1 vccd1 vccd1 net881 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout892 net893 vssd1 vssd1 vccd1 vccd1 net892 sky130_fd_sc_hd__clkbuf_2
XFILLER_18_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15742_ net2076 _01952_ net1237 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[542\]
+ sky130_fd_sc_hd__dfrtp_1
X_12954_ top.CPU.alu.program_counter\[30\] _03409_ _07386_ vssd1 vssd1 vccd1 vccd1
+ _07393_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08868__C1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1090 top.CPU.registers.data\[609\] vssd1 vssd1 vccd1 vccd1 net3647 sky130_fd_sc_hd__dlygate4sd3_1
X_11905_ net3401 net185 net348 _05880_ vssd1 vssd1 vccd1 vccd1 _01661_ sky130_fd_sc_hd__a22o_1
X_15673_ net2007 _01883_ net1245 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[473\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_93_86 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12885_ _07310_ _07329_ _07328_ _07317_ vssd1 vssd1 vccd1 vccd1 _07331_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_193_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_193_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11219__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11836_ net466 _06667_ net243 net154 net2654 vssd1 vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__a32o_1
XANTENNA_clkbuf_leaf_97_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11767_ net470 _06610_ net241 net163 net3367 vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__a32o_1
XFILLER_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13506_ _04459_ _02966_ vssd1 vssd1 vccd1 vccd1 _02973_ sky130_fd_sc_hd__nor2_2
XANTENNA_clkbuf_leaf_140_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10718_ net601 _06331_ _06332_ vssd1 vssd1 vccd1 vccd1 _06333_ sky130_fd_sc_hd__a21oi_4
X_11698_ _06529_ net201 net421 net2986 vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__a22o_1
XFILLER_9_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16225_ clknet_leaf_33_clk _02435_ net1125 vssd1 vssd1 vccd1 vccd1 top.CPU.control_unit.instruction\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_13437_ net888 _02871_ _02937_ _02939_ vssd1 vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__a31o_1
XFILLER_42_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_20_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10649_ _06234_ _06256_ _06260_ _06266_ vssd1 vssd1 vccd1 vccd1 _06267_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_77_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16156_ net2490 _02366_ net1234 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[956\]
+ sky130_fd_sc_hd__dfrtp_1
X_13368_ net889 _02894_ vssd1 vssd1 vccd1 vccd1 _02895_ sky130_fd_sc_hd__and2_1
XANTENNA__09964__C _05367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12671__B _04955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_155_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14940__Q top.CPU.alu.program_counter\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15107_ net1489 _01320_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r2_prev\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11568__A net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11942__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12319_ net2571 _03783_ net1215 vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_110_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16087_ net2421 _02297_ net1182 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[887\]
+ sky130_fd_sc_hd__dfrtp_1
X_13299_ _02838_ _02839_ _02840_ _02841_ vssd1 vssd1 vccd1 vccd1 _02842_ sky130_fd_sc_hd__or4b_1
XANTENNA__09348__A0 top.CPU.alu.program_counter\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13144__A1 top.CPU.data_out\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_35_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15038_ clknet_leaf_91_clk _01283_ net1269 vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11287__B _06471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07860_ top.CPU.registers.data\[445\] net1009 net905 vssd1 vssd1 vccd1 vccd1 _03499_
+ sky130_fd_sc_hd__a21o_1
XFILLER_96_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10902__B1 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07791_ top.CPU.registers.data\[766\] net1384 net996 top.CPU.registers.data\[734\]
+ net920 vssd1 vssd1 vccd1 vccd1 _03430_ sky130_fd_sc_hd__a221o_1
XFILLER_49_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09530_ _05167_ _05168_ net780 vssd1 vssd1 vccd1 vccd1 _05169_ sky130_fd_sc_hd__mux2_1
XANTENNA__11458__B2 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09461_ net795 _05095_ _05096_ net748 vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__o211a_1
XFILLER_64_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_125_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_184_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_184_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11590__X _06749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08412_ _04048_ _04050_ net453 vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__mux2_1
X_09392_ top.CPU.registers.data\[419\] top.CPU.registers.data\[387\] net828 vssd1
+ vssd1 vccd1 vccd1 _05031_ sky130_fd_sc_hd__mux2_1
XANTENNA__12958__A1 top.CPU.alu.program_counter\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14260__430 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 net1899 sky130_fd_sc_hd__inv_2
XFILLER_149_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08343_ net955 _03960_ _03981_ net612 vssd1 vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__a211o_1
XANTENNA__08087__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14557__727 clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 net2196 sky130_fd_sc_hd__inv_2
XANTENNA__08626__A2 net1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout141_A _06105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09823__A1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_108_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout239_A net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08274_ net681 _03897_ _03898_ net923 vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__o211a_1
XANTENNA__07834__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14301__471 clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 net1940 sky130_fd_sc_hd__inv_2
XANTENNA__09036__C1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1050_A _03093_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_840 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout406_A net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12186__A2 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09587__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08551__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11394__B1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07598__C1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1315_A net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11197__B net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11146__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout775_A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1109 net1110 vssd1 vssd1 vccd1 vccd1 net1109 sky130_fd_sc_hd__buf_2
XFILLER_102_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout122 net124 vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__clkbuf_2
Xfanout133 _05990_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__buf_2
XANTENNA__09890__B _03613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout144 _06290_ vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__buf_2
Xfanout155 _06766_ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__buf_4
Xfanout166 _06757_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__buf_6
XANTENNA__08562__A1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout177 _06795_ vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__buf_2
Xfanout188 net191 vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__clkbuf_8
XFILLER_86_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout199 net202 vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout942_A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout563_X net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07989_ net676 _03622_ _03623_ _03627_ vssd1 vssd1 vccd1 vccd1 _03628_ sky130_fd_sc_hd__a31o_1
X_09728_ _05365_ _05366_ vssd1 vssd1 vccd1 vccd1 _05367_ sky130_fd_sc_hd__nand2b_4
XFILLER_47_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12110__A2 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09511__B1 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09659_ _03925_ _04052_ _05296_ _05295_ vssd1 vssd1 vccd1 vccd1 _05298_ sky130_fd_sc_hd__or4b_1
Xclkbuf_leaf_175_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_175_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout730_X net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13632__S net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout828_X net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12670_ top.CPU.alu.program_counter\[3\] _07136_ net1360 vssd1 vssd1 vccd1 vccd1
+ _01166_ sky130_fd_sc_hd__mux2_1
XFILLER_42_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13071__A0 top.CPU.data_out\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11621_ _06354_ net3346 net213 vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__mux2_1
XFILLER_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09275__C1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07825__B1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11552_ net3227 net247 _06740_ net485 vssd1 vssd1 vccd1 vccd1 _01983_ sky130_fd_sc_hd__a22o_1
XANTENNA__09290__A2 net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10503_ net3813 net226 net316 _06127_ vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__a22o_1
X_11483_ _06613_ net260 net256 net3233 vssd1 vssd1 vccd1 vccd1 _02041_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_94_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12177__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16010_ net2344 _02220_ net1084 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[810\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_155_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13222_ _02776_ net3686 _02794_ vssd1 vssd1 vccd1 vccd1 _01348_ sky130_fd_sc_hd__mux2_1
X_10434_ _05583_ _06060_ _05293_ vssd1 vssd1 vccd1 vccd1 _06061_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12491__B _04792_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11385__B1 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07589__C1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11924__A2 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13153_ top.I2C.output_state\[2\] top.I2C.output_state\[13\] top.I2C.output_state\[15\]
+ top.I2C.output_state\[28\] vssd1 vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__or4_1
X_10365_ _03916_ net506 vssd1 vssd1 vccd1 vccd1 _05995_ sky130_fd_sc_hd__nand2_1
X_13925__95 clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 net1564 sky130_fd_sc_hd__inv_2
XFILLER_98_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12104_ net566 net363 _06635_ net178 top.CPU.registers.data\[100\] vssd1 vssd1 vccd1
+ vccd1 _06820_ sky130_fd_sc_hd__a32o_1
X_13084_ top.CPU.data_out\[19\] net2726 net558 vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__mux2_1
X_10296_ _05921_ _05927_ _05928_ vssd1 vssd1 vccd1 vccd1 _05929_ sky130_fd_sc_hd__and3_1
XFILLER_3_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11137__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12035_ net3702 _06780_ _06792_ vssd1 vssd1 vccd1 vccd1 _01552_ sky130_fd_sc_hd__a21o_1
XANTENNA__11688__A1 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08002__B1 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07761__C1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14896__1066 clknet_leaf_199_clk vssd1 vssd1 vccd1 vccd1 net2535 sky130_fd_sc_hd__inv_2
XFILLER_81_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12101__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15725_ net2059 _01935_ net1077 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[525\]
+ sky130_fd_sc_hd__dfrtp_1
X_12937_ _07366_ _07371_ vssd1 vssd1 vccd1 vccd1 _07378_ sky130_fd_sc_hd__nor2_1
XANTENNA__10112__A1 _05399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_166_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_166_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_80_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14244__414 clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 net1883 sky130_fd_sc_hd__inv_2
XFILLER_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15656_ net1990 _01866_ net1098 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[456\]
+ sky130_fd_sc_hd__dfrtp_1
X_12868_ _07315_ _07312_ net126 vssd1 vssd1 vccd1 vccd1 _07316_ sky130_fd_sc_hd__mux2_1
XANTENNA__10738__Y _06352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09321__A net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08069__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11819_ net3379 net142 _06762_ vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__mux2_1
XANTENNA__09266__C1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15587_ net1921 _01797_ net1208 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[387\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08608__A2 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12799_ _07251_ _07252_ vssd1 vssd1 vccd1 vccd1 _07253_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10754__X _06367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12682__A top.CPU.alu.program_counter\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12168__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16208_ net2542 _02418_ net1154 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[1008\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13497__B _02966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08371__S net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09033__A2 net1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11376__B1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11915__A2 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11298__A net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16139_ net2473 _02349_ net1064 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[939\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08241__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16438__RESET_B net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_149_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08792__A1 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07595__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08961_ _04567_ _04599_ vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__and2_1
XFILLER_142_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07912_ net683 _03549_ _03550_ net608 vssd1 vssd1 vccd1 vccd1 _03551_ sky130_fd_sc_hd__a31o_1
XFILLER_68_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08892_ top.CPU.registers.data_out_r1_prev\[11\] net871 net640 _04527_ _04530_ vssd1
+ vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__o221a_4
XANTENNA__10930__A net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1036 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08544__A1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07843_ top.CPU.registers.data\[93\] net1288 net1007 top.CPU.registers.data\[125\]
+ net932 vssd1 vssd1 vccd1 vccd1 _03482_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_162_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_162_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout189_A net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07774_ top.CPU.registers.data\[190\] net1384 net997 top.CPU.registers.data\[158\]
+ vssd1 vssd1 vccd1 vccd1 _03413_ sky130_fd_sc_hd__a22o_1
XFILLER_17_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Left_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09513_ net622 _05147_ _05148_ _05151_ vssd1 vssd1 vccd1 vccd1 _05152_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_157_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_157_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11300__B1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13452__S net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11761__A net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09444_ net612 _05079_ _05082_ net627 vssd1 vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_140_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_166_Right_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09257__C1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09375_ net939 _04992_ _04993_ net956 vssd1 vssd1 vccd1 vccd1 _05014_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout144_X net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08326_ top.CPU.registers.data\[979\] net1295 net1017 top.CPU.registers.data\[1011\]
+ net911 vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__a221o_1
XANTENNA__07807__B1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14028__198 clknet_leaf_195_clk vssd1 vssd1 vccd1 vccd1 net1667 sky130_fd_sc_hd__inv_2
XANTENNA__10096__B net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08257_ top.CPU.registers.data\[470\] net1300 net1021 top.CPU.registers.data\[502\]
+ net917 vssd1 vssd1 vccd1 vccd1 _03896_ sky130_fd_sc_hd__a221o_1
XANTENNA__09009__C1 net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout311_X net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1053_X net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout409_X net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12159__A2 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08188_ top.CPU.registers.data\[151\] net987 _03826_ vssd1 vssd1 vccd1 vccd1 _03827_
+ sky130_fd_sc_hd__a21o_1
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11367__B1 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11906__A2 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08232__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11001__A net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10150_ net390 _05786_ vssd1 vssd1 vccd1 vccd1 _05787_ sky130_fd_sc_hd__nand2_1
XFILLER_134_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11119__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout680_X net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14685__855 clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 net2324 sky130_fd_sc_hd__inv_2
XANTENNA_fanout778_X net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07991__C1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10081_ _04430_ _04532_ net378 vssd1 vssd1 vccd1 vccd1 _05719_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10840__A net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout945_X net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16300__Q top.CPU.data_out\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14726__896 clknet_leaf_125_clk vssd1 vssd1 vccd1 vccd1 net2365 sky130_fd_sc_hd__inv_2
XFILLER_75_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12095__A1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13771_ net30 net1049 net884 net3545 vssd1 vssd1 vccd1 vccd1 _02652_ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_148_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_148_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12767__A top.CPU.alu.program_counter\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10983_ net3751 net217 _06544_ net314 vssd1 vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__a22o_1
XFILLER_83_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15510_ net1844 _01720_ net1229 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[310\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12722_ top.CPU.alu.program_counter\[9\] _04660_ vssd1 vssd1 vccd1 vccd1 _07183_
+ sky130_fd_sc_hd__nand2_1
X_16490_ clknet_leaf_40_clk _02652_ net1115 vssd1 vssd1 vccd1 vccd1 top.mmio.mem_data_i\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08456__S net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_133_Right_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15441_ net1775 _01651_ net1191 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[241\]
+ sky130_fd_sc_hd__dfrtp_1
X_12653_ net1043 _07053_ vssd1 vssd1 vccd1 vccd1 _07121_ sky130_fd_sc_hd__or2_1
XFILLER_130_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11604_ net133 net3579 net214 vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__mux2_1
XFILLER_129_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15372_ net1706 _01582_ net1076 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[172\]
+ sky130_fd_sc_hd__dfrtp_1
X_12584_ _06925_ _07087_ vssd1 vssd1 vccd1 vccd1 _07088_ sky130_fd_sc_hd__nor2_2
XFILLER_12_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09263__A2 net1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11535_ _06657_ net259 net250 net3587 vssd1 vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__a22o_1
XANTENNA__11070__A2 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11610__S net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08044__X _03683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11466_ _06354_ net3646 net263 vssd1 vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__mux2_1
XFILLER_172_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11358__B1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13205_ net892 top.I2C.data_out\[19\] _02782_ vssd1 vssd1 vccd1 vccd1 _02783_ sky130_fd_sc_hd__mux2_1
X_10417_ net406 _06041_ _06043_ _05827_ vssd1 vssd1 vccd1 vccd1 _06045_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_124_331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09420__C1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11397_ net570 net540 _06603_ net1403 vssd1 vssd1 vccd1 vccd1 _06716_ sky130_fd_sc_hd__or4b_1
XFILLER_98_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13136_ top.SPI.command\[1\] _02732_ _02733_ top.SPI.counter\[2\] vssd1 vssd1 vccd1
+ vccd1 _02737_ sky130_fd_sc_hd__a22o_1
XANTENNA__12570__A2 _06081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_727 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10348_ net404 _05663_ _05978_ vssd1 vssd1 vccd1 vccd1 _05979_ sky130_fd_sc_hd__o21a_1
XFILLER_97_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10279_ _05858_ _05911_ net308 vssd1 vssd1 vccd1 vccd1 _05912_ sky130_fd_sc_hd__mux2_1
X_13067_ top.CPU.data_out\[2\] net2702 net559 vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__mux2_1
XFILLER_140_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09723__B1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12018_ net3211 _06781_ vssd1 vssd1 vccd1 vccd1 _06786_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_144_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11530__B1 _06734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10884__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09750__S net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_139_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_139_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_85_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10097__B1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13272__S _06948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15708_ net2042 _01918_ net1194 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[508\]
+ sky130_fd_sc_hd__dfrtp_1
X_07490_ net1346 vssd1 vssd1 vccd1 vccd1 _03130_ sky130_fd_sc_hd__inv_2
XFILLER_94_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11833__A1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08366__S net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15639_ net1973 _01849_ net1180 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[439\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09239__C1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09160_ top.CPU.registers.data\[166\] top.CPU.registers.data\[134\] net814 vssd1
+ vssd1 vccd1 vccd1 _04799_ sky130_fd_sc_hd__mux2_1
XFILLER_148_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09986__A _04765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08890__A net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11597__A0 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08111_ top.CPU.registers.data\[949\] top.CPU.registers.data\[917\] net830 vssd1
+ vssd1 vccd1 vccd1 _03750_ sky130_fd_sc_hd__mux2_1
X_09091_ _04698_ _04729_ vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__nand2_1
XANTENNA__11061__A2 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08462__B1 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10925__A _06333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09197__S net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08042_ top.CPU.registers.data_out_r1_prev\[20\] net873 vssd1 vssd1 vccd1 vccd1 _03681_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__11349__B1 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold901 top.CPU.registers.data\[843\] vssd1 vssd1 vccd1 vccd1 net3458 sky130_fd_sc_hd__dlygate4sd3_1
Xhold912 top.CPU.registers.data\[758\] vssd1 vssd1 vccd1 vccd1 net3469 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap631 _03303_ vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__buf_1
Xhold923 top.CPU.registers.data\[219\] vssd1 vssd1 vccd1 vccd1 net3480 sky130_fd_sc_hd__dlygate4sd3_1
X_14372__542 clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 net2011 sky130_fd_sc_hd__inv_2
Xhold934 top.CPU.registers.data\[958\] vssd1 vssd1 vccd1 vccd1 net3491 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09411__C1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold945 top.CPU.registers.data\[598\] vssd1 vssd1 vccd1 vccd1 net3502 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16612__A net1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14669__839 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 net2308 sky130_fd_sc_hd__inv_2
XFILLER_143_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08765__A1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold956 top.CPU.registers.data\[916\] vssd1 vssd1 vccd1 vccd1 net3513 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold967 top.CPU.registers.data\[743\] vssd1 vssd1 vccd1 vccd1 net3524 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold978 top.CPU.registers.data\[187\] vssd1 vssd1 vccd1 vccd1 net3535 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_164_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09993_ _05624_ _05631_ net386 vssd1 vssd1 vccd1 vccd1 _05632_ sky130_fd_sc_hd__mux2_1
Xhold989 top.CPU.registers.data\[260\] vssd1 vssd1 vccd1 vccd1 net3546 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_164_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08944_ top.CPU.registers.data\[586\] net1374 net971 top.CPU.registers.data\[618\]
+ net902 vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__o221a_1
X_14413__583 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 net2052 sky130_fd_sc_hd__inv_2
XFILLER_103_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1013_A net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10324__A1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08875_ top.CPU.registers.data\[427\] top.CPU.registers.data\[395\] net807 vssd1
+ vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout473_A _03193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07725__C1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09190__A1 _04828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07826_ top.CPU.registers.data\[445\] top.CPU.registers.data\[413\] net816 vssd1
+ vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__mux2_1
XANTENNA__10875__A2 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09478__C1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout261_X net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout640_A net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07757_ top.CPU.registers.data\[62\] top.CPU.registers.data\[30\] net834 vssd1 vssd1
+ vccd1 vccd1 _03396_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout738_A net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout359_X net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1382_A net1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07688_ _03249_ _03259_ _03261_ _03273_ vssd1 vssd1 vccd1 vccd1 _03327_ sky130_fd_sc_hd__a31o_1
XFILLER_25_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10819__B _06428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09427_ net677 _05064_ _05065_ net911 vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__o211a_1
XFILLER_13_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1170_X net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout526_X net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout905_A net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13577__A1 top.CPU.alu.program_counter\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09358_ top.CPU.registers.data\[963\] net1297 net1018 top.CPU.registers.data\[995\]
+ net915 vssd1 vssd1 vccd1 vccd1 _04997_ sky130_fd_sc_hd__a221o_1
XFILLER_100_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11588__B1 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13980__150 clknet_leaf_135_clk vssd1 vssd1 vccd1 vccd1 net1619 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_43_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08309_ top.CPU.registers.data\[659\] net1327 net858 top.CPU.registers.data\[691\]
+ net724 vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_23_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11052__A2 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09289_ top.CPU.registers.data\[324\] net1299 net1020 top.CPU.registers.data\[356\]
+ net940 vssd1 vssd1 vccd1 vccd1 _04928_ sky130_fd_sc_hd__a221o_1
X_11320_ net3444 net292 _06710_ net492 vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__a22o_1
XFILLER_138_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14895__1065 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 net2534 sky130_fd_sc_hd__inv_2
XFILLER_5_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11251_ net516 _06549_ vssd1 vssd1 vccd1 vccd1 _06681_ sky130_fd_sc_hd__nor2_1
XANTENNA__09402__C1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10012__A0 _03476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10202_ net383 _05723_ vssd1 vssd1 vccd1 vccd1 _05838_ sky130_fd_sc_hd__nand2_1
XFILLER_122_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11182_ net3643 net299 _06650_ net317 vssd1 vssd1 vccd1 vccd1 _02263_ sky130_fd_sc_hd__a22o_1
XFILLER_162_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10563__A1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11760__B1 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07964__C1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10133_ _05768_ _05769_ _05770_ net661 vssd1 vssd1 vccd1 vccd1 _05771_ sky130_fd_sc_hd__o31a_1
XFILLER_79_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12261__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15990_ net2324 _02200_ net1229 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[790\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10570__A net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13501__A1 top.CPU.data_out\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09705__B1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14941_ clknet_leaf_73_clk _01187_ net1158 vssd1 vssd1 vccd1 vccd1 top.CPU.alu.program_counter\[24\]
+ sky130_fd_sc_hd__dfrtp_4
X_10064_ net383 _05700_ _05701_ vssd1 vssd1 vccd1 vccd1 _05702_ sky130_fd_sc_hd__or3_1
XANTENNA_input34_A en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11512__B1 _06734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13823_ net3690 net336 net329 top.CPU.data_out\[25\] vssd1 vssd1 vccd1 vccd1 _02703_
+ sky130_fd_sc_hd__a22o_1
XFILLER_29_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13092__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16542_ clknet_leaf_86_clk net3111 net1266 vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__dfrtp_1
X_13754_ _02772_ _02791_ top.I2C.I2C_state\[16\] vssd1 vssd1 vccd1 vccd1 _03088_ sky130_fd_sc_hd__or3b_1
X_10966_ net3512 net219 _06534_ net319 vssd1 vssd1 vccd1 vccd1 _02363_ sky130_fd_sc_hd__a22o_1
XANTENNA__09484__A2 _05120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08141__C1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12705_ top.CPU.alu.program_counter\[7\] _04793_ vssd1 vssd1 vccd1 vccd1 _07168_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_100_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16473_ clknet_leaf_88_clk _02635_ net1273 vssd1 vssd1 vccd1 vccd1 top.SPI.timem\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13685_ net2699 net336 vssd1 vssd1 vccd1 vccd1 _02613_ sky130_fd_sc_hd__and2_1
X_10897_ net132 net437 vssd1 vssd1 vccd1 vccd1 _06492_ sky130_fd_sc_hd__and2_1
X_15424_ net1758 _01634_ net1092 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[224\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12636_ top.I2C.output_state\[14\] net3662 vssd1 vssd1 vccd1 vccd1 _00011_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_80_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11579__B1 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12944__B _03409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15355_ net1689 _01565_ net1213 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[155\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08444__B1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12240__A1 _05771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11043__A2 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12567_ _06268_ _06288_ _07071_ vssd1 vssd1 vccd1 vccd1 _07072_ sky130_fd_sc_hd__or3_1
XFILLER_156_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10251__A0 _05399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14356__526 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 net1995 sky130_fd_sc_hd__inv_2
XFILLER_144_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08995__A1 _04633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11518_ net3914 net253 _06734_ _06480_ vssd1 vssd1 vccd1 vccd1 _02012_ sky130_fd_sc_hd__a22o_1
XFILLER_156_275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15286_ net1620 _01496_ net1230 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[86\]
+ sky130_fd_sc_hd__dfrtp_1
X_12498_ _07005_ _07006_ _07004_ vssd1 vssd1 vccd1 vccd1 _07007_ sky130_fd_sc_hd__a21bo_1
XFILLER_8_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold208 top.SPI.paroutput\[23\] vssd1 vssd1 vccd1 vccd1 net2765 sky130_fd_sc_hd__dlygate4sd3_1
Xhold219 net119 vssd1 vssd1 vccd1 vccd1 net2776 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11449_ net565 net440 _06085_ net538 vssd1 vssd1 vccd1 vccd1 _06724_ sky130_fd_sc_hd__and4_1
XANTENNA__12960__A top.CPU.alu.program_counter\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11279__C net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14100__270 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 net1739 sky130_fd_sc_hd__inv_2
XANTENNA__08747__A1 net1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11751__B1 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13119_ net2686 _02724_ net897 vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__mux2_1
XFILLER_140_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_84_Left_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10480__A _03167_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10911__C _06500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07970__A2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1270 net1275 vssd1 vssd1 vccd1 vccd1 net1270 sky130_fd_sc_hd__clkbuf_4
XANTENNA__15665__RESET_B net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1281 net1282 vssd1 vssd1 vccd1 vccd1 net1281 sky130_fd_sc_hd__clkbuf_4
X_08660_ top.CPU.registers.data\[334\] net1375 net981 top.CPU.registers.data\[366\]
+ net1282 vssd1 vssd1 vccd1 vccd1 _04299_ sky130_fd_sc_hd__o221a_1
Xfanout1292 net1293 vssd1 vssd1 vccd1 vccd1 net1292 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08885__A net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07611_ net1400 _03249_ _03247_ _03246_ vssd1 vssd1 vccd1 vccd1 _03250_ sky130_fd_sc_hd__a211o_1
XANTENNA__10479__X _06105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08591_ top.CPU.registers.data\[335\] net1374 net974 top.CPU.registers.data\[367\]
+ net1281 vssd1 vssd1 vccd1 vccd1 _04230_ sky130_fd_sc_hd__o221a_1
XFILLER_54_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10609__A2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07542_ net1403 net660 vssd1 vssd1 vccd1 vccd1 _03181_ sky130_fd_sc_hd__and2_2
XANTENNA__09475__A2 net1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08132__C1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13008__B1 _07431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07473_ net1371 vssd1 vssd1 vccd1 vccd1 _03113_ sky130_fd_sc_hd__clkinv_4
XPHY_EDGE_ROW_93_Left_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11282__A2 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09880__C1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13964__134 clknet_leaf_191_clk vssd1 vssd1 vccd1 vccd1 net1603 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_157_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13559__A1 _03137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09212_ top.CPU.registers.data\[326\] net1287 net1006 top.CPU.registers.data\[358\]
+ net930 vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_157_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_174_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11034__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09143_ top.CPU.registers.data\[327\] net1302 net1024 top.CPU.registers.data\[359\]
+ net943 vssd1 vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__a221o_1
XANTENNA__12231__A1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16453__RESET_B net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout221_A _06469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10242__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07789__A2 net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout319_A net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09074_ top.CPU.registers.data\[968\] net1376 net975 top.CPU.registers.data\[1000\]
+ net1364 vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__o221a_1
X_14099__269 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 net1738 sky130_fd_sc_hd__inv_2
XFILLER_148_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11990__B1 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08025_ net791 _03658_ _03659_ net743 vssd1 vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout1130_A net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12870__A top.CPU.alu.program_counter\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold720 top.CPU.registers.data\[725\] vssd1 vssd1 vccd1 vccd1 net3277 sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 top.CPU.registers.data\[580\] vssd1 vssd1 vccd1 vccd1 net3288 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08738__A1 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold742 top.CPU.registers.data\[871\] vssd1 vssd1 vccd1 vccd1 net3299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold753 top.CPU.registers.data\[133\] vssd1 vssd1 vccd1 vccd1 net3310 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold764 top.CPU.registers.data\[427\] vssd1 vssd1 vccd1 vccd1 net3321 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout590_A net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold775 top.CPU.registers.data\[158\] vssd1 vssd1 vccd1 vccd1 net3332 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_118_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold786 net71 vssd1 vssd1 vccd1 vccd1 net3343 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout688_A _03332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11742__B1 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07946__C1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold797 net73 vssd1 vssd1 vccd1 vccd1 net3354 sky130_fd_sc_hd__dlygate4sd3_1
X_09976_ _03375_ _05526_ _05614_ _05610_ net445 vssd1 vssd1 vccd1 vccd1 _05615_ sky130_fd_sc_hd__a311o_1
XFILLER_162_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1016_X net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12298__A1 _04566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08927_ _04551_ _04565_ vssd1 vssd1 vccd1 vccd1 _04566_ sky130_fd_sc_hd__nor2_4
XFILLER_76_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout855_A net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09699__C1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1420 top.CPU.addressnew\[14\] vssd1 vssd1 vccd1 vccd1 net3977 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout476_X net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1431 top.CPU.registers.data\[108\] vssd1 vssd1 vccd1 vccd1 net3988 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1442 top.CPU.addressnew\[10\] vssd1 vssd1 vccd1 vccd1 net3999 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08858_ _04483_ _04496_ vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__nor2_4
Xhold1453 top.mmio.mem_data_i\[30\] vssd1 vssd1 vccd1 vccd1 net4010 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09390__S net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1464 top.CPU.registers.data_out_r1_prev\[2\] vssd1 vssd1 vccd1 vccd1 net4021
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08910__A1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11933__B net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07809_ top.CPU.registers.data\[989\] net1318 net849 top.CPU.registers.data\[1021\]
+ net692 vssd1 vssd1 vccd1 vccd1 _03448_ sky130_fd_sc_hd__a221o_1
X_08789_ _04427_ vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout643_X net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1385_X net1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10820_ net574 net518 _06429_ vssd1 vssd1 vccd1 vccd1 _06430_ sky130_fd_sc_hd__and3_1
X_14797__967 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 net2436 sky130_fd_sc_hd__inv_2
XANTENNA__13798__B2 top.CPU.data_out\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10751_ net402 _06199_ vssd1 vssd1 vccd1 vccd1 _06364_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout810_X net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout908_X net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13640__S net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14043__213 clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 net1682 sky130_fd_sc_hd__inv_2
X_13470_ top.CPU.handler.toreg\[24\] _02956_ net123 vssd1 vssd1 vccd1 vccd1 _02490_
+ sky130_fd_sc_hd__mux2_1
X_10682_ net400 _06137_ net411 vssd1 vssd1 vccd1 vccd1 _06298_ sky130_fd_sc_hd__o21a_1
XANTENNA__08734__S net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12421_ net4025 _06941_ _06946_ vssd1 vssd1 vccd1 vccd1 _00069_ sky130_fd_sc_hd__a21bo_1
XANTENNA__09623__C1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12256__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15140_ clknet_leaf_59_clk _01350_ net1140 vssd1 vssd1 vccd1 vccd1 top.I2C.data_out\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_138_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12352_ net1339 top.I2C.output_state\[23\] net2791 vssd1 vssd1 vccd1 vccd1 _06898_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_126_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16123__RESET_B net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11981__B1 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11303_ net3228 net292 _06708_ net496 vssd1 vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__a22o_1
X_15071_ clknet_leaf_50_clk _00049_ net1129 vssd1 vssd1 vccd1 vccd1 top.I2C.output_state\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_126_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12283_ net3808 _03820_ net1184 vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__mux2_1
XFILLER_4_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09077__S1 net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09565__S net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11234_ net530 _06010_ _06523_ vssd1 vssd1 vccd1 vccd1 _06672_ sky130_fd_sc_hd__and3_1
XANTENNA__10536__B2 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11733__B1 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11165_ net458 net429 vssd1 vssd1 vccd1 vccd1 _06644_ sky130_fd_sc_hd__nand2_1
X_10116_ net402 _05642_ vssd1 vssd1 vccd1 vccd1 _05754_ sky130_fd_sc_hd__nand2_4
XFILLER_110_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13486__A0 top.CPU.data_out\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15973_ net2307 _02183_ net1062 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[773\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12289__A1 _04019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11096_ net1407 net577 net532 net137 vssd1 vssd1 vccd1 vccd1 _06606_ sky130_fd_sc_hd__and4_1
XFILLER_110_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09154__A1 top.CPU.control_unit.instruction\[27\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14741__911 clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 net2380 sky130_fd_sc_hd__inv_2
X_10047_ _03286_ _03297_ _03304_ _03310_ vssd1 vssd1 vccd1 vccd1 _05686_ sky130_fd_sc_hd__or4b_1
X_14924_ clknet_leaf_32_clk _01170_ net1125 vssd1 vssd1 vccd1 vccd1 top.CPU.alu.program_counter\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_49_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold80 top.CPU.addressnew\[26\] vssd1 vssd1 vccd1 vccd1 net2637 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09153__X _04792_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08362__C1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold91 top.CPU.registers.data\[545\] vssd1 vssd1 vccd1 vccd1 net2648 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_63_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13806_ net3484 net333 net326 top.CPU.data_out\[8\] vssd1 vssd1 vccd1 vccd1 _02686_
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13948__118 clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 net1587 sky130_fd_sc_hd__inv_2
XANTENNA__09457__A2 net1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11998_ _06566_ net348 net182 net3037 vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__a22o_1
XANTENNA__10459__B net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16525_ clknet_leaf_100_clk _02687_ net1255 vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__dfrtp_1
X_13737_ top.SPI.timem\[17\] _03077_ _07113_ vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_27_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10949_ net1406 _03170_ vssd1 vssd1 vccd1 vccd1 _06524_ sky130_fd_sc_hd__or2_1
XFILLER_31_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_70_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_clk sky130_fd_sc_hd__clkbuf_8
X_16456_ clknet_leaf_58_clk net1346 net1144 vssd1 vssd1 vccd1 vccd1 top.wm.prev_BUSY_O
+ sky130_fd_sc_hd__dfrtp_1
X_13668_ net2859 net331 net330 top.CPU.addressnew\[1\] vssd1 vssd1 vccd1 vccd1 _02596_
+ sky130_fd_sc_hd__a22o_1
XFILLER_31_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14943__Q top.CPU.alu.program_counter\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15407_ net1741 _01617_ net1109 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[207\]
+ sky130_fd_sc_hd__dfrtp_1
X_12619_ _07101_ top.SPI.nextwrx vssd1 vssd1 vccd1 vccd1 _07117_ sky130_fd_sc_hd__nand2_1
XANTENNA__11016__A2 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16387_ clknet_leaf_89_clk _00072_ net1273 vssd1 vssd1 vccd1 vccd1 top.SPI.state\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__13410__B1 net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13599_ net578 _03026_ _03024_ vssd1 vssd1 vccd1 vccd1 _02549_ sky130_fd_sc_hd__o21ai_1
XFILLER_157_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09614__C1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15338_ net1672 _01548_ net1091 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[138\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_117_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11972__B1 net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15269_ net1603 _01479_ net1087 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[69\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_113_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11724__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08196__A2 net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout507 _05676_ vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_130_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09830_ top.CPU.registers.data\[26\] net1000 _05468_ vssd1 vssd1 vccd1 vccd1 _05469_
+ sky130_fd_sc_hd__a21o_1
Xfanout518 net522 vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__buf_4
Xfanout529 net533 vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__clkbuf_2
XFILLER_112_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09761_ top.CPU.registers.data\[827\] top.CPU.registers.data\[795\] net990 vssd1
+ vssd1 vccd1 vccd1 _05400_ sky130_fd_sc_hd__mux2_1
XANTENNA__13477__B1 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13886__56 clknet_leaf_150_clk vssd1 vssd1 vccd1 vccd1 net1525 sky130_fd_sc_hd__inv_2
XFILLER_112_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11593__X _06752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08712_ top.CPU.registers.data\[461\] net1311 net842 top.CPU.registers.data\[493\]
+ net762 vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__a221o_1
XFILLER_39_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14484__654 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 net2123 sky130_fd_sc_hd__inv_2
X_09692_ _05330_ vssd1 vssd1 vccd1 vccd1 _05331_ sky130_fd_sc_hd__inv_2
XFILLER_94_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08643_ net706 _04278_ _04281_ vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__or3_1
X_14894__1064 clknet_leaf_122_clk vssd1 vssd1 vccd1 vccd1 net2533 sky130_fd_sc_hd__inv_2
XFILLER_148_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12568__C _06251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout269_A net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08574_ net740 _04211_ _04212_ net766 vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__o211a_1
XFILLER_25_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14525__695 clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 net2164 sky130_fd_sc_hd__inv_2
XANTENNA__08105__C1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07525_ net1279 _03153_ _03157_ _03144_ vssd1 vssd1 vccd1 vccd1 _03164_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_25_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12865__A top.CPU.alu.program_counter\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_61_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout436_A _06467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1178_A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13401__A0 top.CPU.control_unit.instruction\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07678__B net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout224_X net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09605__C1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1345_A net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09126_ net1034 _04763_ _04733_ vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__a21oi_2
XANTENNA__11963__B1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09057_ top.CPU.registers.data_out_r1_prev\[8\] net871 net635 _04695_ _04681_ vssd1
+ vssd1 vccd1 vccd1 _04696_ sky130_fd_sc_hd__o221ai_2
XANTENNA__09385__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08008_ _03645_ _03646_ net453 vssd1 vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__mux2_1
Xhold550 top.CPU.registers.data\[615\] vssd1 vssd1 vccd1 vccd1 net3107 sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 top.CPU.fetch.current_ra\[0\] vssd1 vssd1 vccd1 vccd1 net3118 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout972_A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold572 top.CPU.fetch.current_ra\[28\] vssd1 vssd1 vccd1 vccd1 net3129 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11715__B1 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07919__C1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09384__A1 _05021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08187__A2 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold583 top.CPU.registers.data\[14\] vssd1 vssd1 vccd1 vccd1 net3140 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold594 top.CPU.registers.data\[630\] vssd1 vssd1 vccd1 vccd1 net3151 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_173_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11191__B2 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08592__C1 net1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13468__A0 top.CPU.handler.toreg\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09959_ _03650_ _05367_ _05594_ _05597_ vssd1 vssd1 vccd1 vccd1 _05598_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout760_X net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout858_X net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13635__S net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12970_ top.I2C.bit_timer_counter\[1\] top.I2C.bit_timer_counter\[0\] top.I2C.bit_timer_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _07406_ sky130_fd_sc_hd__and3_1
XFILLER_46_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08344__C1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1250 top.CPU.registers.data\[654\] vssd1 vssd1 vccd1 vccd1 net3807 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09687__A2 net1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13483__A3 _03200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1261 top.CPU.registers.data\[491\] vssd1 vssd1 vccd1 vccd1 net3818 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11921_ net3780 net184 net343 _06255_ vssd1 vssd1 vccd1 vccd1 _01645_ sky130_fd_sc_hd__a22o_1
Xhold1272 top.CPU.registers.data\[129\] vssd1 vssd1 vccd1 vccd1 net3829 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11494__A2 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1283 top.CPU.registers.data\[858\] vssd1 vssd1 vccd1 vccd1 net3840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1294 top.CPU.registers.data\[131\] vssd1 vssd1 vccd1 vccd1 net3851 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11852_ _06686_ net234 net152 net2858 vssd1 vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__a22o_1
XANTENNA__09439__A2 net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10803_ net3618 net226 net317 _06413_ vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__a22o_1
XFILLER_32_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08647__B1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11783_ _06628_ net199 net160 net3192 vssd1 vssd1 vccd1 vccd1 _01772_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_52_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09844__C1 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16310_ clknet_leaf_96_clk _02519_ net1249 vssd1 vssd1 vccd1 vccd1 top.CPU.data_out\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13522_ top.CPU.data_out\[19\] net591 net339 _02981_ vssd1 vssd1 vccd1 vccd1 _02517_
+ sky130_fd_sc_hd__o22a_1
XFILLER_14_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10734_ _04861_ net508 net503 _04859_ net443 vssd1 vssd1 vccd1 vccd1 _06348_ sky130_fd_sc_hd__o221a_1
XANTENNA__11797__A3 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16241_ clknet_leaf_45_clk _02451_ net1138 vssd1 vssd1 vccd1 vccd1 top.CPU.control_unit.instruction\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07870__A1 _03477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13453_ net1396 net872 _02895_ net419 vssd1 vssd1 vccd1 vccd1 _02948_ sky130_fd_sc_hd__a31o_1
XFILLER_51_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10665_ net408 _06113_ _06281_ net414 vssd1 vssd1 vccd1 vccd1 _06282_ sky130_fd_sc_hd__a211o_1
XFILLER_139_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_149_Left_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12404_ _03125_ top.I2C.I2C_state\[4\] net2620 vssd1 vssd1 vccd1 vccd1 _00034_ sky130_fd_sc_hd__a21o_1
XFILLER_173_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16172_ net2506 _02382_ net1070 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[972\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13384_ net1345 top.mmio.mem_data_i\[21\] net597 vssd1 vssd1 vccd1 vccd1 _02906_
+ sky130_fd_sc_hd__o21a_1
XFILLER_12_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_97_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10596_ _04469_ _05284_ _06215_ vssd1 vssd1 vccd1 vccd1 _06216_ sky130_fd_sc_hd__a21o_1
XFILLER_12_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15123_ clknet_leaf_50_clk _01335_ net1131 vssd1 vssd1 vccd1 vccd1 top.I2C.within_byte_counter_reading\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_127_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12335_ net2588 _04918_ net1083 vssd1 vssd1 vccd1 vccd1 _01306_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15054_ clknet_leaf_55_clk _00042_ net1135 vssd1 vssd1 vccd1 vccd1 top.I2C.output_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_12266_ net2937 _06373_ net431 vssd1 vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__mux2_1
XANTENNA__11706__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10742__B net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09375__A1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11217_ net496 net469 _06663_ net295 net2642 vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__a32o_1
X_12197_ net3764 net654 _06865_ vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__o21a_1
X_14171__341 clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 net1810 sky130_fd_sc_hd__inv_2
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 DAT_O[11] sky130_fd_sc_hd__buf_2
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 DAT_O[21] sky130_fd_sc_hd__buf_2
XANTENNA__11182__B2 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput92 net92 vssd1 vssd1 vccd1 vccd1 DAT_O[31] sky130_fd_sc_hd__buf_2
X_14468__638 clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 net2107 sky130_fd_sc_hd__inv_2
XFILLER_150_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11148_ net483 net459 _06633_ net302 net3314 vssd1 vssd1 vccd1 vccd1 _02280_ sky130_fd_sc_hd__a32o_1
XANTENNA__13459__B1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_158_Left_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11079_ _03190_ net147 net538 net368 net2753 vssd1 vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__a32o_1
X_15956_ net2290 _02166_ net1072 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[756\]
+ sky130_fd_sc_hd__dfrtp_1
X_14212__382 clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 net1851 sky130_fd_sc_hd__inv_2
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09678__A2 net1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08886__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15887_ net2221 _02097_ net1095 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[687\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11485__A2 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14509__679 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 net2148 sky130_fd_sc_hd__inv_2
XANTENNA__11237__A2 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09978__B _05616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08638__B1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_43_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08102__A2 net1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16508_ clknet_leaf_57_clk _02670_ net1144 vssd1 vssd1 vccd1 vccd1 top.mmio.mem_data_i\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_08290_ top.CPU.registers.data\[83\] net1326 net857 top.CPU.registers.data\[115\]
+ net773 vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_154_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10917__B net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_9_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_167_Left_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_171_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16439_ clknet_leaf_80_clk net3607 net1242 vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__dfrtp_1
XFILLER_164_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09063__B1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09602__A2 net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_132_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08169__A2 net1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout304 _06604_ vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16620__A net1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout315 _03195_ vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__buf_4
XFILLER_115_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout326 net327 vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__buf_2
XANTENNA__08574__C1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout337 net338 vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__clkbuf_2
XFILLER_143_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09813_ top.CPU.registers.data\[986\] net1335 net867 top.CPU.registers.data\[1018\]
+ net732 vssd1 vssd1 vccd1 vccd1 _05452_ sky130_fd_sc_hd__a221o_1
XFILLER_86_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout348 net349 vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__clkbuf_4
XFILLER_98_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10920__A1 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout359 _06704_ vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__buf_8
XANTENNA_fanout386_A net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09118__A1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09744_ top.CPU.registers.data\[315\] top.CPU.registers.data\[283\] net827 vssd1
+ vssd1 vccd1 vccd1 _05383_ sky130_fd_sc_hd__mux2_1
XFILLER_55_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08326__C1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12122__B1 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09675_ _05312_ _05313_ net757 vssd1 vssd1 vccd1 vccd1 _05314_ sky130_fd_sc_hd__mux2_1
XFILLER_36_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout174_X net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1295_A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08626_ top.CPU.registers.data\[590\] net1320 net851 top.CPU.registers.data\[622\]
+ net744 vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__a221o_1
XFILLER_55_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08557_ top.CPU.registers.data\[79\] net1314 net845 top.CPU.registers.data\[111\]
+ net747 vssd1 vssd1 vccd1 vccd1 _04196_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout720_A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout341_X net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout439_X net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout818_A net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_34_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_168_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07508_ top.CPU.control_unit.instruction\[6\] net1278 vssd1 vssd1 vccd1 vccd1 _03147_
+ sky130_fd_sc_hd__nor2_1
XFILLER_23_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11779__A3 net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08488_ top.CPU.registers.data\[336\] net1321 net852 top.CPU.registers.data\[368\]
+ net770 vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__a221o_1
XFILLER_168_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07852__A1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_58 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout606_X net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12189__B1 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10450_ _05753_ _05866_ _05870_ _05981_ _06076_ vssd1 vssd1 vccd1 vccd1 _06077_ sky130_fd_sc_hd__a221o_1
XANTENNA__11936__B1 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09109_ _04744_ _04747_ net638 vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__a21o_1
X_10381_ net574 net520 _06010_ vssd1 vssd1 vccd1 vccd1 _06011_ sky130_fd_sc_hd__and3_1
XANTENNA__11400__A2 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12120_ top.CPU.registers.data\[92\] net657 net245 vssd1 vssd1 vccd1 vccd1 _06828_
+ sky130_fd_sc_hd__o21a_1
X_14155__325 clknet_leaf_134_clk vssd1 vssd1 vccd1 vccd1 net1794 sky130_fd_sc_hd__inv_2
XANTENNA_fanout975_X net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12051_ _06597_ _06779_ _06781_ net2867 vssd1 vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__a22o_1
Xhold380 top.CPU.registers.data\[5\] vssd1 vssd1 vccd1 vccd1 net2937 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold391 top.CPU.registers.data\[801\] vssd1 vssd1 vccd1 vccd1 net2948 sky130_fd_sc_hd__dlygate4sd3_1
X_11002_ net525 _06555_ vssd1 vssd1 vccd1 vccd1 _06556_ sky130_fd_sc_hd__nor2_2
XANTENNA__08565__C1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_1036 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07907__A2 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11096__D net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13365__S net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout860 net862 vssd1 vssd1 vccd1 vccd1 net860 sky130_fd_sc_hd__clkbuf_4
X_15810_ net2144 _02020_ net1174 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[610\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_70_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout871 net877 vssd1 vssd1 vccd1 vccd1 net871 sky130_fd_sc_hd__buf_8
Xfanout882 net883 vssd1 vssd1 vccd1 vccd1 net882 sky130_fd_sc_hd__clkbuf_4
Xfanout893 _02777_ vssd1 vssd1 vccd1 vccd1 net893 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15741_ net2075 _01951_ net1121 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[541\]
+ sky130_fd_sc_hd__dfrtp_1
X_12953_ top.CPU.alu.program_counter\[30\] _07392_ net1361 vssd1 vssd1 vccd1 vccd1
+ _01193_ sky130_fd_sc_hd__mux2_1
XANTENNA__11467__A2 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1080 top.CPU.registers.data\[367\] vssd1 vssd1 vccd1 vccd1 net3637 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08332__A2 net1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1091 top.CPU.registers.data\[943\] vssd1 vssd1 vccd1 vccd1 net3648 sky130_fd_sc_hd__dlygate4sd3_1
X_11904_ net3639 net186 net350 _05849_ vssd1 vssd1 vccd1 vccd1 _01662_ sky130_fd_sc_hd__a22o_1
X_15672_ net2006 _01882_ net1148 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[472\]
+ sky130_fd_sc_hd__dfrtp_1
X_12884_ _07310_ _07329_ _07317_ vssd1 vssd1 vccd1 vccd1 _07330_ sky130_fd_sc_hd__o21a_1
XFILLER_33_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07540__B1 _03118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13613__A0 top.CPU.alu.program_counter\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11835_ _06666_ net207 net155 net3073 vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__a22o_1
XANTENNA__11219__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12709__S net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_25_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07599__A net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ net466 _06609_ net239 net162 net3181 vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__a32o_1
XANTENNA__10737__B net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09832__A2 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13505_ top.CPU.data_out\[11\] net588 _02969_ _02972_ vssd1 vssd1 vccd1 vccd1 _02509_
+ sky130_fd_sc_hd__o22a_1
X_10717_ top.CPU.fetch.current_ra\[7\] net1040 net633 top.CPU.handler.toreg\[7\] vssd1
+ vssd1 vccd1 vccd1 _06332_ sky130_fd_sc_hd__a22o_2
X_11697_ _06527_ net207 net422 net2966 vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__a22o_1
X_16224_ clknet_leaf_30_clk _02434_ net1152 vssd1 vssd1 vccd1 vccd1 top.CPU.control_unit.instruction\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_13436_ _03200_ _03266_ _02935_ vssd1 vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__o21a_2
X_10648_ net416 _06264_ _06265_ vssd1 vssd1 vccd1 vccd1 _06266_ sky130_fd_sc_hd__o21a_1
XFILLER_139_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11927__B1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09596__A1 _05232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08399__A2 net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13392__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16155_ net2489 _02365_ net1214 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[955\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_154_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13367_ top.I2C.data_out\[16\] net556 _02893_ net597 vssd1 vssd1 vccd1 vccd1 _02894_
+ sky130_fd_sc_hd__a22o_1
X_10579_ net408 _06199_ vssd1 vssd1 vccd1 vccd1 _06200_ sky130_fd_sc_hd__or2_1
XANTENNA__10753__A _05672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09964__D _03650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14893__1063 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 net2532 sky130_fd_sc_hd__inv_2
XFILLER_115_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15438__RESET_B net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15106_ net1488 _01319_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r2_prev\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_170_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12318_ net2570 _03915_ net1227 vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_110_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16086_ net2420 _02296_ net1221 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[886\]
+ sky130_fd_sc_hd__dfrtp_1
X_13298_ top.mmio.mem_data_i\[30\] top.mmio.mem_data_i\[31\] top.mmio.mem_data_i\[28\]
+ top.mmio.mem_data_i\[29\] vssd1 vssd1 vccd1 vccd1 _02841_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_110_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09348__A1 _04986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15037_ clknet_leaf_89_clk _01282_ net1273 vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__dfrtp_1
X_12249_ net661 _06010_ net434 _06886_ vssd1 vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__a31o_1
XANTENNA__11287__C net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11155__B2 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08556__C1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10902__A1 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08571__A2 net1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13856__26 clknet_leaf_112_clk vssd1 vssd1 vccd1 vccd1 net1495 sky130_fd_sc_hd__inv_2
XANTENNA__08369__S net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07790_ top.CPU.registers.data\[606\] net1303 net1025 top.CPU.registers.data\[638\]
+ net944 vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__a221o_1
XANTENNA__12104__B1 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_147_Right_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_108_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15939_ net2273 _02149_ net1183 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[739\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11458__A2 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08323__A2 net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09989__A _04891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09460_ net795 _05093_ _05094_ net723 vssd1 vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__o211a_1
XFILLER_97_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_125_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16226__RESET_B net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08411_ _04049_ vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__inv_2
XFILLER_24_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09391_ top.CPU.registers.data\[227\] net1391 net828 top.CPU.registers.data\[195\]
+ net775 vssd1 vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__a221o_1
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10928__A net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_16_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__10418__B1 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12958__A2 _03409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08342_ net677 _03964_ _03965_ vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__and3_1
X_14596__766 clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 net2235 sky130_fd_sc_hd__inv_2
XFILLER_20_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08273_ top.CPU.registers.data_out_r2_prev\[22\] net687 net622 _03911_ vssd1 vssd1
+ vccd1 vccd1 _03912_ sky130_fd_sc_hd__o211a_1
XANTENNA__11630__A2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16615__A net1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout134_A _05990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09036__B1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08832__S net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11918__B1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14139__309 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 net1778 sky130_fd_sc_hd__inv_2
XANTENNA_fanout301_A _06604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1043_A _03165_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07598__B1 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_362 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08795__C1 net1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09339__A1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1210_A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11146__A1 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1308_A _03110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08547__C1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07972__A _03610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout123 net124 vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__clkbuf_4
XFILLER_114_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout134 _05990_ vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11697__A2 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout670_A net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout145 _06270_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__buf_2
XANTENNA_fanout291_X net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout156 net159 vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__clkbuf_8
Xfanout167 _06757_ vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout768_A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout178 _06795_ vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__buf_4
Xfanout189 net191 vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__buf_4
X_07988_ net953 _03625_ _03626_ net611 vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__a31o_1
XANTENNA__07770__B1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_114_Right_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09727_ _05332_ _05363_ vssd1 vssd1 vccd1 vccd1 _05366_ sky130_fd_sc_hd__nand2_2
XANTENNA_clkbuf_leaf_200_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout556_X net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12102__B net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout935_A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09899__A _04430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10657__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09658_ _04052_ _05296_ vssd1 vssd1 vccd1 vccd1 _05297_ sky130_fd_sc_hd__or2_2
X_14540__710 clknet_leaf_195_clk vssd1 vssd1 vccd1 vccd1 net2179 sky130_fd_sc_hd__inv_2
XFILLER_70_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10121__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08609_ net903 _04245_ _04247_ net1367 vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__a211o_1
X_13870__40 clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 net1509 sky130_fd_sc_hd__inv_2
XFILLER_82_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09589_ net1378 _03162_ vssd1 vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout723_X net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11620_ _06509_ net428 net206 net214 net2714 vssd1 vssd1 vccd1 vccd1 _01929_ sky130_fd_sc_hd__a32o_1
XFILLER_168_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09814__A2 net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11551_ net563 net526 _06528_ vssd1 vssd1 vccd1 vccd1 _06740_ sky130_fd_sc_hd__and3_1
XFILLER_156_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10502_ net1405 net576 net518 net139 vssd1 vssd1 vccd1 vccd1 _06127_ sky130_fd_sc_hd__and4_1
X_11482_ net485 net473 _06612_ net255 net3403 vssd1 vssd1 vccd1 vccd1 _02042_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_94_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11909__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13221_ _06948_ _02792_ vssd1 vssd1 vccd1 vccd1 _02794_ sky130_fd_sc_hd__nand2_1
X_10433_ _04193_ _05575_ vssd1 vssd1 vccd1 vccd1 _06060_ sky130_fd_sc_hd__or2_1
XANTENNA__13374__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12177__A3 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12264__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07589__B1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13152_ net1359 net126 _02742_ _02739_ top.CPU.alu.program_counter\[1\] vssd1 vssd1
+ vccd1 vccd1 _01298_ sky130_fd_sc_hd__a32o_1
X_10364_ _03923_ _05972_ net445 vssd1 vssd1 vccd1 vccd1 _05994_ sky130_fd_sc_hd__a21oi_1
XFILLER_124_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12103_ _06634_ _06770_ _06819_ net176 net3630 vssd1 vssd1 vccd1 vccd1 _01511_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_72_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_888 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13083_ top.CPU.data_out\[18\] net2751 net559 vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__mux2_1
XFILLER_2_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10295_ net550 _05367_ _05923_ net413 _05917_ vssd1 vssd1 vccd1 vccd1 _05928_ sky130_fd_sc_hd__o221a_1
XANTENNA__11137__A1 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07882__A net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08538__C1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12034_ top.CPU.registers.data\[142\] net649 net361 _06727_ vssd1 vssd1 vccd1 vccd1
+ _06792_ sky130_fd_sc_hd__o211a_1
XFILLER_104_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11608__S net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10896__B1 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout690 net691 vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__buf_4
XFILLER_92_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12012__B net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08305__A2 net1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12936_ _07375_ _07376_ vssd1 vssd1 vccd1 vccd1 _07377_ sky130_fd_sc_hd__and2b_1
X_15724_ net2058 _01934_ net1078 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[524\]
+ sky130_fd_sc_hd__dfrtp_1
X_14283__453 clknet_leaf_134_clk vssd1 vssd1 vccd1 vccd1 net1922 sky130_fd_sc_hd__inv_2
XFILLER_18_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12867_ _07313_ _07314_ vssd1 vssd1 vccd1 vccd1 _07315_ sky130_fd_sc_hd__nor2_1
X_15655_ net1989 _01865_ net1197 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[455\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11860__A2 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11818_ _06231_ net3847 net156 vssd1 vssd1 vccd1 vccd1 _01742_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13062__A1 top.CPU.data_out\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09266__B1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15586_ net1920 _01796_ net1172 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[386\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_159_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12798_ top.CPU.alu.program_counter\[16\] _04189_ vssd1 vssd1 vccd1 vccd1 _07252_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__08218__A _03822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10467__B _05680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09805__A2 net1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14324__494 clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 net1963 sky130_fd_sc_hd__inv_2
XANTENNA__07816__A1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11749_ net142 net534 net498 net192 net2660 vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__a32o_1
XFILLER_119_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12682__B _04919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09569__A1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13419_ _02830_ _02931_ vssd1 vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__nor2_1
X_16207_ net2541 _02417_ net1097 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[1007\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_128_896 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16138_ net2472 _02348_ net1084 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[938\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_154_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_149_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08792__A2 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08960_ _04594_ _04598_ net452 vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__mux2_1
X_16069_ net2403 _02279_ net1087 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[869\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_5_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_166_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07911_ top.CPU.registers.data\[252\] net1384 net995 top.CPU.registers.data\[220\]
+ net919 vssd1 vssd1 vccd1 vccd1 _03550_ sky130_fd_sc_hd__a221o_1
XFILLER_142_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08891_ _04528_ _04529_ net635 vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__a21o_1
XANTENNA__11679__A2 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10930__B _06354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07842_ top.CPU.registers.data\[157\] net979 _03480_ vssd1 vssd1 vccd1 vccd1 _03481_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__16407__RESET_B net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_162_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07773_ top.CPU.registers.data\[414\] net1303 net1025 top.CPU.registers.data\[446\]
+ vssd1 vssd1 vccd1 vccd1 _03412_ sky130_fd_sc_hd__a22o_1
XANTENNA__13825__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09512_ net629 _05149_ _05150_ net608 vssd1 vssd1 vccd1 vccd1 _05151_ sky130_fd_sc_hd__a31o_1
XFILLER_17_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08701__C1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09443_ net936 _05080_ _05081_ net954 vssd1 vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__o211a_1
XANTENNA__11761__B net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11851__A2 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout251_A _06733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout349_A net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09257__B1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09374_ net679 _04998_ _04999_ vssd1 vssd1 vccd1 vccd1 _05013_ sky130_fd_sc_hd__and3_1
XFILLER_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08325_ top.CPU.registers.data\[851\] net1294 net1015 top.CPU.registers.data\[883\]
+ net936 vssd1 vssd1 vccd1 vccd1 _03964_ sky130_fd_sc_hd__a221o_1
XFILLER_21_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1160_A net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout137_X net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout516_A net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1258_A net1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09009__B1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08256_ top.CPU.registers.data\[342\] net1307 net1030 top.CPU.registers.data\[374\]
+ net941 vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__a221o_1
XANTENNA__08480__A1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08187_ top.CPU.registers.data\[183\] net1014 net912 vssd1 vssd1 vccd1 vccd1 _03826_
+ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout304_X net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_81_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_104_Left_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08768__C1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08232__A1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout885_A _03095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11001__B net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11119__A1 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10590__A2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07991__B1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10080_ _04294_ _04363_ net378 vssd1 vssd1 vccd1 vccd1 _05718_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_96_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout673_X net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08940__C1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout840_X net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14267__437 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 net1906 sky130_fd_sc_hd__inv_2
XANTENNA_fanout938_X net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13643__S net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Left_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13770_ net29 net1051 net886 net3921 vssd1 vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__a22o_1
XANTENNA__08299__A1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10982_ net527 _06543_ vssd1 vssd1 vccd1 vccd1 _06544_ sky130_fd_sc_hd__nor2_1
XFILLER_90_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12767__B _04392_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12721_ top.CPU.alu.program_counter\[8\] _07182_ net1360 vssd1 vssd1 vccd1 vccd1
+ _01171_ sky130_fd_sc_hd__mux2_1
XANTENNA__09422__A net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14892__1062 clknet_leaf_189_clk vssd1 vssd1 vccd1 vccd1 net2531 sky130_fd_sc_hd__inv_2
XFILLER_55_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_154_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14011__181 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 net1650 sky130_fd_sc_hd__inv_2
XANTENNA__11842__A2 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12259__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14308__478 clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 net1947 sky130_fd_sc_hd__inv_2
X_15440_ net1774 _01650_ net1156 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[240\]
+ sky130_fd_sc_hd__dfrtp_1
X_12652_ _03138_ top.CPU.busy vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__nor2_1
XFILLER_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_34_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11603_ _05961_ net3399 net212 vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__mux2_1
XANTENNA__13595__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15371_ net1705 _01581_ net1064 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[171\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_168_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12583_ top.CPU.addressnew\[19\] top.CPU.addressnew\[18\] _07085_ _07086_ vssd1 vssd1
+ vccd1 vccd1 _07087_ sky130_fd_sc_hd__or4_1
XFILLER_129_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_169_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11534_ _06656_ net259 net250 net3197 vssd1 vssd1 vccd1 vccd1 _01997_ sky130_fd_sc_hd__a22o_1
XFILLER_12_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_122_Left_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13347__A2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_49_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11465_ net492 net477 _06592_ net266 net3019 vssd1 vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__a32o_1
XFILLER_99_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13204_ top.I2C.within_byte_counter_reading\[1\] top.I2C.within_byte_counter_reading\[0\]
+ top.I2C.within_byte_counter_reading\[2\] vssd1 vssd1 vccd1 vccd1 _02782_ sky130_fd_sc_hd__or3b_2
X_10416_ _06043_ vssd1 vssd1 vccd1 vccd1 _06044_ sky130_fd_sc_hd__inv_2
XANTENNA__09420__B1 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11396_ _06522_ net276 net271 net3593 vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__a22o_1
XFILLER_124_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13135_ net2700 _02736_ _02734_ vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__mux2_1
XFILLER_48_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08774__A2 net1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10347_ net404 _05977_ vssd1 vssd1 vccd1 vccd1 _05978_ sky130_fd_sc_hd__nand2_1
XFILLER_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_92 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13066_ top.CPU.data_out\[1\] net2669 net560 vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__mux2_1
X_10278_ _05332_ _05467_ net379 vssd1 vssd1 vccd1 vccd1 _05911_ sky130_fd_sc_hd__mux2_1
XFILLER_140_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09184__C1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09723__A1 top.CPU.control_unit.instruction\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12017_ net3778 net151 _06785_ vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__a21o_1
XANTENNA__08526__A2 net1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_107_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10869__B1 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08995__X _04634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08931__C1 net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_105_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12086__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14946__Q top.CPU.alu.program_counter\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10097__B2 _03409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15707_ net2041 _01917_ net1213 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[507\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11581__B _06731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11294__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12919_ top.CPU.alu.program_counter\[27\] top.CPU.alu.program_counter\[26\] _07337_
+ vssd1 vssd1 vccd1 vccd1 _07362_ sky130_fd_sc_hd__and3_1
XFILLER_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09239__B1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15638_ net1972 _01848_ net1228 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[438\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_148_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12693__A top.CPU.alu.program_counter\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15569_ net1903 _01779_ net1189 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[369\]
+ sky130_fd_sc_hd__dfrtp_1
X_08110_ net798 _03747_ _03748_ net728 vssd1 vssd1 vccd1 vccd1 _03749_ sky130_fd_sc_hd__o211a_1
XANTENNA__08998__C1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09090_ _04727_ _04728_ net452 vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__mux2_1
XANTENNA__10925__B _06472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08041_ top.CPU.control_unit.instruction\[16\] _03672_ net641 vssd1 vssd1 vccd1 vccd1
+ _03680_ sky130_fd_sc_hd__a21oi_1
XFILLER_31_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11102__A net1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold902 top.CPU.registers.data\[795\] vssd1 vssd1 vccd1 vccd1 net3459 sky130_fd_sc_hd__dlygate4sd3_1
Xhold913 top.CPU.registers.data\[770\] vssd1 vssd1 vccd1 vccd1 net3470 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09411__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold924 top.CPU.registers.data\[286\] vssd1 vssd1 vccd1 vccd1 net3481 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_127_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_6_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold935 top.CPU.registers.data\[463\] vssd1 vssd1 vccd1 vccd1 net3492 sky130_fd_sc_hd__dlygate4sd3_1
Xhold946 top.CPU.registers.data\[607\] vssd1 vssd1 vccd1 vccd1 net3503 sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 top.CPU.registers.data\[896\] vssd1 vssd1 vccd1 vccd1 net3514 sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 top.CPU.registers.data\[601\] vssd1 vssd1 vccd1 vccd1 net3525 sky130_fd_sc_hd__dlygate4sd3_1
X_09992_ _05627_ _05630_ net381 vssd1 vssd1 vccd1 vccd1 _05631_ sky130_fd_sc_hd__mux2_1
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold979 net65 vssd1 vssd1 vccd1 vccd1 net3536 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_164_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10572__A2 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08943_ net928 _04580_ _04581_ net951 vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__o211a_1
XFILLER_130_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08411__A _04049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_15_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_15_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout299_A _06645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09714__A1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08874_ net784 _04511_ _04512_ net714 vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__o211a_1
XFILLER_56_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1006_A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08922__C1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07825_ top.CPU.registers.data\[253\] net1389 net816 top.CPU.registers.data\[221\]
+ net768 vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout466_A net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07756_ top.CPU.registers.data\[478\] net1333 net864 top.CPU.registers.data\[510\]
+ net778 vssd1 vssd1 vccd1 vccd1 _03395_ sky130_fd_sc_hd__a221o_1
XANTENNA__10659__Y _06276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07687_ _03271_ _03314_ _03284_ _03304_ vssd1 vssd1 vccd1 vccd1 _03326_ sky130_fd_sc_hd__and4bb_1
XANTENNA_fanout633_A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout254_X net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1375_A net1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09426_ top.CPU.registers.data\[66\] net1294 net1015 top.CPU.registers.data\[98\]
+ net954 vssd1 vssd1 vccd1 vccd1 _05065_ sky130_fd_sc_hd__a221o_1
X_13840__10 clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 net1479 sky130_fd_sc_hd__inv_2
X_09357_ top.CPU.registers.data\[835\] net1297 net1018 top.CPU.registers.data\[867\]
+ net939 vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__a221o_1
XANTENNA__09896__B _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout421_X net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout800_A net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout519_X net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08989__C1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09388__S net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08308_ top.CPU.registers.data\[563\] top.CPU.registers.data\[531\] net826 vssd1
+ vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09288_ top.CPU.registers.data\[964\] net1299 net1020 top.CPU.registers.data\[996\]
+ net918 vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__a221o_1
XFILLER_166_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14652__822 clknet_leaf_137_clk vssd1 vssd1 vccd1 vccd1 net2291 sky130_fd_sc_hd__inv_2
XFILLER_126_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07504__1 clknet_leaf_183_clk vssd1 vssd1 vccd1 vccd1 net1470 sky130_fd_sc_hd__inv_2
XFILLER_126_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08239_ top.CPU.registers.data\[662\] net1334 net866 top.CPU.registers.data\[694\]
+ net731 vssd1 vssd1 vccd1 vccd1 _03878_ sky130_fd_sc_hd__a221o_1
XFILLER_138_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1330_X net1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11012__A net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08205__A1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11250_ net2820 net293 _06680_ net481 vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__a22o_1
XFILLER_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09402__B1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12001__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout790_X net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10012__A1 _03544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10201_ _05718_ _05724_ net306 vssd1 vssd1 vccd1 vccd1 _05837_ sky130_fd_sc_hd__mux2_1
XANTENNA__13638__S net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11181_ _06035_ net430 vssd1 vssd1 vccd1 vccd1 _06650_ sky130_fd_sc_hd__and2_1
XFILLER_69_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07964__B1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09417__A net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10132_ top.CPU.fetch.current_ra\[30\] net1042 vssd1 vssd1 vccd1 vccd1 _05770_ sky130_fd_sc_hd__and2_1
XFILLER_122_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10570__B _06190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12114__Y _06825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_89_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14940_ clknet_leaf_72_clk _01186_ net1158 vssd1 vssd1 vccd1 vccd1 top.CPU.alu.program_counter\[23\]
+ sky130_fd_sc_hd__dfrtp_4
X_10063_ _05192_ net372 vssd1 vssd1 vccd1 vccd1 _05701_ sky130_fd_sc_hd__nor2_1
XANTENNA__12170__D1 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09181__A2 net1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input27_A DAT_I[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13822_ net3496 net337 net329 top.CPU.data_out\[24\] vssd1 vssd1 vccd1 vccd1 _02702_
+ sky130_fd_sc_hd__a22o_1
XFILLER_75_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13265__B2 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16541_ clknet_leaf_85_clk net3691 net1266 vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__dfrtp_1
X_13753_ net2630 _03087_ vssd1 vssd1 vccd1 vccd1 _02642_ sky130_fd_sc_hd__xnor2_1
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10965_ net530 _05933_ net541 vssd1 vssd1 vccd1 vccd1 _06534_ sky130_fd_sc_hd__nor3_2
X_12704_ top.CPU.alu.program_counter\[7\] _04793_ vssd1 vssd1 vccd1 vccd1 _07167_
+ sky130_fd_sc_hd__nor2_1
X_16472_ clknet_leaf_88_clk _02634_ net1274 vssd1 vssd1 vccd1 vccd1 top.SPI.timem\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13684_ net2649 net332 vssd1 vssd1 vccd1 vccd1 _02612_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_100_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10896_ net484 net460 _06491_ net221 net3103 vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_100_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12635_ top.I2C.output_state\[14\] net3626 vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__and2_1
X_15423_ net1757 _01633_ net1221 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[223\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_130_Left_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11621__S net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15354_ net1688 _01564_ net1251 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[154\]
+ sky130_fd_sc_hd__dfrtp_1
X_12566_ _06309_ _06331_ _06352_ _07070_ vssd1 vssd1 vccd1 vccd1 _07071_ sky130_fd_sc_hd__or4b_1
XFILLER_7_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14395__565 clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 net2034 sky130_fd_sc_hd__inv_2
X_11517_ net489 net136 net356 net252 net2945 vssd1 vssd1 vccd1 vccd1 _02013_ sky130_fd_sc_hd__a32o_1
XANTENNA__10237__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15285_ net1619 _01495_ net1210 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[85\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_144_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12497_ _05154_ _05190_ _05227_ _05265_ vssd1 vssd1 vccd1 vccd1 _07006_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_156_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold209 top.CPU.registers.data\[418\] vssd1 vssd1 vccd1 vccd1 net2766 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11448_ _06056_ net3856 net263 vssd1 vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__mux2_1
XFILLER_109_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11200__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10761__A net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11379_ _06494_ net281 net273 net3092 vssd1 vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__a22o_1
XFILLER_4_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07955__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13118_ top.SPI.command\[5\] net1410 top.SPI.paroutput\[29\] net1358 vssd1 vssd1
+ vccd1 vccd1 _02724_ sky130_fd_sc_hd__a22o_1
XANTENNA__10480__B net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_1012 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13049_ top.SPI.parameters\[26\] top.SPI.paroutput\[18\] net1357 vssd1 vssd1 vccd1
+ vccd1 _07450_ sky130_fd_sc_hd__mux2_1
XFILLER_140_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1260 net1262 vssd1 vssd1 vccd1 vccd1 net1260 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09761__S net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1271 net1275 vssd1 vssd1 vccd1 vccd1 net1271 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09172__A2 net1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1282 _03115_ vssd1 vssd1 vccd1 vccd1 net1282 sky130_fd_sc_hd__buf_4
XANTENNA__12688__A top.CPU.alu.program_counter\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1293 _03113_ vssd1 vssd1 vccd1 vccd1 net1293 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08380__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07610_ top.CPU.control_unit.instruction\[14\] net1398 vssd1 vssd1 vccd1 vccd1 _03249_
+ sky130_fd_sc_hd__or2_1
XANTENNA__11592__A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08590_ net1367 _04228_ vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__or2_1
XFILLER_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13256__B2 _02803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07541_ top.CPU.control_unit.instruction\[7\] net1407 net662 vssd1 vssd1 vccd1 vccd1
+ _03180_ sky130_fd_sc_hd__o21a_4
XFILLER_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12200__B net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08132__B1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08683__A1 _03116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07472_ top.CPU.control_unit.instruction\[18\] vssd1 vssd1 vccd1 vccd1 _03112_ sky130_fd_sc_hd__inv_2
XFILLER_14_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09211_ top.CPU.registers.data\[230\] net1379 net978 top.CPU.registers.data\[198\]
+ net904 vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__a221o_1
XFILLER_14_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14636__806 clknet_leaf_189_clk vssd1 vssd1 vccd1 vccd1 net2275 sky130_fd_sc_hd__inv_2
XFILLER_50_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10936__A net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire591_X net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09142_ net943 _04779_ _04780_ net958 vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_174_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12231__A2 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11034__A3 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09001__S net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09073_ net617 _04704_ _04711_ net611 vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__o211a_1
XFILLER_163_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout214_A _06752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08024_ net791 _03652_ _03653_ net719 vssd1 vssd1 vccd1 vccd1 _03663_ sky130_fd_sc_hd__o211a_1
XANTENNA__08840__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold710 top.CPU.registers.data\[720\] vssd1 vssd1 vccd1 vccd1 net3267 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12870__B _03823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold721 top.CPU.registers.data\[498\] vssd1 vssd1 vccd1 vccd1 net3278 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10942__Y _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold732 top.CPU.registers.data\[42\] vssd1 vssd1 vccd1 vccd1 net3289 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08199__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13458__S net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold743 top.CPU.registers.data\[197\] vssd1 vssd1 vccd1 vccd1 net3300 sky130_fd_sc_hd__dlygate4sd3_1
X_14891__1061 clknet_leaf_148_clk vssd1 vssd1 vccd1 vccd1 net2530 sky130_fd_sc_hd__inv_2
XFILLER_162_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold754 top.CPU.registers.data\[276\] vssd1 vssd1 vccd1 vccd1 net3311 sky130_fd_sc_hd__dlygate4sd3_1
Xhold765 top.CPU.registers.data\[512\] vssd1 vssd1 vccd1 vccd1 net3322 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10545__A2 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold776 top.CPU.registers.data\[891\] vssd1 vssd1 vccd1 vccd1 net3333 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11742__A1 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07946__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold787 top.CPU.registers.data\[702\] vssd1 vssd1 vccd1 vccd1 net3344 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09975_ _05524_ _05613_ _03444_ vssd1 vssd1 vccd1 vccd1 _05614_ sky130_fd_sc_hd__a21o_1
Xhold798 top.CPU.registers.data\[696\] vssd1 vssd1 vccd1 vccd1 net3355 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09148__C1 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08926_ net641 _04561_ _04564_ net703 _04558_ vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__o311a_1
XFILLER_130_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13495__A1 net1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12298__A2 _06887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09699__B1 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1410 top.SPI.paroutput\[20\] vssd1 vssd1 vccd1 vccd1 net3967 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09671__S net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1009_X net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1421 top.CPU.handler.toreg\[28\] vssd1 vssd1 vccd1 vccd1 net3978 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1432 top.I2C.within_byte_counter_writing\[1\] vssd1 vssd1 vccd1 vccd1 net3989
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08857_ net617 _04495_ _04490_ net611 vssd1 vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__o211a_1
Xhold1443 top.SPI.busy vssd1 vssd1 vccd1 vccd1 net4000 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout371_X net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout750_A net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1454 top.SPI.count\[1\] vssd1 vssd1 vccd1 vccd1 net4011 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1465 top.CPU.fetch.current_ra\[23\] vssd1 vssd1 vccd1 vccd1 net4022 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout469_X net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout848_A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07808_ top.CPU.registers.data\[925\] net1319 net850 top.CPU.registers.data\[957\]
+ net692 vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__a221o_1
XANTENNA__08287__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08788_ top.CPU.registers.data_out_r1_prev\[12\] net871 net641 _04411_ _04426_ vssd1
+ vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__o221ai_4
X_07739_ net700 _03377_ vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout1280_X net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08123__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout636_X net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1378_X net1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11007__A net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10750_ net389 _06362_ _06360_ net406 vssd1 vssd1 vccd1 vccd1 _06363_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_45_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14082__252 clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 net1721 sky130_fd_sc_hd__inv_2
X_09409_ net751 _05046_ _05047_ net696 vssd1 vssd1 vccd1 vccd1 _05048_ sky130_fd_sc_hd__o211a_1
XFILLER_158_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10681_ net400 _06296_ vssd1 vssd1 vccd1 vccd1 _06297_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout803_X net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14379__549 clknet_leaf_135_clk vssd1 vssd1 vccd1 vccd1 net2018 sky130_fd_sc_hd__inv_2
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12420_ net1354 top.SPI.state\[5\] vssd1 vssd1 vccd1 vccd1 _06946_ sky130_fd_sc_hd__nand2_2
XANTENNA__12222__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12351_ net37 net3892 net898 net1054 net3975 vssd1 vssd1 vccd1 vccd1 _00064_ sky130_fd_sc_hd__a32o_1
XANTENNA__16306__Q top.CPU.data_out\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14123__293 clknet_leaf_148_clk vssd1 vssd1 vccd1 vccd1 net1762 sky130_fd_sc_hd__inv_2
XFILLER_126_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11302_ net475 net520 _05694_ _06487_ vssd1 vssd1 vccd1 vccd1 _06708_ sky130_fd_sc_hd__and4_1
XANTENNA__09846__S net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15070_ clknet_leaf_49_clk _00048_ net1129 vssd1 vssd1 vccd1 vccd1 top.I2C.output_state\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12282_ net2599 _03611_ net1150 vssd1 vssd1 vccd1 vccd1 _01399_ sky130_fd_sc_hd__mux2_1
XANTENNA__09387__C1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11233_ net2833 net295 _06671_ net488 vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__a22o_1
XANTENNA__10581__A _06141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07937__B1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11164_ net566 net517 vssd1 vssd1 vccd1 vccd1 _06643_ sky130_fd_sc_hd__nor2_1
XFILLER_106_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10115_ net409 _05643_ vssd1 vssd1 vccd1 vccd1 _05753_ sky130_fd_sc_hd__nor2_2
XFILLER_122_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13486__A1 _05226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15972_ net2306 _02182_ net1186 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[772\]
+ sky130_fd_sc_hd__dfrtp_1
X_11095_ net496 net469 _06605_ net304 net2806 vssd1 vssd1 vccd1 vccd1 _02305_ sky130_fd_sc_hd__a32o_1
XANTENNA__08986__A net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_720 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14780__950 clknet_leaf_136_clk vssd1 vssd1 vccd1 vccd1 net2419 sky130_fd_sc_hd__inv_2
X_10046_ _03306_ _03310_ _03323_ _03329_ vssd1 vssd1 vccd1 vccd1 _05685_ sky130_fd_sc_hd__a31oi_4
X_14923_ clknet_leaf_30_clk _01169_ net1152 vssd1 vssd1 vccd1 vccd1 top.CPU.alu.program_counter\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11497__B1 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold70 top.I2C.I2C_state\[6\] vssd1 vssd1 vccd1 vccd1 net2627 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08362__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold81 net49 vssd1 vssd1 vccd1 vccd1 net2638 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11616__S net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold92 net47 vssd1 vssd1 vccd1 vccd1 net2649 sky130_fd_sc_hd__dlygate4sd3_1
X_13805_ net3641 net333 net326 net3532 vssd1 vssd1 vccd1 vccd1 _02685_ sky130_fd_sc_hd__a22o_1
X_14821__991 clknet_leaf_110_clk vssd1 vssd1 vccd1 vccd1 net2460 sky130_fd_sc_hd__inv_2
XANTENNA__13789__A2 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11997_ _06564_ net341 net180 net3551 vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__a22o_1
XFILLER_63_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13987__157 clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 net1626 sky130_fd_sc_hd__inv_2
XANTENNA__08114__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10459__C net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09311__C1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16524_ clknet_leaf_100_clk _02686_ net1255 vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__dfrtp_1
XFILLER_91_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13736_ _03076_ _03077_ vssd1 vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_27_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10948_ net1406 _03170_ vssd1 vssd1 vccd1 vccd1 _06523_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_27_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12955__B net1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09610__A net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16455_ clknet_leaf_86_clk _02618_ net1265 vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__dfrtp_1
XFILLER_149_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13667_ net2795 net331 net330 top.CPU.addressnew\[0\] vssd1 vssd1 vccd1 vccd1 _02595_
+ sky130_fd_sc_hd__a22o_1
X_10879_ net521 _05693_ _06479_ vssd1 vssd1 vccd1 vccd1 _06481_ sky130_fd_sc_hd__and3_1
X_15406_ net1740 _01616_ net1105 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[206\]
+ sky130_fd_sc_hd__dfrtp_1
X_12618_ top.SPI.state\[3\] top.SPI.state\[4\] top.SPI.register\[1\] vssd1 vssd1 vccd1
+ vccd1 _07116_ sky130_fd_sc_hd__o21a_1
X_16386_ clknet_leaf_89_clk _00071_ net1273 vssd1 vssd1 vccd1 vccd1 top.SPI.state\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_13598_ net1349 _06067_ _06081_ _03025_ vssd1 vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__a31o_1
XANTENNA__09614__B1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12213__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12549_ top.CPU.handler.state\[5\] _03152_ _07055_ _07057_ net3998 vssd1 vssd1 vccd1
+ vccd1 _07058_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_117_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15337_ net1671 _01547_ net1060 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[137\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11421__B1 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09090__A1 _04728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1 _03047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15268_ net1602 _01478_ net1185 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[68\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09917__B2 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15199_ clknet_leaf_87_clk _01409_ net1271 vssd1 vssd1 vccd1 vccd1 top.SPI.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_113_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09393__A2 net1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout508 net510 vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_130_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout519 net522 vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__clkbuf_4
XFILLER_99_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09760_ net1037 net448 _05398_ vssd1 vssd1 vccd1 vccd1 _05399_ sky130_fd_sc_hd__a21oi_4
XANTENNA__12910__S net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13477__A1 net1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08711_ net784 _04349_ vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__or2_1
XANTENNA__11488__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13931__101 clknet_leaf_135_clk vssd1 vssd1 vccd1 vccd1 net1570 sky130_fd_sc_hd__inv_2
X_09691_ _05308_ _05316_ _05329_ vssd1 vssd1 vccd1 vccd1 _05330_ sky130_fd_sc_hd__a21oi_4
Xfanout1090 net1093 vssd1 vssd1 vccd1 vccd1 net1090 sky130_fd_sc_hd__clkbuf_4
X_08642_ net793 _04279_ _04280_ net744 vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__o211a_1
XFILLER_82_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10160__B1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_159_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08573_ top.CPU.registers.data\[911\] net1314 net846 top.CPU.registers.data\[943\]
+ net716 vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__a221o_1
XANTENNA__16618__A net1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout164_A _06757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08105__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14066__236 clknet_leaf_193_clk vssd1 vssd1 vccd1 vccd1 net1705 sky130_fd_sc_hd__inv_2
X_07524_ net1279 _03153_ _03157_ _03144_ vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__a22oi_4
XFILLER_25_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09520__A top.CPU.alu.program_counter\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11660__B1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07864__C1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout331_A net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout429_A _06642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1073_A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08408__A1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14107__277 clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 net1746 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_40_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12204__A2 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09125_ _04763_ vssd1 vssd1 vccd1 vccd1 _04764_ sky130_fd_sc_hd__inv_2
XANTENNA__11412__B1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09081__A1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12881__A top.CPU.alu.program_counter\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1240_A net1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout217_X net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1338_A _03109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09056_ net702 _04690_ _04692_ _04693_ _04694_ vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__o32a_1
XFILLER_135_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08007_ top.CPU.control_unit.instruction\[24\] net1046 _03408_ vssd1 vssd1 vccd1
+ vccd1 _03646_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout798_A net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold540 top.SPI.counter\[0\] vssd1 vssd1 vccd1 vccd1 net3097 sky130_fd_sc_hd__dlygate4sd3_1
Xhold551 top.CPU.registers.data\[878\] vssd1 vssd1 vccd1 vccd1 net3108 sky130_fd_sc_hd__dlygate4sd3_1
Xhold562 top.CPU.registers.data\[188\] vssd1 vssd1 vccd1 vccd1 net3119 sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 top.CPU.registers.data\[968\] vssd1 vssd1 vccd1 vccd1 net3130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold584 top.CPU.registers.data\[13\] vssd1 vssd1 vccd1 vccd1 net3141 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold595 top.CPU.registers.data\[456\] vssd1 vssd1 vccd1 vccd1 net3152 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout965_A net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14764__934 clknet_leaf_191_clk vssd1 vssd1 vccd1 vccd1 net2403 sky130_fd_sc_hd__inv_2
XFILLER_1_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11191__A2 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12820__S net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09958_ _05332_ _05364_ _05367_ _05529_ vssd1 vssd1 vccd1 vccd1 _05597_ sky130_fd_sc_hd__a22o_1
XANTENNA__09136__A2 net1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08909_ top.CPU.registers.data\[74\] net1313 net844 top.CPU.registers.data\[106\]
+ net765 vssd1 vssd1 vccd1 vccd1 _04548_ sky130_fd_sc_hd__a221o_1
XANTENNA__11479__B1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11944__B net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout753_X net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09889_ _05500_ _05467_ vssd1 vssd1 vccd1 vccd1 _05528_ sky130_fd_sc_hd__and2b_1
Xhold1240 top.I2C.data_out\[21\] vssd1 vssd1 vccd1 vccd1 net3797 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1251 top.CPU.registers.data_out_r1_prev\[23\] vssd1 vssd1 vccd1 vccd1 net3808
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14805__975 clknet_leaf_172_clk vssd1 vssd1 vccd1 vccd1 net2444 sky130_fd_sc_hd__inv_2
XANTENNA__09541__C1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1262 top.CPU.registers.data\[650\] vssd1 vssd1 vccd1 vccd1 net3819 sky130_fd_sc_hd__dlygate4sd3_1
X_11920_ net3787 net184 net344 _06233_ vssd1 vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__a22o_1
XANTENNA__07698__A2 _03154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1273 top.CPU.registers.data\[544\] vssd1 vssd1 vccd1 vccd1 net3830 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1284 top.wm.curr_state\[2\] vssd1 vssd1 vccd1 vccd1 net3841 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1295 top.SPI.dcx vssd1 vssd1 vccd1 vccd1 net3852 sky130_fd_sc_hd__dlygate4sd3_1
X_11851_ _06684_ net234 net152 net2698 vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout920_X net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13651__S net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10802_ net1406 net577 net517 net148 vssd1 vssd1 vccd1 vccd1 _06413_ sky130_fd_sc_hd__and4_1
X_11782_ _06627_ net196 net160 net3387 vssd1 vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__a22o_1
XFILLER_54_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10454__A1 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13521_ _03984_ net584 vssd1 vssd1 vccd1 vccd1 _02981_ sky130_fd_sc_hd__and2_1
X_10733_ net416 _06340_ _06341_ _06346_ vssd1 vssd1 vccd1 vccd1 _06347_ sky130_fd_sc_hd__a22o_1
XFILLER_158_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07855__C1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11651__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12267__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08742__S1 net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13452_ net3981 _02947_ net123 vssd1 vssd1 vccd1 vccd1 _02481_ sky130_fd_sc_hd__mux2_1
X_16240_ clknet_leaf_45_clk _02450_ net1138 vssd1 vssd1 vccd1 vccd1 top.CPU.control_unit.instruction\[16\]
+ sky130_fd_sc_hd__dfrtp_4
X_10664_ net397 _06279_ _06280_ net402 vssd1 vssd1 vccd1 vccd1 _06281_ sky130_fd_sc_hd__o211a_1
XFILLER_139_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_14_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12403_ _03120_ top.I2C.I2C_state\[11\] net2565 vssd1 vssd1 vccd1 vccd1 _00028_ sky130_fd_sc_hd__a21o_1
XANTENNA__10206__A1 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11403__B1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13383_ net1379 _02905_ net668 vssd1 vssd1 vccd1 vccd1 _02454_ sky130_fd_sc_hd__mux2_1
X_16171_ net2505 _02381_ net1057 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[971\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09072__A1 net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10595_ _04469_ _05284_ net446 vssd1 vssd1 vccd1 vccd1 _06215_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_97_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09576__S net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11954__A1 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15122_ clknet_leaf_50_clk _01334_ net1130 vssd1 vssd1 vccd1 vccd1 top.I2C.within_byte_counter_reading\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_11_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12334_ net2575 _04855_ net1080 vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__mux2_1
XFILLER_127_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15053_ clknet_leaf_73_clk _01298_ net1158 vssd1 vssd1 vccd1 vccd1 top.CPU.alu.program_counter\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_142_728 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12265_ net2984 _06354_ net432 vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__mux2_1
XANTENNA__10509__A2 _05939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_128_Right_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11216_ net530 net138 net545 vssd1 vssd1 vccd1 vccd1 _06663_ sky130_fd_sc_hd__and3_1
XANTENNA__08032__C1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12196_ net566 net363 _06673_ net170 top.CPU.registers.data\[53\] vssd1 vssd1 vccd1
+ vccd1 _06865_ sky130_fd_sc_hd__a32o_1
Xoutput60 net60 vssd1 vssd1 vccd1 vccd1 ADR_O[3] sky130_fd_sc_hd__buf_2
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 DAT_O[12] sky130_fd_sc_hd__buf_2
XANTENNA__11182__A2 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput82 net82 vssd1 vssd1 vccd1 vccd1 DAT_O[22] sky130_fd_sc_hd__buf_2
Xoutput93 net93 vssd1 vssd1 vccd1 vccd1 DAT_O[3] sky130_fd_sc_hd__buf_2
XFILLER_122_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09780__C1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11147_ net515 _06356_ vssd1 vssd1 vccd1 vccd1 _06633_ sky130_fd_sc_hd__nor2_1
XANTENNA__12730__S net1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13459__A1 net1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09127__A2 net1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07824__S net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15955_ net2289 _02165_ net1184 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[755\]
+ sky130_fd_sc_hd__dfrtp_1
X_11078_ net3697 net366 _06594_ net311 vssd1 vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__a22o_1
XANTENNA__09532__C1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10029_ _05663_ _05667_ vssd1 vssd1 vccd1 vccd1 _05668_ sky130_fd_sc_hd__nor2_1
XFILLER_64_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15886_ net2220 _02096_ net1193 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[686\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_64_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10693__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11890__B1 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08099__C1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14890__1060 clknet_leaf_151_clk vssd1 vssd1 vccd1 vccd1 net2529 sky130_fd_sc_hd__inv_2
XANTENNA__09835__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16507_ clknet_leaf_49_clk _02669_ net1128 vssd1 vssd1 vccd1 vccd1 top.mmio.mem_data_i\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_13719_ net4013 _03064_ _07113_ vssd1 vssd1 vccd1 vccd1 _03067_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11642__B1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16438_ clknet_leaf_80_clk _02601_ net1242 vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__dfrtp_1
XFILLER_32_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07861__A2 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16369_ clknet_leaf_70_clk _02578_ net1169 vssd1 vssd1 vccd1 vccd1 top.CPU.fetch.current_ra\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11945__A1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13147__B1 net1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14451__621 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 net2090 sky130_fd_sc_hd__inv_2
XFILLER_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14748__918 clknet_leaf_136_clk vssd1 vssd1 vccd1 vccd1 net2387 sky130_fd_sc_hd__inv_2
XFILLER_126_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11110__A net1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09366__A2 net1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout305 net307 vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__clkbuf_4
XFILLER_99_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout316 net322 vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__buf_4
Xfanout327 net328 vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09771__C1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09812_ top.CPU.registers.data_out_r1_prev\[26\] net876 _05440_ _05443_ vssd1 vssd1
+ vccd1 vccd1 _05451_ sky130_fd_sc_hd__o22a_1
Xfanout338 _03047_ vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__buf_2
XFILLER_141_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout349 net353 vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__buf_2
XFILLER_86_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10920__A2 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09743_ net797 _05380_ _05381_ net751 vssd1 vssd1 vccd1 vccd1 _05382_ sky130_fd_sc_hd__o211a_1
XANTENNA__08326__B1 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout281_A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout379_A net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09674_ top.CPU.registers.data\[441\] top.CPU.registers.data\[409\] net837 vssd1
+ vssd1 vccd1 vccd1 _05313_ sky130_fd_sc_hd__mux2_1
XFILLER_55_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10133__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08625_ top.CPU.registers.data\[750\] net1390 net818 top.CPU.registers.data\[718\]
+ net720 vssd1 vssd1 vccd1 vccd1 _04264_ sky130_fd_sc_hd__a221o_1
XANTENNA__11881__A0 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12876__A top.CPU.alu.program_counter\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout546_A _06523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout167_X net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1288_A net1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08556_ top.CPU.registers.data\[239\] net1387 net812 top.CPU.registers.data\[207\]
+ net717 vssd1 vssd1 vccd1 vccd1 _04195_ sky130_fd_sc_hd__a221o_1
XANTENNA__08629__A1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10667__Y _06284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07507_ top.CPU.control_unit.instruction\[3\] top.CPU.control_unit.instruction\[2\]
+ top.CPU.control_unit.instruction\[0\] top.CPU.control_unit.instruction\[1\] vssd1
+ vssd1 vccd1 vccd1 _03146_ sky130_fd_sc_hd__or4bb_1
XFILLER_52_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11633__B1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08487_ top.CPU.registers.data\[304\] top.CPU.registers.data\[272\] net821 vssd1
+ vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout713_A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12189__A1 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11004__B net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout501_X net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13500__A _04656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09108_ net700 _04745_ _04746_ vssd1 vssd1 vccd1 vccd1 _04747_ sky130_fd_sc_hd__or3_1
XFILLER_148_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10380_ net601 _06008_ _06009_ vssd1 vssd1 vccd1 vccd1 _06010_ sky130_fd_sc_hd__a21o_4
XFILLER_164_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09039_ net740 _04671_ _04670_ net766 vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout1410_X net1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14194__364 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 net1833 sky130_fd_sc_hd__inv_2
XFILLER_151_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11020__A net1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09357__A2 net1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12050_ net3829 net655 _06794_ vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_92_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold370 net91 vssd1 vssd1 vccd1 vccd1 net2927 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08014__C1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold381 top.CPU.registers.data\[639\] vssd1 vssd1 vccd1 vccd1 net2938 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout870_X net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11001_ net540 net501 _06271_ vssd1 vssd1 vccd1 vccd1 _06555_ sky130_fd_sc_hd__or3b_1
Xhold392 top.CPU.registers.data\[827\] vssd1 vssd1 vccd1 vccd1 net2949 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13646__S net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09762__C1 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout850 net854 vssd1 vssd1 vccd1 vccd1 net850 sky130_fd_sc_hd__clkbuf_4
Xfanout861 net862 vssd1 vssd1 vccd1 vccd1 net861 sky130_fd_sc_hd__buf_2
Xfanout872 net873 vssd1 vssd1 vccd1 vccd1 net872 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout883 _03166_ vssd1 vssd1 vccd1 vccd1 net883 sky130_fd_sc_hd__buf_2
Xfanout894 net896 vssd1 vssd1 vccd1 vccd1 net894 sky130_fd_sc_hd__clkbuf_4
XFILLER_92_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15740_ net2074 _01950_ net1235 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[540\]
+ sky130_fd_sc_hd__dfrtp_1
X_12952_ _07391_ _07387_ net128 vssd1 vssd1 vccd1 vccd1 _07392_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1070 top.CPU.handler.toreg\[6\] vssd1 vssd1 vccd1 vccd1 net3627 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1081 top.CPU.registers.data\[335\] vssd1 vssd1 vccd1 vccd1 net3638 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1092 top.CPU.registers.data\[323\] vssd1 vssd1 vccd1 vccd1 net3649 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11903_ net3721 net184 net344 _05811_ vssd1 vssd1 vccd1 vccd1 _01663_ sky130_fd_sc_hd__a22o_1
XFILLER_18_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15671_ net2005 _01881_ net1181 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[471\]
+ sky130_fd_sc_hd__dfrtp_1
X_12883_ top.CPU.alu.program_counter\[23\] _03823_ _03916_ top.CPU.alu.program_counter\[22\]
+ vssd1 vssd1 vccd1 vccd1 _07329_ sky130_fd_sc_hd__a22o_1
XFILLER_73_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11834_ _06665_ net235 net153 net3063 vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__a22o_1
XANTENNA__09817__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11624__A0 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11765_ _06608_ net206 net163 net3370 vssd1 vssd1 vccd1 vccd1 _01790_ sky130_fd_sc_hd__a22o_1
XANTENNA__07828__C1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10716_ net511 _05562_ _06315_ _06330_ vssd1 vssd1 vccd1 vccd1 _06331_ sky130_fd_sc_hd__a31o_1
X_13504_ _04497_ _02966_ vssd1 vssd1 vccd1 vccd1 _02972_ sky130_fd_sc_hd__nor2_1
XFILLER_9_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11696_ _06526_ net208 net422 net2912 vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__a22o_1
XFILLER_13_196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16223_ net2557 _02433_ net1220 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[1023\]
+ sky130_fd_sc_hd__dfrtp_1
X_10647_ _05666_ _05887_ _05900_ _05672_ _06202_ vssd1 vssd1 vccd1 vccd1 _06265_ sky130_fd_sc_hd__a221o_1
X_13435_ _03200_ _03248_ _02935_ vssd1 vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__o21a_1
X_14435__605 clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 net2074 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_77_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13366_ top.mmio.mem_data_i\[16\] net592 net1345 vssd1 vssd1 vccd1 vccd1 _02893_
+ sky130_fd_sc_hd__a21o_1
X_16154_ net2488 _02364_ net1251 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[954\]
+ sky130_fd_sc_hd__dfrtp_1
X_10578_ _06112_ _06198_ net390 vssd1 vssd1 vccd1 vccd1 _06199_ sky130_fd_sc_hd__mux2_1
X_15105_ net1487 _01318_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r2_prev\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_12317_ net2584 _03854_ net1183 vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__mux2_1
X_13297_ top.mmio.mem_data_i\[24\] top.mmio.mem_data_i\[26\] top.mmio.mem_data_i\[27\]
+ top.mmio.mem_data_i\[25\] vssd1 vssd1 vccd1 vccd1 _02840_ sky130_fd_sc_hd__or4bb_1
X_16085_ net2419 _02295_ net1211 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[885\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_138_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_110_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15036_ clknet_leaf_91_clk _01281_ net1270 vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__dfrtp_1
X_12248_ net433 top.CPU.registers.data\[22\] vssd1 vssd1 vccd1 vccd1 _06886_ sky130_fd_sc_hd__and2b_1
XFILLER_170_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11155__A2 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08556__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12179_ _06663_ net351 net170 net2679 vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__a22o_1
XFILLER_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10902__A2 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15407__RESET_B net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12104__A1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09505__C1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15938_ net2272 _02148_ net1173 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[738\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16549__CLK clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10666__A1 _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11863__B1 net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_125_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15869_ net2203 _02079_ net1121 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[669\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_88_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08410_ top.CPU.control_unit.instruction\[18\] _03160_ _03985_ vssd1 vssd1 vccd1
+ vccd1 _04049_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_125_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09390_ top.CPU.registers.data\[163\] top.CPU.registers.data\[131\] net828 vssd1
+ vssd1 vccd1 vccd1 _05029_ sky130_fd_sc_hd__mux2_1
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10928__B net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10418__A1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08341_ net678 _03962_ _03963_ vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__and3_1
XANTENNA__11615__A0 _06230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08087__A2 net1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08272_ net959 _03910_ _03907_ net615 vssd1 vssd1 vccd1 vccd1 _03911_ sky130_fd_sc_hd__a211o_1
XANTENNA__08492__C1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Left_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10944__A net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout127_A net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14178__348 clknet_leaf_140_clk vssd1 vssd1 vccd1 vccd1 net1817 sky130_fd_sc_hd__inv_2
XFILLER_164_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09587__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12040__B1 _06781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08244__C1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08414__A _04020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11394__A2 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08795__B1 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1036_A net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14219__389 clknet_leaf_163_clk vssd1 vssd1 vccd1 vccd1 net1858 sky130_fd_sc_hd__inv_2
XANTENNA__11146__A2 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout496_A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout124 _02936_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__buf_2
XFILLER_87_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout135 _05879_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__buf_2
Xfanout146 _06149_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__buf_2
XANTENNA_input1_A ACK_I vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout157 net159 vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__buf_6
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout168 net169 vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__buf_4
Xfanout179 _06795_ vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__clkbuf_4
X_07987_ top.CPU.registers.data\[664\] net1290 net1010 top.CPU.registers.data\[696\]
+ net907 vssd1 vssd1 vccd1 vccd1 _03626_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout663_A net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout284_X net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09726_ _05332_ _05363_ vssd1 vssd1 vccd1 vccd1 _05365_ sky130_fd_sc_hd__nor2_1
XFILLER_86_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09511__A2 net1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09657_ _04020_ _04051_ vssd1 vssd1 vccd1 vccd1 _05296_ sky130_fd_sc_hd__nor2_1
XANTENNA__08346__A_N net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11854__B1 net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout830_A net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout549_X net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout928_A net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08608_ top.CPU.registers.data\[655\] net1004 net929 _04246_ vssd1 vssd1 vccd1 vccd1
+ _04247_ sky130_fd_sc_hd__o211a_1
X_09588_ _05226_ vssd1 vssd1 vccd1 vccd1 _05227_ sky130_fd_sc_hd__inv_2
XFILLER_63_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11606__A0 _06033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08539_ top.CPU.registers.data\[592\] net1291 net1011 top.CPU.registers.data\[624\]
+ net935 vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__a221o_1
XANTENNA__09275__A1 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1360_X net1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14620__790 clknet_leaf_137_clk vssd1 vssd1 vccd1 vccd1 net2259 sky130_fd_sc_hd__inv_2
XANTENNA_fanout716_X net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11015__A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11550_ _06664_ net261 net248 net3113 vssd1 vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__a22o_1
XANTENNA__11082__B2 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07825__A2 net1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10501_ top.CPU.fetch.current_ra\[17\] net1044 net633 top.CPU.handler.toreg\[17\]
+ _06125_ vssd1 vssd1 vccd1 vccd1 _06126_ sky130_fd_sc_hd__a221o_2
X_11481_ _06611_ net261 net257 net3493 vssd1 vssd1 vccd1 vccd1 _02043_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_94_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13220_ top.I2C.output_state\[28\] _02791_ vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__nand2_1
XFILLER_7_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12031__A0 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10432_ _04052_ _05964_ net446 vssd1 vssd1 vccd1 vccd1 _06059_ sky130_fd_sc_hd__o21a_1
XANTENNA__08235__C1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11385__A2 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13151_ _07125_ _07126_ vssd1 vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__xnor2_1
X_10363_ _03923_ _05972_ vssd1 vssd1 vccd1 vccd1 _05993_ sky130_fd_sc_hd__or2_1
XFILLER_164_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08250__A2 _03887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12102_ top.CPU.registers.data\[101\] net645 vssd1 vssd1 vccd1 vccd1 _06819_ sky130_fd_sc_hd__or2_1
XFILLER_152_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13082_ top.CPU.data_out\[17\] net3257 net560 vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10294_ _05642_ _05926_ _05915_ vssd1 vssd1 vccd1 vccd1 _05927_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10860__Y _06467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11137__A2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12334__A1 _04855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08538__B1 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12033_ _06587_ _06779_ net150 net3078 vssd1 vssd1 vccd1 vccd1 _01553_ sky130_fd_sc_hd__a22o_1
XFILLER_105_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08002__A2 net1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11688__A3 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10896__A1 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_8_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout680 net684 vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__clkbuf_4
XFILLER_78_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07761__A1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout691 net701 vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__buf_4
XANTENNA__12098__B1 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10648__A1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15723_ net2057 _01933_ net1065 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[523\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09502__A2 net1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12935_ top.CPU.alu.program_counter\[29\] _03477_ vssd1 vssd1 vccd1 vccd1 _07376_
+ sky130_fd_sc_hd__or2_1
XANTENNA__11845__B1 net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11624__S net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15654_ net1988 _01864_ net1072 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[454\]
+ sky130_fd_sc_hd__dfrtp_1
X_12866_ top.CPU.alu.program_counter\[21\] _07298_ top.CPU.alu.program_counter\[22\]
+ vssd1 vssd1 vccd1 vccd1 _07314_ sky130_fd_sc_hd__a21oi_1
XFILLER_61_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11817_ net3429 _06213_ _06762_ vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15585_ net1919 _01795_ net1231 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[385\]
+ sky130_fd_sc_hd__dfrtp_1
X_12797_ top.CPU.alu.program_counter\[16\] _04189_ vssd1 vssd1 vccd1 vccd1 _07251_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_120_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11748_ _06230_ net536 net499 net192 net2788 vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__a32o_1
XANTENNA__10480__D_N _06105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11679_ _06496_ net199 net164 net3492 vssd1 vssd1 vccd1 vccd1 _01873_ sky130_fd_sc_hd__a22o_1
X_16206_ net2540 _02416_ net1107 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[1006\]
+ sky130_fd_sc_hd__dfrtp_1
X_13418_ top.I2C.data_out\[30\] net555 _02930_ vssd1 vssd1 vccd1 vccd1 _02931_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08226__C1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11376__A2 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16137_ net2471 _02347_ net1060 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[937\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_127_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13349_ net889 _02880_ vssd1 vssd1 vccd1 vccd1 _02881_ sky130_fd_sc_hd__and2_1
XANTENNA__08241__A2 net1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11298__C net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13916__86 clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 net1555 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_149_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16068_ net2402 _02278_ net1185 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[868\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_103_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12325__A1 _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13522__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11595__A net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15019_ clknet_leaf_96_clk _01264_ net1247 vssd1 vssd1 vccd1 vccd1 top.SPI.parameters\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_07910_ top.CPU.registers.data\[92\] net1302 net1023 top.CPU.registers.data\[124\]
+ net943 vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__a221o_1
X_08890_ net690 _04516_ _04519_ vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__or3_1
XFILLER_69_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10930__C net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07841_ top.CPU.registers.data\[189\] net1007 net905 vssd1 vssd1 vccd1 vccd1 _03480_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_127_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14563__733 clknet_leaf_114_clk vssd1 vssd1 vccd1 vccd1 net2202 sky130_fd_sc_hd__inv_2
XANTENNA__12089__B1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07772_ net920 _03410_ vssd1 vssd1 vccd1 vccd1 _03411_ sky130_fd_sc_hd__nand2_1
XANTENNA__10004__A net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09511_ top.CPU.registers.data\[449\] net1307 net1030 top.CPU.registers.data\[481\]
+ net923 vssd1 vssd1 vccd1 vccd1 _05150_ sky130_fd_sc_hd__a221o_1
XANTENNA__11836__B1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16447__RESET_B net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08701__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09442_ top.CPU.registers.data\[898\] net1294 net1015 top.CPU.registers.data\[930\]
+ net911 vssd1 vssd1 vccd1 vccd1 _05081_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_4_2_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14604__774 clknet_leaf_189_clk vssd1 vssd1 vccd1 vccd1 net2243 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_140_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09004__S net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09373_ top.CPU.registers.data_out_r2_prev\[3\] net687 _05010_ _05011_ net620 vssd1
+ vssd1 vccd1 vccd1 _05012_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout244_A _06748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_25_Left_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08324_ top.CPU.registers.data\[467\] net1301 net1017 top.CPU.registers.data\[499\]
+ net913 vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__a221o_1
XFILLER_21_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08465__C1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07807__A2 net1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08255_ top.CPU.registers.data\[854\] net1300 net1021 top.CPU.registers.data\[886\]
+ net941 vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout411_A net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10674__A net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout509_A net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1153_A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08186_ top.CPU.registers.data\[23\] net986 _03824_ vssd1 vssd1 vccd1 vccd1 _03825_
+ sky130_fd_sc_hd__a21o_1
XFILLER_146_661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11367__A2 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1320_A net1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09674__S net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout780_A net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11119__A2 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12316__A1 _03645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout878_A net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout499_X net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10327__B1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout666_X net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11827__A0 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09709_ net682 _05346_ _05347_ vssd1 vssd1 vccd1 vccd1 _05348_ sky130_fd_sc_hd__and3_1
X_10981_ _03167_ net501 net540 net141 vssd1 vssd1 vccd1 vccd1 _06543_ sky130_fd_sc_hd__or4b_1
XFILLER_74_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout833_X net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12095__A3 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13225__A _02780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12720_ _07175_ _07181_ net125 vssd1 vssd1 vccd1 vccd1 _07182_ sky130_fd_sc_hd__mux2_1
XFILLER_167_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12651_ top.CPU.done top.CPU.handler.state\[2\] _07055_ vssd1 vssd1 vccd1 vccd1 _00000_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09248__A1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11602_ _06482_ net428 net209 net214 net2804 vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__a32o_1
X_12582_ top.CPU.addressnew\[12\] top.CPU.addressnew\[17\] top.CPU.addressnew\[16\]
+ _06918_ vssd1 vssd1 vccd1 vccd1 _07086_ sky130_fd_sc_hd__or4_1
X_15370_ net1704 _01580_ net1091 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[170\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10263__C1 _05643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11533_ net483 _06231_ net354 net250 net2879 vssd1 vssd1 vccd1 vccd1 _01998_ sky130_fd_sc_hd__a32o_1
XANTENNA__11032__X _06575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11464_ _06311_ net3364 net263 vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__mux2_1
XFILLER_171_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11358__A2 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10415_ _03242_ net396 net403 vssd1 vssd1 vccd1 vccd1 _06043_ sky130_fd_sc_hd__a21oi_1
X_13203_ net3784 _02779_ _02781_ _02773_ vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__a22o_1
XFILLER_87_1032 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11395_ _06521_ net282 net274 net3380 vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__a22o_1
XFILLER_125_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09584__S net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10346_ _05859_ _05976_ net390 vssd1 vssd1 vccd1 vccd1 _05977_ sky130_fd_sc_hd__mux2_1
X_13134_ top.SPI.counter\[1\] net594 _02728_ vssd1 vssd1 vccd1 vccd1 _02736_ sky130_fd_sc_hd__a21o_1
XFILLER_48_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07982__A1 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11619__S net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09708__C1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13065_ top.CPU.data_out\[0\] net2718 net560 vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__mux2_1
X_10277_ _03649_ _05300_ _05367_ net371 _05909_ vssd1 vssd1 vccd1 vccd1 _05910_ sky130_fd_sc_hd__a311o_1
X_14250__420 clknet_leaf_145_clk vssd1 vssd1 vccd1 vccd1 net1889 sky130_fd_sc_hd__inv_2
X_12016_ top.CPU.registers.data\[153\] net656 _06581_ net364 net568 vssd1 vssd1 vccd1
+ vccd1 _06785_ sky130_fd_sc_hd__o2111a_1
X_14547__717 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 net2186 sky130_fd_sc_hd__inv_2
XANTENNA__10869__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08931__B1 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11530__A2 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13807__B2 top.CPU.data_out\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10759__A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10097__A2 _05670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15706_ net2040 _01916_ net1252 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[506\]
+ sky130_fd_sc_hd__dfrtp_1
X_12918_ top.CPU.alu.program_counter\[27\] _07346_ vssd1 vssd1 vccd1 vccd1 _07361_
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_122_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08695__C1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11294__B2 _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11833__A3 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15637_ net1971 _01847_ net1217 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[437\]
+ sky130_fd_sc_hd__dfrtp_1
X_12849_ top.CPU.alu.program_counter\[20\] _07287_ vssd1 vssd1 vccd1 vccd1 _07299_
+ sky130_fd_sc_hd__nor2_1
XFILLER_21_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08447__C1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08663__S net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15568_ net1902 _01778_ net1107 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[368\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12693__B _04856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08998__B1 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15499_ net1833 _01709_ net1064 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[299\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08462__A2 net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08040_ _03675_ _03678_ net1308 vssd1 vssd1 vccd1 vccd1 _03679_ sky130_fd_sc_hd__o21ai_1
XFILLER_174_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11349__A2 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11102__B net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold903 top.CPU.registers.data\[776\] vssd1 vssd1 vccd1 vccd1 net3460 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold914 top.CPU.registers.data\[1016\] vssd1 vssd1 vccd1 vccd1 net3471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold925 top.CPU.registers.data\[308\] vssd1 vssd1 vccd1 vccd1 net3482 sky130_fd_sc_hd__dlygate4sd3_1
Xhold936 top.CPU.registers.data\[633\] vssd1 vssd1 vccd1 vccd1 net3493 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold947 top.CPU.registers.data\[695\] vssd1 vssd1 vccd1 vccd1 net3504 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09347__X _04986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold958 top.CPU.registers.data\[917\] vssd1 vssd1 vccd1 vccd1 net3515 sky130_fd_sc_hd__dlygate4sd3_1
X_09991_ _05628_ _05629_ vssd1 vssd1 vccd1 vccd1 _05630_ sky130_fd_sc_hd__nor2_1
XFILLER_115_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold969 top.CPU.registers.data\[734\] vssd1 vssd1 vccd1 vccd1 net3526 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10309__A0 _03613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08942_ top.CPU.registers.data\[682\] net1374 net971 top.CPU.registers.data\[650\]
+ net902 vssd1 vssd1 vccd1 vccd1 _04581_ sky130_fd_sc_hd__a221o_1
X_08873_ top.CPU.registers.data\[75\] net1311 net842 top.CPU.registers.data\[107\]
+ net762 vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__a221o_1
XFILLER_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07725__A1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout194_A net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07824_ top.CPU.registers.data\[189\] top.CPU.registers.data\[157\] net816 vssd1
+ vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__mux2_1
X_13838__8 clknet_leaf_121_clk vssd1 vssd1 vccd1 vccd1 net1477 sky130_fd_sc_hd__inv_2
XANTENNA__09478__A1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07755_ top.CPU.registers.data\[446\] top.CPU.registers.data\[414\] net834 vssd1
+ vssd1 vccd1 vccd1 _03394_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout361_A net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout459_A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07686_ _03285_ net632 _03306_ vssd1 vssd1 vccd1 vccd1 _03325_ sky130_fd_sc_hd__and3_1
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09425_ top.CPU.registers.data\[34\] top.CPU.registers.data\[2\] net986 vssd1 vssd1
+ vccd1 vccd1 _05064_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1270_A net1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout247_X net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout626_A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12234__B1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09356_ top.CPU.registers.data\[899\] net1297 net1018 top.CPU.registers.data\[931\]
+ net915 vssd1 vssd1 vccd1 vccd1 _04995_ sky130_fd_sc_hd__a221o_1
XFILLER_40_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08307_ net707 _03944_ _03945_ _03943_ vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_43_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09287_ top.CPU.registers.data\[836\] net1299 net1020 top.CPU.registers.data\[868\]
+ net940 vssd1 vssd1 vccd1 vccd1 _04926_ sky130_fd_sc_hd__a221o_1
XFILLER_20_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14691__861 clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 net2330 sky130_fd_sc_hd__inv_2
XFILLER_138_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08238_ top.CPU.registers.data\[566\] top.CPU.registers.data\[534\] net835 vssd1
+ vssd1 vccd1 vccd1 _03877_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout995_A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11012__B net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08169_ top.CPU.registers.data\[983\] net1325 net856 top.CPU.registers.data\[1015\]
+ net723 vssd1 vssd1 vccd1 vccd1 _03808_ sky130_fd_sc_hd__a221o_1
XFILLER_134_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1323_X net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10200_ _05833_ _05834_ _05835_ net395 _05754_ vssd1 vssd1 vccd1 vccd1 _05836_ sky130_fd_sc_hd__a221o_1
XFILLER_162_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14234__404 clknet_leaf_161_clk vssd1 vssd1 vccd1 vccd1 net1873 sky130_fd_sc_hd__inv_2
X_11180_ net490 _06488_ _06643_ net300 net2872 vssd1 vssd1 vccd1 vccd1 _02264_ sky130_fd_sc_hd__a32o_1
XANTENNA__08610__C1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10131_ top.CPU.handler.toreg\[30\] net881 vssd1 vssd1 vccd1 vccd1 _05769_ sky130_fd_sc_hd__and2_1
XANTENNA__11760__A2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09166__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10062_ _05123_ net377 vssd1 vssd1 vccd1 vccd1 _05700_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_89_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09705__A2 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout950_X net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16369__RESET_B net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12170__C1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13654__S net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11512__A2 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13821_ net3091 net334 net327 top.CPU.data_out\[23\] vssd1 vssd1 vccd1 vccd1 _02701_
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10579__A net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16540_ clknet_leaf_85_clk net3497 net1265 vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__dfrtp_1
XFILLER_62_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13752_ _03086_ _03087_ vssd1 vssd1 vccd1 vccd1 _02641_ sky130_fd_sc_hd__and2_1
XANTENNA__11276__B2 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10964_ net3890 net218 _06533_ net320 vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__a22o_1
X_12703_ _07164_ _07165_ vssd1 vssd1 vccd1 vccd1 _07166_ sky130_fd_sc_hd__nor2_1
X_16471_ clknet_leaf_88_clk _02633_ net1272 vssd1 vssd1 vccd1 vccd1 top.SPI.timem\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13683_ net2655 net332 vssd1 vssd1 vccd1 vccd1 _02611_ sky130_fd_sc_hd__and2_1
XFILLER_71_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10895_ net659 _06056_ net436 vssd1 vssd1 vccd1 vccd1 _06491_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_100_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09579__S net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15422_ net1756 _01632_ net1238 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[222\]
+ sky130_fd_sc_hd__dfrtp_1
X_12634_ top.I2C.output_state\[26\] net2782 vssd1 vssd1 vccd1 vccd1 _00013_ sky130_fd_sc_hd__and2_1
XANTENNA__08429__C1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12225__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15933__RESET_B net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15353_ net1687 _01563_ net1239 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[153\]
+ sky130_fd_sc_hd__dfrtp_1
X_12565_ _06371_ _06389_ _07069_ vssd1 vssd1 vccd1 vccd1 _07070_ sky130_fd_sc_hd__and3_1
XFILLER_12_773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08444__A2 net1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11516_ _06647_ net262 net253 net3461 vssd1 vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_22_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15284_ net1618 _01494_ net1074 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[84\]
+ sky130_fd_sc_hd__dfrtp_1
X_12496_ _05154_ _05190_ vssd1 vssd1 vccd1 vccd1 _07005_ sky130_fd_sc_hd__nand2_1
XFILLER_138_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12018__B _06781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11447_ net3337 net265 _06723_ net490 vssd1 vssd1 vccd1 vccd1 _02071_ sky130_fd_sc_hd__a22o_1
XFILLER_171_247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11200__A1 net1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11378_ _06493_ net277 net272 net3352 vssd1 vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__a22o_1
XFILLER_98_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10761__B _06373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07955__A1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11751__A2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13117_ net2672 _02723_ net897 vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__mux2_1
X_10329_ _03167_ _05960_ vssd1 vssd1 vccd1 vccd1 _05961_ sky130_fd_sc_hd__nor2_1
XANTENNA__10480__C net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13048_ net2994 _07449_ net895 vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__mux2_1
XFILLER_61_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14018__188 clknet_leaf_147_clk vssd1 vssd1 vccd1 vccd1 net1657 sky130_fd_sc_hd__inv_2
XFILLER_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12700__A1 top.CPU.alu.program_counter\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1250 net1259 vssd1 vssd1 vccd1 vccd1 net1250 sky130_fd_sc_hd__clkbuf_4
Xfanout1261 net1262 vssd1 vssd1 vccd1 vccd1 net1261 sky130_fd_sc_hd__clkbuf_4
Xfanout1272 net1275 vssd1 vssd1 vccd1 vccd1 net1272 sky130_fd_sc_hd__clkbuf_2
Xfanout1283 net1285 vssd1 vssd1 vccd1 vccd1 net1283 sky130_fd_sc_hd__buf_4
Xfanout1294 net1301 vssd1 vssd1 vccd1 vccd1 net1294 sky130_fd_sc_hd__clkbuf_4
XFILLER_38_158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11592__B net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14999_ clknet_leaf_93_clk _01244_ net1262 vssd1 vssd1 vccd1 vccd1 top.SPI.parameters\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_80_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07540_ _03160_ _03163_ net1038 _03118_ vssd1 vssd1 vccd1 vccd1 _03179_ sky130_fd_sc_hd__a31oi_1
X_07471_ top.CPU.control_unit.instruction\[17\] vssd1 vssd1 vccd1 vccd1 _03111_ sky130_fd_sc_hd__inv_2
XANTENNA__13008__A2 _07429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11812__S _06762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09489__S net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09210_ top.CPU.registers.data\[70\] net1287 net1006 top.CPU.registers.data\[102\]
+ net930 vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__a221o_1
XANTENNA__11019__B2 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14675__845 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 net2314 sky130_fd_sc_hd__inv_2
XANTENNA__10936__B net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_95_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09141_ top.CPU.registers.data\[391\] net1304 net1024 top.CPU.registers.data\[423\]
+ net919 vssd1 vssd1 vccd1 vccd1 _04780_ sky130_fd_sc_hd__a221o_1
XANTENNA__15674__RESET_B net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10778__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10242__A2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09072_ net951 _04707_ _04710_ net624 vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_135_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14716__886 clknet_leaf_139_clk vssd1 vssd1 vccd1 vccd1 net2355 sky130_fd_sc_hd__inv_2
XFILLER_30_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08023_ net705 _03660_ _03661_ vssd1 vssd1 vccd1 vccd1 _03662_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_135_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11990__A2 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold700 top.SPI.parameters\[17\] vssd1 vssd1 vccd1 vccd1 net3257 sky130_fd_sc_hd__dlygate4sd3_1
Xhold711 top.CPU.registers.data\[397\] vssd1 vssd1 vccd1 vccd1 net3268 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout207_A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold722 top.CPU.registers.data\[460\] vssd1 vssd1 vccd1 vccd1 net3279 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold733 top.CPU.registers.data\[894\] vssd1 vssd1 vccd1 vccd1 net3290 sky130_fd_sc_hd__dlygate4sd3_1
Xhold744 top.CPU.registers.data\[525\] vssd1 vssd1 vccd1 vccd1 net3301 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold755 top.CPU.registers.data\[614\] vssd1 vssd1 vccd1 vccd1 net3312 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_153_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold766 top.CPU.registers.data\[490\] vssd1 vssd1 vccd1 vccd1 net3323 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold777 top.CPU.registers.data\[489\] vssd1 vssd1 vccd1 vccd1 net3334 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11742__A2 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold788 top.CPU.registers.data\[288\] vssd1 vssd1 vccd1 vccd1 net3345 sky130_fd_sc_hd__dlygate4sd3_1
X_09974_ _05602_ _05603_ _03580_ _05512_ vssd1 vssd1 vccd1 vccd1 _05613_ sky130_fd_sc_hd__a211o_1
XFILLER_130_111 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold799 top.CPU.registers.data\[203\] vssd1 vssd1 vccd1 vccd1 net3356 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09148__B1 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_33_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08925_ net787 _04562_ _04563_ net741 vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__o211a_1
XANTENNA__13474__S net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13495__A2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout576_A _03169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout197_X net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1400 top.CPU.registers.data\[89\] vssd1 vssd1 vccd1 vccd1 net3957 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1411 top.mmio.mem_data_i\[4\] vssd1 vssd1 vccd1 vccd1 net3968 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1422 top.CPU.registers.data\[66\] vssd1 vssd1 vccd1 vccd1 net3979 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1433 top.SPI.timem\[9\] vssd1 vssd1 vccd1 vccd1 net3990 sky130_fd_sc_hd__dlygate4sd3_1
X_08856_ net1366 _04491_ _04494_ vssd1 vssd1 vccd1 vccd1 _04495_ sky130_fd_sc_hd__o21a_1
X_13900__70 clknet_leaf_193_clk vssd1 vssd1 vccd1 vccd1 net1539 sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_168_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1444 top.CPU.registers.data\[122\] vssd1 vssd1 vccd1 vccd1 net4001 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1455 top.SPI.register\[0\] vssd1 vssd1 vccd1 vccd1 net4012 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09253__A _04891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1466 top.I2C.I2C_state\[2\] vssd1 vssd1 vccd1 vccd1 net4023 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_55_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07807_ top.CPU.registers.data\[669\] net1319 net850 top.CPU.registers.data\[701\]
+ net704 vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__a221o_1
XFILLER_84_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout364_X net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08787_ _04422_ _04425_ net635 vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout743_A net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_48_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07738_ top.CPU.registers.data\[958\] top.CPU.registers.data\[926\] top.CPU.registers.data\[830\]
+ top.CPU.registers.data\[798\] net833 net730 vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__mux4_1
XANTENNA__08659__C1 net1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08123__A1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout531_X net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout910_A _03353_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07669_ net632 _03298_ _03305_ vssd1 vssd1 vccd1 vccd1 _03308_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout629_X net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_9_Left_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09408_ top.CPU.registers.data\[643\] net1328 net859 top.CPU.registers.data\[675\]
+ net727 vssd1 vssd1 vccd1 vccd1 _05047_ sky130_fd_sc_hd__a221o_1
X_10680_ _06218_ _06295_ net388 vssd1 vssd1 vccd1 vccd1 _06296_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12207__B1 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09339_ net696 _04975_ _04976_ _04977_ vssd1 vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_109_Right_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09623__A1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_106_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11023__A net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12350_ net898 net2969 vssd1 vssd1 vccd1 vccd1 _00065_ sky130_fd_sc_hd__nor2_1
XFILLER_127_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout998_X net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13649__S net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11301_ net3463 net291 net359 net133 vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__a22o_1
XANTENNA__11981__A2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12281_ net2601 _05331_ net1240 vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__mux2_1
XFILLER_4_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10862__A net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09387__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11232_ net571 net528 net134 net546 vssd1 vssd1 vccd1 vccd1 _06671_ sky130_fd_sc_hd__and4_1
XFILLER_106_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11733__A2 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10073__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11163_ net513 _06466_ vssd1 vssd1 vccd1 vccd1 _06642_ sky130_fd_sc_hd__nor2_1
XFILLER_84_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09139__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10114_ net409 _05616_ vssd1 vssd1 vccd1 vccd1 _05752_ sky130_fd_sc_hd__or2_2
XFILLER_136_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15971_ net2305 _02181_ net1208 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[771\]
+ sky130_fd_sc_hd__dfrtp_1
X_11094_ net574 net530 net138 vssd1 vssd1 vccd1 vccd1 _06605_ sky130_fd_sc_hd__and3_1
XFILLER_49_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10045_ _03306_ _03310_ _03322_ _03319_ vssd1 vssd1 vccd1 vccd1 _05684_ sky130_fd_sc_hd__a31oi_2
X_14922_ clknet_leaf_30_clk _01168_ net1152 vssd1 vssd1 vccd1 vccd1 top.CPU.alu.program_counter\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__11497__A1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_10_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold60 top.CPU.handler.state\[4\] vssd1 vssd1 vccd1 vccd1 net2617 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 _00036_ vssd1 vssd1 vccd1 vccd1 net2628 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 net41 vssd1 vssd1 vccd1 vccd1 net2639 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold93 top.CPU.registers.data\[806\] vssd1 vssd1 vccd1 vccd1 net2650 sky130_fd_sc_hd__dlygate4sd3_1
X_13804_ net3155 net334 net327 top.CPU.data_out\[6\] vssd1 vssd1 vccd1 vccd1 _02684_
+ sky130_fd_sc_hd__a22o_1
XFILLER_17_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10102__A net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14362__532 clknet_leaf_162_clk vssd1 vssd1 vccd1 vccd1 net2001 sky130_fd_sc_hd__inv_2
XANTENNA__08114__A1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11996_ _06563_ net344 net181 net2840 vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__a22o_1
XFILLER_17_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16523_ clknet_leaf_100_clk _02685_ net1255 vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__dfrtp_1
X_14659__829 clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 net2298 sky130_fd_sc_hd__inv_2
X_13735_ top.SPI.timem\[15\] top.SPI.timem\[16\] _03074_ vssd1 vssd1 vccd1 vccd1 _03077_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10459__D net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10947_ net3529 net222 _06522_ net312 vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_27_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16454_ clknet_leaf_81_clk _02617_ net1242 vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__dfrtp_1
XFILLER_71_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13666_ _06919_ net890 _03045_ _07089_ vssd1 vssd1 vccd1 vccd1 _03048_ sky130_fd_sc_hd__o211a_1
X_10878_ _05693_ _06479_ vssd1 vssd1 vccd1 vccd1 _06480_ sky130_fd_sc_hd__and2_1
X_14403__573 clknet_leaf_171_clk vssd1 vssd1 vccd1 vccd1 net2042 sky130_fd_sc_hd__inv_2
X_15405_ net1739 _01615_ net1059 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[205\]
+ sky130_fd_sc_hd__dfrtp_1
X_12617_ _07095_ _07096_ _07103_ _07115_ top.SPI.state\[4\] vssd1 vssd1 vccd1 vccd1
+ _00072_ sky130_fd_sc_hd__a32o_1
X_16385_ clknet_leaf_65_clk _02594_ net1163 vssd1 vssd1 vccd1 vccd1 top.CPU.handler.writeout
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09075__C1 net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13597_ top.CPU.alu.program_counter\[19\] net1349 vssd1 vssd1 vccd1 vccd1 _03025_
+ sky130_fd_sc_hd__nor2_1
Xclkbuf_4_14_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_14_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__15085__RESET_B net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15336_ net1670 _01546_ net1089 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[136\]
+ sky130_fd_sc_hd__dfrtp_1
X_12548_ _07053_ _07056_ vssd1 vssd1 vccd1 vccd1 _07057_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_117_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11972__A2 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15267_ net1601 _01477_ net1210 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[67\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_172_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10772__A _05754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_2 _06645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ _06983_ _06984_ _06985_ _06986_ _06987_ vssd1 vssd1 vccd1 vccd1 _06988_ sky130_fd_sc_hd__a311o_1
XFILLER_6_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15198_ clknet_leaf_90_clk _01408_ net1271 vssd1 vssd1 vccd1 vccd1 top.SPI.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_113_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11185__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11724__A2 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout509 net510 vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_130_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09772__S net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_807 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13477__A2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08710_ top.CPU.registers.data\[429\] top.CPU.registers.data\[397\] net807 vssd1
+ vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__mux2_1
X_13970__140 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 net1609 sky130_fd_sc_hd__inv_2
XANTENNA__08889__C1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09690_ net803 _05322_ _05328_ vssd1 vssd1 vccd1 vccd1 _05329_ sky130_fd_sc_hd__and3_1
XFILLER_6_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1080 net1082 vssd1 vssd1 vccd1 vccd1 net1080 sky130_fd_sc_hd__clkbuf_4
Xfanout1091 net1093 vssd1 vssd1 vccd1 vccd1 net1091 sky130_fd_sc_hd__clkbuf_2
XFILLER_55_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08641_ top.CPU.registers.data\[206\] net818 net769 _04263_ vssd1 vssd1 vccd1 vccd1
+ _04280_ sky130_fd_sc_hd__a211o_1
XFILLER_66_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11108__A net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08572_ top.CPU.registers.data\[815\] top.CPU.registers.data\[783\] net811 vssd1
+ vssd1 vccd1 vccd1 _04211_ sky130_fd_sc_hd__mux2_1
XFILLER_23_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07523_ _03144_ _03157_ vssd1 vssd1 vccd1 vccd1 _03162_ sky130_fd_sc_hd__nand2_2
XANTENNA__08656__A2 _04291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout157_A net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09520__B net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09605__A1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout324_A net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09124_ top.CPU.registers.data_out_r1_prev\[7\] net875 _04748_ _04762_ vssd1 vssd1
+ vccd1 vccd1 _04763_ sky130_fd_sc_hd__o211ai_4
XFILLER_108_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09055_ net738 _04684_ _04685_ net690 vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__a31o_1
XANTENNA__11963__A2 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1233_A net1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08006_ _03629_ _03644_ vssd1 vssd1 vccd1 vccd1 _03645_ sky130_fd_sc_hd__or2_4
XFILLER_163_578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold530 top.CPU.registers.data\[306\] vssd1 vssd1 vccd1 vccd1 net3087 sky130_fd_sc_hd__dlygate4sd3_1
X_14839__1009 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 net2478 sky130_fd_sc_hd__inv_2
XFILLER_151_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold541 top.CPU.registers.data\[990\] vssd1 vssd1 vccd1 vccd1 net3098 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout693_A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold552 top.CPU.registers.data\[419\] vssd1 vssd1 vccd1 vccd1 net3109 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07919__A1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11715__A2 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold563 top.CPU.registers.data\[788\] vssd1 vssd1 vccd1 vccd1 net3120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 top.CPU.registers.data\[972\] vssd1 vssd1 vccd1 vccd1 net3131 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08041__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold585 net75 vssd1 vssd1 vccd1 vccd1 net3142 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold596 top.CPU.registers.data\[542\] vssd1 vssd1 vccd1 vccd1 net3153 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09957_ _03650_ _05594_ _05529_ vssd1 vssd1 vccd1 vccd1 _05596_ sky130_fd_sc_hd__a21o_1
XFILLER_132_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout481_X net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout860_A net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13877__47 clknet_leaf_171_clk vssd1 vssd1 vccd1 vccd1 net1516 sky130_fd_sc_hd__inv_2
XFILLER_131_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout958_A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout579_X net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08908_ top.CPU.registers.data\[42\] top.CPU.registers.data\[10\] net809 vssd1 vssd1
+ vccd1 vccd1 _04547_ sky130_fd_sc_hd__mux2_1
X_09888_ _03374_ _03445_ _03581_ _05513_ vssd1 vssd1 vccd1 vccd1 _05527_ sky130_fd_sc_hd__and4_1
XANTENNA__08344__A1 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1230 top.CPU.registers.data\[236\] vssd1 vssd1 vccd1 vccd1 net3787 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1241 top.CPU.handler.toreg\[10\] vssd1 vssd1 vccd1 vccd1 net3798 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09541__B1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1252 top.CPU.registers.data\[237\] vssd1 vssd1 vccd1 vccd1 net3809 sky130_fd_sc_hd__dlygate4sd3_1
X_08839_ top.CPU.registers.data\[939\] top.CPU.registers.data\[907\] net964 vssd1
+ vssd1 vccd1 vccd1 _04478_ sky130_fd_sc_hd__mux2_1
X_14346__516 clknet_leaf_145_clk vssd1 vssd1 vccd1 vccd1 net1985 sky130_fd_sc_hd__inv_2
XANTENNA_fanout1390_X net1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1263 top.CPU.registers.data\[742\] vssd1 vssd1 vccd1 vccd1 net3820 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1274 top.CPU.fetch.current_ra\[11\] vssd1 vssd1 vccd1 vccd1 net3831 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout746_X net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1285 top.CPU.registers.data\[35\] vssd1 vssd1 vccd1 vccd1 net3842 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11018__A net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1296 top.CPU.registers.data\[1012\] vssd1 vssd1 vccd1 vccd1 net3853 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12428__B1 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11850_ _06682_ net196 net152 net2917 vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__a22o_1
XFILLER_167_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10801_ net601 _06410_ _06411_ vssd1 vssd1 vccd1 vccd1 _06412_ sky130_fd_sc_hd__a21o_2
XFILLER_122_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13504__Y _02972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10857__A net1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11781_ _06626_ net234 net160 net3309 vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout913_X net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08647__A2 net1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11452__S net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13520_ top.CPU.data_out\[18\] net589 net339 _02980_ vssd1 vssd1 vccd1 vccd1 _02516_
+ sky130_fd_sc_hd__o22a_1
X_10732_ net409 _06344_ _06345_ vssd1 vssd1 vccd1 vccd1 _06346_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_24_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13451_ _02892_ _02937_ _02939_ vssd1 vssd1 vccd1 vccd1 _02947_ sky130_fd_sc_hd__a21o_1
X_10663_ net397 _06198_ vssd1 vssd1 vccd1 vccd1 _06280_ sky130_fd_sc_hd__nand2_1
X_12402_ _03120_ top.I2C.I2C_state\[8\] net2613 vssd1 vssd1 vccd1 vccd1 _00038_ sky130_fd_sc_hd__a21o_1
X_16170_ net2504 _02380_ net1084 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[970\]
+ sky130_fd_sc_hd__dfrtp_1
X_13382_ net888 _02904_ vssd1 vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__and2_1
X_10594_ net3858 net225 net311 _06214_ vssd1 vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_97_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15121_ clknet_leaf_51_clk net3937 net1132 vssd1 vssd1 vccd1 vccd1 top.I2C.scl_out
+ sky130_fd_sc_hd__dfstp_1
XFILLER_139_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11954__A2 _06500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12333_ net2572 _04792_ net1199 vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__mux2_1
XANTENNA__10592__A net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09158__A _04765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15052_ clknet_leaf_73_clk _01297_ net1158 vssd1 vssd1 vccd1 vccd1 top.CPU.alu.program_counter\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_12264_ net2880 _06334_ net433 vssd1 vssd1 vccd1 vccd1 _01417_ sky130_fd_sc_hd__mux2_1
XANTENNA__11167__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11706__A2 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11215_ net1403 net472 net540 _06603_ vssd1 vssd1 vccd1 vccd1 _06662_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_75_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12195_ net475 _06672_ _06864_ net171 net3553 vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__a32o_1
Xoutput50 net50 vssd1 vssd1 vccd1 vccd1 ADR_O[1] sky130_fd_sc_hd__buf_2
Xoutput61 net61 vssd1 vssd1 vccd1 vccd1 ADR_O[4] sky130_fd_sc_hd__buf_2
XANTENNA__10914__B1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 DAT_O[13] sky130_fd_sc_hd__buf_2
XANTENNA__09445__X _05084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput83 net83 vssd1 vssd1 vccd1 vccd1 DAT_O[23] sky130_fd_sc_hd__buf_2
X_13954__124 clknet_leaf_140_clk vssd1 vssd1 vccd1 vccd1 net1593 sky130_fd_sc_hd__inv_2
X_11146_ net487 net464 _06632_ net303 net3299 vssd1 vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__a32o_1
XFILLER_96_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10390__A1 _05733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput94 net94 vssd1 vssd1 vccd1 vccd1 DAT_O[4] sky130_fd_sc_hd__buf_2
XANTENNA__13459__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11627__S net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07791__C1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13408__A net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11077_ net438 _06373_ net534 vssd1 vssd1 vccd1 vccd1 _06594_ sky130_fd_sc_hd__and3_1
X_15954_ net2288 _02164_ net1081 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[754\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12131__A2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10028_ net404 _05665_ vssd1 vssd1 vccd1 vccd1 _05667_ sky130_fd_sc_hd__nand2_2
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09532__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_196_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_196_clk
+ sky130_fd_sc_hd__clkbuf_8
X_15885_ net2219 _02095_ net1077 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[685\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_64_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08886__A2 net1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14089__259 clknet_leaf_155_clk vssd1 vssd1 vccd1 vccd1 net1728 sky130_fd_sc_hd__inv_2
XANTENNA__08936__S net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13891__61 clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 net1530 sky130_fd_sc_hd__inv_2
XFILLER_64_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09296__C1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11979_ _06536_ net347 net182 net3569 vssd1 vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__a22o_1
XANTENNA__08638__A2 net1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09835__A1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16506_ clknet_leaf_49_clk _02668_ net1128 vssd1 vssd1 vccd1 vccd1 top.mmio.mem_data_i\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11215__X _06662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13718_ top.SPI.timem\[9\] top.SPI.timem\[10\] _03062_ vssd1 vssd1 vccd1 vccd1 _03066_
+ sky130_fd_sc_hd__and3_1
XFILLER_16_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16437_ clknet_leaf_80_clk _02600_ net1241 vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__dfrtp_1
X_13649_ net3259 _07305_ net663 vssd1 vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__mux2_1
XANTENNA__09048__C1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16368_ clknet_leaf_62_clk _02577_ net1164 vssd1 vssd1 vccd1 vccd1 top.CPU.fetch.current_ra\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_157_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09063__A2 net1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15319_ net1653 _01529_ net1183 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[119\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_132_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16299_ clknet_leaf_108_clk _02508_ net1246 vssd1 vssd1 vccd1 vccd1 top.CPU.data_out\[10\]
+ sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_120_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_120_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13147__A1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14490__660 clknet_leaf_162_clk vssd1 vssd1 vccd1 vccd1 net2129 sky130_fd_sc_hd__inv_2
XFILLER_145_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14787__957 clknet_leaf_170_clk vssd1 vssd1 vccd1 vccd1 net2426 sky130_fd_sc_hd__inv_2
XFILLER_67_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11110__B net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12921__S net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout306 net307 vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08574__A1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09811_ net758 _05444_ _05445_ _05449_ vssd1 vssd1 vccd1 vccd1 _05450_ sky130_fd_sc_hd__a31o_1
XANTENNA__09771__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout317 net322 vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__clkbuf_4
Xfanout328 net329 vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__clkbuf_2
Xfanout339 _02978_ vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__buf_2
X_14033__203 clknet_leaf_187_clk vssd1 vssd1 vccd1 vccd1 net1672 sky130_fd_sc_hd__inv_2
XANTENNA_clkload11_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14828__998 clknet_leaf_195_clk vssd1 vssd1 vccd1 vccd1 net2467 sky130_fd_sc_hd__inv_2
XANTENNA__10441__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13318__A _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09742_ top.CPU.registers.data\[475\] net1331 net862 top.CPU.registers.data\[507\]
+ net775 vssd1 vssd1 vccd1 vccd1 _05381_ sky130_fd_sc_hd__a221o_1
XANTENNA__12122__A2 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09523__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10669__C1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09673_ top.CPU.registers.data\[313\] top.CPU.registers.data\[281\] net837 vssd1
+ vssd1 vccd1 vccd1 _05312_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_187_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_187_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout274_A _06714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11330__B1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08624_ top.CPU.registers.data\[238\] net1387 vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__and2_1
XANTENNA__08846__S net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10948__Y _06523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07603__X _03242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08555_ _04193_ vssd1 vssd1 vccd1 vccd1 _04194_ sky130_fd_sc_hd__inv_2
XANTENNA__09826__A1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09287__C1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout441_A net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1183_A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07837__A0 top.CPU.alu.program_counter\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07506_ top.CPU.control_unit.instruction\[3\] top.CPU.control_unit.instruction\[2\]
+ top.CPU.control_unit.instruction\[0\] top.CPU.control_unit.instruction\[1\] vssd1
+ vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__and4bb_1
X_08486_ _04093_ _04124_ vssd1 vssd1 vccd1 vccd1 _04125_ sky130_fd_sc_hd__nor2_1
XANTENNA__08147__A _03755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09039__C1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12892__A top.CPU.alu.program_counter\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout706_A _03212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07986__A net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_99_Left_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14731__901 clknet_leaf_149_clk vssd1 vssd1 vccd1 vccd1 net2370 sky130_fd_sc_hd__inv_2
X_09107_ net800 _04740_ _04741_ net754 vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__o211a_1
XANTENNA__11936__A2 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13500__B _02967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_111_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_111_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13138__A1 top.CPU.data_out\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1236_X net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09038_ net788 _04674_ _04675_ _04676_ net691 vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__a311o_1
XFILLER_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout696_X net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13938__108 clknet_leaf_193_clk vssd1 vssd1 vccd1 vccd1 net1577 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_92_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11020__B _03170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12831__S net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold360 top.CPU.registers.data\[301\] vssd1 vssd1 vccd1 vccd1 net2917 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09211__C1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold371 top.CPU.registers.data\[803\] vssd1 vssd1 vccd1 vccd1 net2928 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1403_X net1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold382 top.CPU.registers.data\[986\] vssd1 vssd1 vccd1 vccd1 net2939 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08565__A1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold393 top.CPU.registers.data\[441\] vssd1 vssd1 vccd1 vccd1 net2950 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ net3046 net216 _06554_ net311 vssd1 vssd1 vccd1 vccd1 _02349_ sky130_fd_sc_hd__a22o_1
XFILLER_78_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09762__B1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10372__A1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout863_X net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout840 net854 vssd1 vssd1 vccd1 vccd1 net840 sky130_fd_sc_hd__clkbuf_4
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout851 net853 vssd1 vssd1 vccd1 vccd1 net851 sky130_fd_sc_hd__clkbuf_4
XFILLER_131_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout862 _03203_ vssd1 vssd1 vccd1 vccd1 net862 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout873 net874 vssd1 vssd1 vccd1 vccd1 net873 sky130_fd_sc_hd__clkbuf_4
Xfanout884 _03095_ vssd1 vssd1 vccd1 vccd1 net884 sky130_fd_sc_hd__buf_2
XANTENNA__12113__A2 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09514__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout895 net896 vssd1 vssd1 vccd1 vccd1 net895 sky130_fd_sc_hd__clkbuf_4
XANTENNA__15777__RESET_B net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12951_ _07388_ _07390_ vssd1 vssd1 vccd1 vccd1 _07391_ sky130_fd_sc_hd__nor2_1
XFILLER_46_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_178_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_178_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold1060 top.SPI.paroutput\[29\] vssd1 vssd1 vccd1 vccd1 net3617 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_19_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11321__B1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1071 top.CPU.registers.data\[634\] vssd1 vssd1 vccd1 vccd1 net3628 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_133_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11902_ net3505 net186 net350 _05772_ vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__a22o_1
XANTENNA__15706__RESET_B net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15670_ net2004 _01880_ net1227 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[470\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1082 top.CPU.registers.data\[252\] vssd1 vssd1 vccd1 vccd1 net3639 sky130_fd_sc_hd__dlygate4sd3_1
X_12882_ _07326_ _07327_ vssd1 vssd1 vccd1 vccd1 _07328_ sky130_fd_sc_hd__nor2_1
Xhold1093 top.CPU.registers.data\[469\] vssd1 vssd1 vccd1 vccd1 net3650 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07513__X _03152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13074__A0 top.CPU.data_out\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11833_ net470 _06664_ net240 net154 net2724 vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__a32o_1
XANTENNA__09817__A1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11035__X _06577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11764_ _06607_ net235 net160 net3516 vssd1 vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_99_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_161_Right_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13503_ top.CPU.data_out\[10\] net587 _02969_ _02971_ vssd1 vssd1 vccd1 vccd1 _02508_
+ sky130_fd_sc_hd__o22a_1
X_10715_ _06328_ _06329_ _06327_ vssd1 vssd1 vccd1 vccd1 _06330_ sky130_fd_sc_hd__o21ai_1
XFILLER_159_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11695_ net1403 net542 net498 vssd1 vssd1 vccd1 vccd1 _06758_ sky130_fd_sc_hd__nand3_1
XFILLER_9_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16222_ net2556 _02432_ net1204 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[1022\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_146_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13434_ top.CPU.control_unit.instruction\[12\] net1399 net872 vssd1 vssd1 vccd1 vccd1
+ _02937_ sky130_fd_sc_hd__o21a_2
XFILLER_173_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10646_ _06090_ _06263_ net399 vssd1 vssd1 vccd1 vccd1 _06264_ sky130_fd_sc_hd__mux2_1
XANTENNA__08491__S net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14474__644 clknet_leaf_151_clk vssd1 vssd1 vccd1 vccd1 net2113 sky130_fd_sc_hd__inv_2
XANTENNA__11388__B1 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11927__A2 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16153_ net2487 _02363_ net1245 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[953\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_155_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13365_ net1389 _02892_ net671 vssd1 vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_102_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_102_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_154_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10577_ _06162_ _06197_ net310 vssd1 vssd1 vccd1 vccd1 _06198_ sky130_fd_sc_hd__mux2_1
XANTENNA__11211__A _06428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15104_ net1486 _01317_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r2_prev\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_12316_ net2574 _03645_ net1149 vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__mux2_1
X_16084_ net2418 _02294_ net1072 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[884\]
+ sky130_fd_sc_hd__dfrtp_1
X_13296_ top.mmio.mem_data_i\[17\] top.mmio.mem_data_i\[19\] top.mmio.mem_data_i\[18\]
+ top.mmio.mem_data_i\[16\] vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_110_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15035_ clknet_leaf_91_clk _01280_ net1270 vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_110_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14515__685 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 net2154 sky130_fd_sc_hd__inv_2
XANTENNA__12741__S net1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12247_ net3390 net134 net433 vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__mux2_1
XANTENNA__09202__C1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12178_ _03181_ net462 net540 _06751_ vssd1 vssd1 vccd1 vccd1 _06857_ sky130_fd_sc_hd__or4_1
XANTENNA__11560__B1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07764__C1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11129_ net497 net461 _06622_ net301 net3108 vssd1 vssd1 vccd1 vccd1 _02288_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_147_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12104__A2 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09505__B1 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_169_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_169_clk
+ sky130_fd_sc_hd__clkbuf_8
X_15937_ net2271 _02147_ net1230 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[737\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_37_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15868_ net2202 _02078_ net1235 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[668\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13065__A0 top.CPU.data_out\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14838__1008 clknet_leaf_180_clk vssd1 vssd1 vccd1 vccd1 net2477 sky130_fd_sc_hd__inv_2
X_15799_ net2133 _02009_ net1185 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[599\]
+ sky130_fd_sc_hd__dfrtp_1
X_08340_ top.CPU.registers.data_out_r2_prev\[19\] net687 net620 _03976_ _03978_ vssd1
+ vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__o2111a_1
XFILLER_149_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08271_ _03908_ _03909_ net947 vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08492__B1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09036__A2 net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11379__B1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10944__B _05693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11918__A2 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13320__B net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07598__A2 net1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10051__B1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12879__A0 top.CPU.alu.program_counter\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10960__A net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08547__A1 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1029_A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout391_A net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout125 net127 vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__buf_2
XFILLER_102_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout136 _05879_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout489_A net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout147 _06391_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__buf_2
Xfanout158 net159 vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__buf_2
Xfanout169 net171 vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__clkbuf_8
X_07986_ net933 _03624_ vssd1 vssd1 vccd1 vccd1 _03625_ sky130_fd_sc_hd__or2_1
X_13847__17 clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 net1486 sky130_fd_sc_hd__inv_2
X_09725_ _05363_ vssd1 vssd1 vccd1 vccd1 _05364_ sky130_fd_sc_hd__inv_2
XFILLER_28_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout656_A net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout277_X net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1398_A net1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09656_ _03988_ _03989_ vssd1 vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__and2_1
XFILLER_16_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08607_ top.CPU.registers.data\[687\] net1286 vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__or2_1
XFILLER_63_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout823_A net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09587_ top.CPU.registers.data_out_r2_prev\[0\] net686 net605 _05225_ _05209_ vssd1
+ vssd1 vccd1 vccd1 _05226_ sky130_fd_sc_hd__o221a_4
XANTENNA_fanout444_X net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08538_ top.CPU.registers.data\[752\] net1378 net984 top.CPU.registers.data\[720\]
+ net909 vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__a221o_1
XFILLER_169_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14161__331 clknet_leaf_179_clk vssd1 vssd1 vccd1 vccd1 net1800 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11082__A2 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08469_ top.CPU.registers.data\[561\] top.CPU.registers.data\[529\] net995 vssd1
+ vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout611_X net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14458__628 clknet_leaf_164_clk vssd1 vssd1 vccd1 vccd1 net2097 sky130_fd_sc_hd__inv_2
XANTENNA__09680__C1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout709_X net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10500_ net600 _06124_ vssd1 vssd1 vccd1 vccd1 _06125_ sky130_fd_sc_hd__nor2_1
XFILLER_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12016__D1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11480_ _06610_ net261 net257 net3628 vssd1 vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__a22o_1
XANTENNA__11909__A2 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14202__372 clknet_leaf_166_clk vssd1 vssd1 vccd1 vccd1 net1841 sky130_fd_sc_hd__inv_2
XANTENNA__08235__B1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10431_ net3853 net228 net313 _06058_ vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__a22o_1
XFILLER_109_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10042__B1 _05680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11031__A _03180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07589__A2 net1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13150_ net126 _02740_ _02741_ _02739_ top.CPU.alu.program_counter\[0\] vssd1 vssd1
+ vccd1 vccd1 _01297_ sky130_fd_sc_hd__a32o_1
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10362_ _03922_ _04057_ _05966_ _05967_ net446 vssd1 vssd1 vccd1 vccd1 _05992_ sky130_fd_sc_hd__o311a_1
XANTENNA_fanout980_X net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13657__S net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11790__B1 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12101_ net3960 net649 _06818_ vssd1 vssd1 vccd1 vccd1 _01512_ sky130_fd_sc_hd__o21a_1
XANTENNA__07994__C1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10293_ _05924_ _05925_ net402 vssd1 vssd1 vccd1 vccd1 _05926_ sky130_fd_sc_hd__mux2_1
X_13081_ top.CPU.data_out\[16\] net2898 net560 vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10870__A net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12032_ _06149_ net3574 net150 vssd1 vssd1 vccd1 vccd1 _01554_ sky130_fd_sc_hd__mux2_1
Xhold190 top.CPU.registers.data\[681\] vssd1 vssd1 vccd1 vccd1 net2747 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10896__A2 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout670 net671 vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09723__X _05362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout681 net684 vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12098__A1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout692 net694 vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__buf_4
XFILLER_46_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15722_ net2056 _01932_ net1090 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[522\]
+ sky130_fd_sc_hd__dfrtp_1
X_12934_ top.CPU.alu.program_counter\[29\] _03477_ vssd1 vssd1 vccd1 vccd1 _07375_
+ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09171__A net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13861__31 clknet_leaf_109_clk vssd1 vssd1 vccd1 vccd1 net1500 sky130_fd_sc_hd__inv_2
X_15653_ net1987 _01863_ net1083 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[453\]
+ sky130_fd_sc_hd__dfrtp_1
X_12865_ top.CPU.alu.program_counter\[22\] top.CPU.alu.program_counter\[21\] _07298_
+ vssd1 vssd1 vccd1 vccd1 _07313_ sky130_fd_sc_hd__and3_1
XANTENNA__11206__A net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11816_ _06500_ _06648_ net236 net156 net3136 vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__a32o_1
XANTENNA__10110__A _03476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15584_ net1918 _01794_ net1092 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[384\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ top.CPU.alu.program_counter\[15\] _07250_ net1362 vssd1 vssd1 vccd1 vccd1
+ _01178_ sky130_fd_sc_hd__mux2_1
XANTENNA__09266__A2 net1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _06589_ net498 net192 net3268 vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__a22o_1
XFILLER_53_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11678_ net462 _06495_ net237 net165 net2958 vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__a32o_1
X_16205_ net2539 _02415_ net1069 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[1005\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_146_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13417_ net67 top.mmio.mem_data_i\[30\] net598 vssd1 vssd1 vccd1 vccd1 _02930_ sky130_fd_sc_hd__o21a_1
X_10629_ _04533_ net508 net503 _04535_ net443 vssd1 vssd1 vccd1 vccd1 _06248_ sky130_fd_sc_hd__o221a_1
XANTENNA__08226__B1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08321__S0 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16136_ net2470 _02346_ net1088 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[936\]
+ sky130_fd_sc_hd__dfrtp_1
X_13348_ top.I2C.data_out\[11\] net553 _02879_ net596 vssd1 vssd1 vccd1 vccd1 _02880_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10584__A1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11781__B1 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16067_ net2401 _02277_ net1207 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[867\]
+ sky130_fd_sc_hd__dfrtp_1
X_13279_ _07054_ _02825_ net634 vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_149_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10780__A net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15018_ clknet_leaf_98_clk _01263_ net1254 vssd1 vssd1 vccd1 vccd1 top.SPI.parameters\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09346__A net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11595__B net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11533__B1 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16240__Q top.CPU.control_unit.instruction\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_68_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07840_ top.CPU.registers.data\[29\] net979 _03478_ vssd1 vssd1 vccd1 vccd1 _03479_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_127_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12089__A1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07771_ top.CPU.registers.data\[318\] top.CPU.registers.data\[286\] top.CPU.registers.data\[62\]
+ top.CPU.registers.data\[30\] net996 net621 vssd1 vssd1 vccd1 vccd1 _03410_ sky130_fd_sc_hd__mux4_1
XANTENNA__10004__B _05616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10779__X _06391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13825__A2 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11815__S net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15281__RESET_B net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09510_ top.CPU.registers.data\[321\] net1307 net1030 top.CPU.registers.data\[353\]
+ net947 vssd1 vssd1 vccd1 vccd1 _05149_ sky130_fd_sc_hd__a221o_1
XANTENNA__11836__A1 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08162__C1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09441_ top.CPU.registers.data\[802\] top.CPU.registers.data\[770\] net986 vssd1
+ vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_140_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14145__315 clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 net1784 sky130_fd_sc_hd__inv_2
XANTENNA__11116__A net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09372_ net939 _05003_ _05004_ net607 vssd1 vssd1 vccd1 vccd1 _05011_ sky130_fd_sc_hd__a31o_1
XANTENNA__09257__A2 net1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08323_ top.CPU.registers.data\[339\] net1296 net1016 top.CPU.registers.data\[371\]
+ net938 vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__a221o_1
XANTENNA__12261__A1 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08465__B1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10955__A net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout237_A net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08254_ top.CPU.registers.data\[982\] net1299 net1021 top.CPU.registers.data\[1014\]
+ net918 vssd1 vssd1 vccd1 vccd1 _03893_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_31_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10674__B _06290_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12013__A1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08185_ top.CPU.registers.data\[55\] net1017 net936 vssd1 vssd1 vccd1 vccd1 _03824_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__09414__C1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout404_A net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1146_A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08768__A1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11772__B1 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1313_A net1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13513__B2 _02976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07991__A2 net1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10327__B2 top.CPU.handler.toreg\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout773_A net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11524__B1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07728__C1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08940__A1 net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout561_X net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout940_A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07969_ top.CPU.control_unit.instruction\[16\] _03607_ _03605_ vssd1 vssd1 vccd1
+ vccd1 _03608_ sky130_fd_sc_hd__o21a_1
XFILLER_75_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout659_X net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13506__A _04459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09708_ top.CPU.registers.data\[761\] net1385 net1001 top.CPU.registers.data\[729\]
+ net922 vssd1 vssd1 vccd1 vccd1 _05347_ sky130_fd_sc_hd__a221o_1
XFILLER_114_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10980_ net3326 net218 _06542_ net316 vssd1 vssd1 vccd1 vccd1 _02357_ sky130_fd_sc_hd__a22o_1
XFILLER_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09639_ _04664_ _04730_ _04665_ vssd1 vssd1 vccd1 vccd1 _05278_ sky130_fd_sc_hd__a21o_1
XFILLER_16_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11026__A net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12650_ _07118_ net3982 top.I2C.output_state\[7\] vssd1 vssd1 vccd1 vccd1 _00004_
+ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_48_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11601_ _06479_ net428 net209 net215 net2817 vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__a32o_1
XANTENNA__13512__Y _02976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12252__A1 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12581_ top.CPU.addressnew\[11\] top.CPU.addressnew\[13\] top.CPU.addressnew\[15\]
+ top.CPU.addressnew\[14\] vssd1 vssd1 vccd1 vccd1 _07085_ sky130_fd_sc_hd__or4_1
XANTENNA__14933__RESET_B net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10865__A net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14909__1079 clknet_leaf_134_clk vssd1 vssd1 vccd1 vccd1 net2548 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11460__S net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13241__A top.I2C.output_state\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11532_ _06655_ net259 net250 net3385 vssd1 vssd1 vccd1 vccd1 _01999_ sky130_fd_sc_hd__a22o_1
XFILLER_157_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09405__C1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11463_ net144 net3404 net264 vssd1 vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__mux2_1
XFILLER_137_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13202_ top.I2C.data_out\[18\] net892 _02780_ vssd1 vssd1 vccd1 vccd1 _02781_ sky130_fd_sc_hd__mux2_1
X_10414_ net406 _06041_ vssd1 vssd1 vccd1 vccd1 _06042_ sky130_fd_sc_hd__nor2_1
XFILLER_171_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10566__A1 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11394_ _06516_ net280 net273 net3365 vssd1 vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__a22o_1
XFILLER_87_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09420__A2 net1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11763__B1 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07967__C1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13133_ net2653 _02735_ _02734_ vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__mux2_1
XANTENNA__12497__A1_N _05154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10345_ _05911_ _05975_ net308 vssd1 vssd1 vccd1 vccd1 _05976_ sky130_fd_sc_hd__mux2_1
XFILLER_152_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14837__1007 clknet_leaf_172_clk vssd1 vssd1 vccd1 vccd1 net2476 sky130_fd_sc_hd__inv_2
XANTENNA__09708__B1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13064_ net3077 top.CPU.data_out\[11\] net557 vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__mux2_1
X_10276_ _03649_ _05300_ _05367_ vssd1 vssd1 vccd1 vccd1 _05909_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14586__756 clknet_leaf_163_clk vssd1 vssd1 vccd1 vccd1 net2225 sky130_fd_sc_hd__inv_2
XANTENNA__09184__A1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1410 top.SPI.state\[0\] vssd1 vssd1 vccd1 vccd1 net1410 sky130_fd_sc_hd__clkbuf_4
X_12015_ net4002 net656 _06784_ vssd1 vssd1 vccd1 vccd1 _01564_ sky130_fd_sc_hd__o21a_1
XFILLER_78_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10869__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_161_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14627__797 clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 net2266 sky130_fd_sc_hd__inv_2
XFILLER_93_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10759__B _06371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12917_ _07355_ _07359_ vssd1 vssd1 vccd1 vccd1 _07360_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_122_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15705_ net2039 _01915_ net1238 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[505\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08695__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11294__A2 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12848_ top.CPU.alu.program_counter\[20\] _07287_ vssd1 vssd1 vccd1 vccd1 _07298_
+ sky130_fd_sc_hd__and2_1
X_15636_ net1970 _01846_ net1119 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[436\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09239__A2 net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15567_ net1901 _01777_ net1096 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[367\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08447__B1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12779_ _07213_ _07224_ vssd1 vssd1 vccd1 vccd1 _07235_ sky130_fd_sc_hd__nor2_1
XFILLER_9_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08516__Y _04155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15498_ net1832 _01708_ net1088 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[298\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_174_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16235__Q top.CPU.control_unit.instruction\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_80_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_662 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold904 top.CPU.registers.data\[604\] vssd1 vssd1 vccd1 vccd1 net3461 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_156_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11102__C net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold915 top.CPU.registers.data\[279\] vssd1 vssd1 vccd1 vccd1 net3472 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09411__A2 net1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14530__700 clknet_leaf_146_clk vssd1 vssd1 vccd1 vccd1 net2169 sky130_fd_sc_hd__inv_2
XANTENNA__11754__B1 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07958__C1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold926 top.CPU.registers.data\[760\] vssd1 vssd1 vccd1 vccd1 net3483 sky130_fd_sc_hd__dlygate4sd3_1
X_16119_ net2453 _02329_ net1173 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[919\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold937 top.CPU.registers.data\[766\] vssd1 vssd1 vccd1 vccd1 net3494 sky130_fd_sc_hd__dlygate4sd3_1
Xhold948 top.CPU.registers.data\[254\] vssd1 vssd1 vccd1 vccd1 net3505 sky130_fd_sc_hd__dlygate4sd3_1
X_09990_ _04987_ net372 vssd1 vssd1 vccd1 vccd1 _05629_ sky130_fd_sc_hd__nor2_1
Xhold959 top.CPU.registers.data\[381\] vssd1 vssd1 vccd1 vccd1 net3516 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_170_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09076__A net1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08941_ top.CPU.registers.data\[554\] top.CPU.registers.data\[522\] net971 vssd1
+ vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__mux2_1
XANTENNA__10309__A1 _05332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11506__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12214__B net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15462__RESET_B net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08872_ top.CPU.registers.data\[43\] top.CPU.registers.data\[11\] net808 vssd1 vssd1
+ vccd1 vccd1 _04511_ sky130_fd_sc_hd__mux2_1
XANTENNA__08922__A1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07823_ top.CPU.registers.data\[93\] net1319 net849 top.CPU.registers.data\[125\]
+ net768 vssd1 vssd1 vccd1 vccd1 _03462_ sky130_fd_sc_hd__a221o_1
XANTENNA__13326__A _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07754_ top.CPU.registers.data\[254\] net1394 net834 top.CPU.registers.data\[222\]
+ net781 vssd1 vssd1 vccd1 vccd1 _03393_ sky130_fd_sc_hd__a221o_1
XANTENNA__08135__C1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07685_ net632 _03318_ _03323_ vssd1 vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout354_A net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_91_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_91_clk sky130_fd_sc_hd__clkbuf_8
X_09424_ net954 _05062_ _05061_ net612 vssd1 vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__a211o_1
X_09355_ top.CPU.registers.data\[803\] top.CPU.registers.data\[771\] net990 vssd1
+ vssd1 vccd1 vccd1 _04994_ sky130_fd_sc_hd__mux2_1
XANTENNA__08438__B1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout142_X net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout521_A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout619_A net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08306_ top.CPU.registers.data\[979\] net1325 net856 top.CPU.registers.data\[1011\]
+ net724 vssd1 vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__a221o_1
XFILLER_139_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09286_ top.CPU.registers.data\[932\] top.CPU.registers.data\[900\] top.CPU.registers.data\[804\]
+ top.CPU.registers.data\[772\] net989 net914 vssd1 vssd1 vccd1 vccd1 _04925_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_43_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10796__A1 _05754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_7_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11993__B1 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08237_ top.CPU.registers.data\[982\] net1330 net861 top.CPU.registers.data\[1014\]
+ net728 vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_60_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout407_X net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12203__C_N _06796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08168_ top.CPU.registers.data\[855\] net1325 net856 top.CPU.registers.data\[887\]
+ net749 vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__a221o_1
XANTENNA__09402__A2 net1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11745__B1 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout988_A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14273__443 clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 net1912 sky130_fd_sc_hd__inv_2
XFILLER_134_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08610__B1 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08099_ net752 _03733_ _03734_ _03737_ net637 vssd1 vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__a311o_1
XFILLER_133_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1316_X net1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10130_ net601 _05767_ vssd1 vssd1 vccd1 vccd1 _05768_ sky130_fd_sc_hd__and2_1
XFILLER_0_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07964__A2 net1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout776_X net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10061_ _05514_ net447 _05698_ vssd1 vssd1 vccd1 vccd1 _05699_ sky130_fd_sc_hd__and3_1
XFILLER_0_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14314__484 clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 net1953 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_89_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08374__C1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout943_X net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13820_ net2894 net334 net328 top.CPU.data_out\[22\] vssd1 vssd1 vccd1 vccd1 _02700_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12140__A net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13751_ top.SPI.timem\[22\] _03085_ vssd1 vssd1 vccd1 vccd1 _03087_ sky130_fd_sc_hd__nand2_1
XANTENNA__11276__A2 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08677__B1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10963_ net530 _06532_ vssd1 vssd1 vccd1 vccd1 _06533_ sky130_fd_sc_hd__nor2_1
XANTENNA__13670__B1 _03048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12702_ top.CPU.alu.program_counter\[6\] _07152_ top.CPU.alu.program_counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 _07165_ sky130_fd_sc_hd__a21oi_1
X_16470_ clknet_leaf_88_clk _02632_ net1272 vssd1 vssd1 vccd1 vccd1 top.SPI.timem\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_13682_ net2634 net336 vssd1 vssd1 vccd1 vccd1 _02610_ sky130_fd_sc_hd__and2_1
XANTENNA__08764__S net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08617__X _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10894_ net3732 net222 _06490_ net466 vssd1 vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__a22o_1
XFILLER_44_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15421_ net1755 _01631_ net1112 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[221\]
+ sky130_fd_sc_hd__dfrtp_1
X_12633_ top.I2C.byte_manager_state\[2\] top.I2C.output_state\[14\] _06912_ vssd1
+ vssd1 vccd1 vccd1 _00014_ sky130_fd_sc_hd__and3_1
XANTENNA__08429__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15352_ net1686 _01562_ net1150 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[152\]
+ sky130_fd_sc_hd__dfrtp_1
X_12564_ _06410_ _06426_ _06445_ vssd1 vssd1 vccd1 vccd1 _07069_ sky130_fd_sc_hd__and3b_1
XFILLER_8_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11984__B1 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11515_ _05809_ net429 net258 _06735_ vssd1 vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__a31o_1
XANTENNA__07652__A1 net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15283_ net1617 _01493_ net1175 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[83\]
+ sky130_fd_sc_hd__dfrtp_1
X_12495_ _05084_ _05120_ vssd1 vssd1 vccd1 vccd1 _07004_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_22_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09595__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09448__X _05087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_44_Left_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11446_ _03193_ _06033_ net538 vssd1 vssd1 vccd1 vccd1 _06723_ sky130_fd_sc_hd__and3_1
XFILLER_109_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11736__B1 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11200__A2 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11377_ _06492_ net280 net273 net3298 vssd1 vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__a22o_1
XFILLER_153_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13116_ top.SPI.command\[4\] net1410 top.SPI.paroutput\[28\] net1358 vssd1 vssd1
+ vccd1 vccd1 _02723_ sky130_fd_sc_hd__a22o_1
XFILLER_98_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10328_ _05690_ _05958_ _05959_ vssd1 vssd1 vccd1 vccd1 _05960_ sky130_fd_sc_hd__o21ba_2
XANTENNA__13489__A0 top.CPU.data_out\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_163_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ top.SPI.parameters\[25\] top.SPI.paroutput\[17\] net1357 vssd1 vssd1 vccd1
+ vccd1 _07449_ sky130_fd_sc_hd__mux2_1
X_10259_ net413 _05888_ _05892_ _05618_ _05884_ vssd1 vssd1 vccd1 vccd1 _05893_ sky130_fd_sc_hd__o221a_1
XFILLER_79_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1240 net1276 vssd1 vssd1 vccd1 vccd1 net1240 sky130_fd_sc_hd__buf_2
XFILLER_61_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12700__A2 _03118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1251 net1252 vssd1 vssd1 vccd1 vccd1 net1251 sky130_fd_sc_hd__buf_2
Xfanout1262 net1276 vssd1 vssd1 vccd1 vccd1 net1262 sky130_fd_sc_hd__clkbuf_2
Xfanout1273 net1275 vssd1 vssd1 vccd1 vccd1 net1273 sky130_fd_sc_hd__clkbuf_4
XFILLER_38_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_53_Left_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1284 net1285 vssd1 vssd1 vccd1 vccd1 net1284 sky130_fd_sc_hd__buf_2
XANTENNA__08380__A2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13146__A top.CPU.alu.program_counter\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1295 net1301 vssd1 vssd1 vccd1 vccd1 net1295 sky130_fd_sc_hd__buf_2
X_14998_ clknet_leaf_94_clk _01243_ net1261 vssd1 vssd1 vccd1 vccd1 top.SPI.parameters\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12464__A1 _05330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08668__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12464__B2 _05498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_73_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_35_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08132__A2 net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07470_ top.CPU.control_unit.instruction\[16\] vssd1 vssd1 vccd1 vccd1 _03110_ sky130_fd_sc_hd__inv_2
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15619_ net1953 _01829_ net1208 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[419\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11019__A2 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09617__C1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09140_ top.CPU.registers.data\[295\] top.CPU.registers.data\[263\] net997 vssd1
+ vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_174_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11975__B1 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_62_Left_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09071_ _04708_ _04709_ net672 vssd1 vssd1 vccd1 vccd1 _04710_ sky130_fd_sc_hd__o21a_1
XFILLER_163_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14257__427 clknet_leaf_190_clk vssd1 vssd1 vccd1 vccd1 net1896 sky130_fd_sc_hd__inv_2
X_08022_ net791 _03656_ _03657_ net743 vssd1 vssd1 vccd1 vccd1 _03661_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_135_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold701 top.CPU.registers.data\[949\] vssd1 vssd1 vccd1 vccd1 net3258 sky130_fd_sc_hd__dlygate4sd3_1
Xhold712 top.CPU.registers.data\[202\] vssd1 vssd1 vccd1 vccd1 net3269 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11727__B1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold723 top.SPI.counter\[2\] vssd1 vssd1 vccd1 vccd1 net3280 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08199__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold734 top.CPU.registers.data\[249\] vssd1 vssd1 vccd1 vccd1 net3291 sky130_fd_sc_hd__dlygate4sd3_1
X_14001__171 clknet_leaf_190_clk vssd1 vssd1 vccd1 vccd1 net1640 sky130_fd_sc_hd__inv_2
Xhold745 top.CPU.registers.data\[231\] vssd1 vssd1 vccd1 vccd1 net3302 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold756 net63 vssd1 vssd1 vccd1 vccd1 net3313 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07946__A2 net1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold767 top.CPU.registers.data\[724\] vssd1 vssd1 vccd1 vccd1 net3324 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11742__A3 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold778 top.CPU.registers.data\[284\] vssd1 vssd1 vccd1 vccd1 net3335 sky130_fd_sc_hd__dlygate4sd3_1
X_09973_ _05512_ _05611_ vssd1 vssd1 vccd1 vccd1 _05612_ sky130_fd_sc_hd__nor2_1
XFILLER_118_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold789 top.CPU.registers.data\[518\] vssd1 vssd1 vccd1 vccd1 net3346 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08924_ top.CPU.registers.data\[970\] net1313 net844 top.CPU.registers.data\[1002\]
+ net765 vssd1 vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__a221o_1
XFILLER_39_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1011_A net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12152__B1 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09699__A2 net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1401 top.CPU.registers.data\[599\] vssd1 vssd1 vccd1 vccd1 net3958 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1109_A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14908__1078 clknet_leaf_137_clk vssd1 vssd1 vccd1 vccd1 net2547 sky130_fd_sc_hd__inv_2
XFILLER_58_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_71_Left_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1412 top.I2C.output_state\[13\] vssd1 vssd1 vccd1 vccd1 net3969 sky130_fd_sc_hd__dlygate4sd3_1
X_08855_ net1283 _04492_ _04493_ vssd1 vssd1 vccd1 vccd1 _04494_ sky130_fd_sc_hd__or3_1
XANTENNA__10702__A1 _05664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1423 top.I2C.data_out\[6\] vssd1 vssd1 vccd1 vccd1 net3980 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout471_A net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1434 top.CPU.registers.data\[97\] vssd1 vssd1 vccd1 vccd1 net3991 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1445 top.CPU.registers.data\[154\] vssd1 vssd1 vccd1 vccd1 net4002 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1456 top.SPI.timem\[10\] vssd1 vssd1 vccd1 vccd1 net4013 sky130_fd_sc_hd__dlygate4sd3_1
X_07806_ _03442_ _03443_ vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1467 top.SPI.command\[0\] vssd1 vssd1 vccd1 vccd1 net4024 sky130_fd_sc_hd__dlygate4sd3_1
X_08786_ net692 _04423_ _04424_ vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__or3_1
XFILLER_55_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07737_ top.CPU.alu.program_counter\[30\] net1036 vssd1 vssd1 vccd1 vccd1 _03376_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__08659__B1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12895__A top.CPU.alu.program_counter\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1380_A net1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_64_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout357_X net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07668_ _03271_ _03283_ net632 _03297_ _03304_ vssd1 vssd1 vccd1 vccd1 _03307_ sky130_fd_sc_hd__o2111a_1
XANTENNA__11007__C net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09407_ top.CPU.registers.data\[547\] top.CPU.registers.data\[515\] net828 vssd1
+ vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__mux2_1
X_14836__1006 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 net2475 sky130_fd_sc_hd__inv_2
XFILLER_71_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12207__A1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09608__C1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout903_A net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout524_X net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07599_ net779 _03236_ _03237_ vssd1 vssd1 vccd1 vccd1 _03238_ sky130_fd_sc_hd__or3_1
X_09338_ net708 _04973_ _04974_ net643 vssd1 vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_80_Left_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11966__B1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09269_ top.CPU.registers.data\[677\] top.CPU.registers.data\[645\] top.CPU.registers.data\[549\]
+ top.CPU.registers.data\[517\] net966 net901 vssd1 vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__mux4_1
X_11300_ _05960_ _06705_ net290 net3412 vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__a2bb2o_1
X_12280_ net2609 _05465_ net1253 vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__mux2_1
XANTENNA__09709__A net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11718__B1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10862__B net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11231_ net3585 net294 _06670_ net314 vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__a22o_1
XFILLER_20_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15313__RESET_B net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11162_ net480 net457 _06641_ net301 net3026 vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__a32o_1
XANTENNA__11733__A3 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10113_ net384 _05750_ _05749_ net396 vssd1 vssd1 vccd1 vccd1 _05751_ sky130_fd_sc_hd__a211oi_1
XFILLER_1_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15970_ net2304 _02180_ net1173 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[770\]
+ sky130_fd_sc_hd__dfrtp_1
X_11093_ net1404 net551 net472 _06603_ vssd1 vssd1 vccd1 vccd1 _06604_ sky130_fd_sc_hd__or4_4
XANTENNA__12789__B _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input32_A DAT_I[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10044_ _05617_ _05641_ _05642_ _05662_ _05682_ vssd1 vssd1 vccd1 vccd1 _05683_ sky130_fd_sc_hd__a221o_1
X_14921_ clknet_leaf_30_clk _01167_ net1152 vssd1 vssd1 vccd1 vccd1 top.CPU.alu.program_counter\[4\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold50 top.mmio.m1 vssd1 vssd1 vccd1 vccd1 net2607 sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 top.CPU.registers.data_out_r2_prev\[4\] vssd1 vssd1 vccd1 vccd1 net2618 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08362__A2 net1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold72 top.CPU.registers.data_out_r1_prev\[13\] vssd1 vssd1 vccd1 vccd1 net2629 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold83 net43 vssd1 vssd1 vccd1 vccd1 net2640 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_21_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold94 top.CPU.registers.data\[294\] vssd1 vssd1 vccd1 vccd1 net2651 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07570__B1 _03111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13803_ net3834 net333 net326 net3666 vssd1 vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__a22o_1
XFILLER_28_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11995_ _06561_ net350 net182 net2868 vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__a22o_1
XANTENNA__09847__C1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_55_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_16_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09311__A1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13734_ top.SPI.timem\[15\] _03074_ net3896 vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__a21oi_1
X_16522_ clknet_leaf_99_clk _02684_ net1256 vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__dfrtp_1
X_14698__868 clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 net2337 sky130_fd_sc_hd__inv_2
X_10946_ net130 net437 vssd1 vssd1 vccd1 vccd1 _06522_ sky130_fd_sc_hd__and2_1
XANTENNA__08347__X _03986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_119_Left_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16453_ clknet_leaf_81_clk _02616_ net1242 vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__dfrtp_1
X_13665_ _03045_ _03046_ vssd1 vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__nor2_4
X_10877_ net661 _05906_ _06471_ vssd1 vssd1 vccd1 vccd1 _06479_ sky130_fd_sc_hd__and3_1
X_12616_ _07101_ _07111_ net1354 vssd1 vssd1 vccd1 vccd1 _07115_ sky130_fd_sc_hd__o21ai_1
X_15404_ net1738 _01614_ net1070 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[204\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_156_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16384_ clknet_leaf_62_clk _02593_ net1163 vssd1 vssd1 vccd1 vccd1 top.CPU.fetch.current_ra\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09075__B1 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13596_ top.CPU.addressnew\[19\] net578 vssd1 vssd1 vccd1 vccd1 _03024_ sky130_fd_sc_hd__nand2_1
XFILLER_129_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09614__A2 net1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11957__B1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15335_ net1669 _01545_ net1198 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[135\]
+ sky130_fd_sc_hd__dfrtp_1
X_12547_ net1353 _03246_ vssd1 vssd1 vccd1 vccd1 _07056_ sky130_fd_sc_hd__nand2_1
XFILLER_12_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11421__A2 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15266_ net1600 _01476_ net1177 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[66\]
+ sky130_fd_sc_hd__dfrtp_1
X_12478_ _06980_ _06981_ vssd1 vssd1 vccd1 vccd1 _06987_ sky130_fd_sc_hd__nor2_1
XANTENNA_3 _06714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11709__B1 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09378__A1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11429_ _06573_ net276 net267 net3733 vssd1 vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__a22o_1
XFILLER_6_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15197_ clknet_leaf_87_clk _01407_ net1271 vssd1 vssd1 vccd1 vccd1 top.SPI.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11185__A1 net1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07928__A2 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08338__C1 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12134__B1 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11488__A2 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14642__812 clknet_leaf_201_clk vssd1 vssd1 vccd1 vccd1 net2281 sky130_fd_sc_hd__inv_2
Xfanout1070 net1075 vssd1 vssd1 vccd1 vccd1 net1070 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09550__A1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08640_ top.CPU.registers.data\[174\] top.CPU.registers.data\[142\] net819 vssd1
+ vssd1 vccd1 vccd1 _04279_ sky130_fd_sc_hd__mux2_1
XFILLER_67_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1081 net1082 vssd1 vssd1 vccd1 vccd1 net1081 sky130_fd_sc_hd__clkbuf_4
Xfanout1092 net1093 vssd1 vssd1 vccd1 vccd1 net1092 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10160__A2 _05667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08571_ top.CPU.registers.data\[975\] net1315 net846 top.CPU.registers.data\[1007\]
+ net716 vssd1 vssd1 vccd1 vccd1 _04210_ sky130_fd_sc_hd__a221o_1
XANTENNA__11108__B net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09838__C1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_46_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08105__A2 net1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10448__B1 _05733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07522_ net1279 _03153_ vssd1 vssd1 vccd1 vccd1 _03161_ sky130_fd_sc_hd__nand2_2
XFILLER_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08510__C1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09853__A2 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11660__A2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11124__A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11948__B1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09123_ net800 _04754_ _04761_ net642 vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__a211o_1
XFILLER_157_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11412__A2 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08813__B1 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10963__A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout317_A net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1059_A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10620__B1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09054_ net785 _04688_ _04689_ net716 vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__o211a_1
X_08005_ net625 _03635_ _03643_ vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__and3_1
Xhold520 top.SPI.counter\[3\] vssd1 vssd1 vccd1 vccd1 net3077 sky130_fd_sc_hd__dlygate4sd3_1
Xhold531 top.SPI.paroutput\[18\] vssd1 vssd1 vccd1 vccd1 net3088 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold542 top.CPU.registers.data\[134\] vssd1 vssd1 vccd1 vccd1 net3099 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1226_A net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08577__C1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11176__B2 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold553 net86 vssd1 vssd1 vccd1 vccd1 net3110 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08041__A1 top.CPU.control_unit.instruction\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold564 net80 vssd1 vssd1 vccd1 vccd1 net3121 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10384__C1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold575 top.CPU.registers.data\[673\] vssd1 vssd1 vccd1 vccd1 net3132 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold586 _02694_ vssd1 vssd1 vccd1 vccd1 net3143 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold597 top.CPU.registers.data\[860\] vssd1 vssd1 vccd1 vccd1 net3154 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout686_A _03332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11794__A net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08592__A2 net1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09956_ _03650_ _05594_ vssd1 vssd1 vccd1 vccd1 _05595_ sky130_fd_sc_hd__nand2_1
XFILLER_89_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1014_X net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08329__C1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08907_ top.CPU.registers.data\[234\] net1387 net809 top.CPU.registers.data\[202\]
+ net765 vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__a221o_1
XFILLER_66_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09887_ _03407_ _03441_ vssd1 vssd1 vccd1 vccd1 _05526_ sky130_fd_sc_hd__nand2_1
XANTENNA__11479__A2 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1220 top.CPU.registers.data\[73\] vssd1 vssd1 vccd1 vccd1 net3777 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout474_X net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout853_A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1231 top.mmio.mem_data_i\[19\] vssd1 vssd1 vccd1 vccd1 net3788 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10687__B1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08838_ net624 _04473_ _04476_ vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__or3_1
X_14385__555 clknet_leaf_190_clk vssd1 vssd1 vccd1 vccd1 net2024 sky130_fd_sc_hd__inv_2
Xhold1242 top.CPU.registers.data\[698\] vssd1 vssd1 vccd1 vccd1 net3799 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_142_Right_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1253 top.I2C.data_out\[22\] vssd1 vssd1 vccd1 vccd1 net3810 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1264 top.CPU.registers.data\[46\] vssd1 vssd1 vccd1 vccd1 net3821 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1275 top.CPU.registers.data_out_r1_prev\[16\] vssd1 vssd1 vccd1 vccd1 net3832
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13625__A0 top.CPU.alu.program_counter\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1286 top.CPU.registers.data\[708\] vssd1 vssd1 vccd1 vccd1 net3843 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1297 top.CPU.registers.data\[763\] vssd1 vssd1 vccd1 vccd1 net3854 sky130_fd_sc_hd__dlygate4sd3_1
X_08769_ top.CPU.registers.data\[844\] net1316 net847 top.CPU.registers.data\[876\]
+ net742 vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout641_X net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12428__B2 top.I2C.output_state\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1383_X net1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout739_X net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_37_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__13514__A _04188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10439__B1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10800_ top.CPU.fetch.current_ra\[3\] net1040 net633 top.CPU.handler.toreg\[3\] vssd1
+ vssd1 vccd1 vccd1 _06411_ sky130_fd_sc_hd__a22o_1
X_11780_ _06623_ net196 net160 net3415 vssd1 vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__a22o_1
XFILLER_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14426__596 clknet_leaf_164_clk vssd1 vssd1 vccd1 vccd1 net2065 sky130_fd_sc_hd__inv_2
XFILLER_54_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10857__B net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09844__A2 net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10731_ net399 _06179_ _06139_ vssd1 vssd1 vccd1 vccd1 _06345_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_24_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11651__A2 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout906_X net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13450_ net3717 _02946_ net123 vssd1 vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__mux2_1
X_10662_ _06241_ _06278_ net306 vssd1 vssd1 vccd1 vccd1 _06279_ sky130_fd_sc_hd__mux2_1
XANTENNA__09057__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12401_ _03122_ net2632 net2608 vssd1 vssd1 vccd1 vccd1 _00037_ sky130_fd_sc_hd__a21o_1
X_13381_ top.I2C.data_out\[20\] net555 _02859_ top.mmio.mem_data_i\[20\] vssd1 vssd1
+ vccd1 vccd1 _02904_ sky130_fd_sc_hd__a22o_1
XANTENNA__08804__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11403__A2 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10593_ net572 net514 _06213_ vssd1 vssd1 vccd1 vccd1 _06214_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_97_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15120_ clknet_leaf_56_clk top.I2C.inter_received_n net1141 vssd1 vssd1 vccd1 vccd1
+ top.I2C.inter_received sky130_fd_sc_hd__dfrtp_1
X_12332_ net2573 _04727_ net1234 vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__mux2_1
XFILLER_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11954__A3 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10592__B net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15051_ clknet_leaf_91_clk _01296_ net1269 vssd1 vssd1 vccd1 vccd1 top.SPI.command\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_108_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12263_ net2999 _06311_ net431 vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__mux2_1
XFILLER_147_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11167__A1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11214_ net130 net3562 net297 vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_112_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12194_ top.CPU.registers.data\[54\] net655 net364 vssd1 vssd1 vccd1 vccd1 _06864_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_75_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput40 net40 vssd1 vssd1 vccd1 vccd1 ADR_O[10] sky130_fd_sc_hd__buf_2
XANTENNA__10914__A1 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput51 net51 vssd1 vssd1 vccd1 vccd1 ADR_O[20] sky130_fd_sc_hd__buf_2
XFILLER_150_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput62 net62 vssd1 vssd1 vccd1 vccd1 ADR_O[5] sky130_fd_sc_hd__buf_2
XANTENNA__09780__A1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 DAT_O[14] sky130_fd_sc_hd__buf_2
X_13993__163 clknet_leaf_157_clk vssd1 vssd1 vccd1 vccd1 net1632 sky130_fd_sc_hd__inv_2
X_11145_ net519 _06335_ vssd1 vssd1 vccd1 vccd1 _06632_ sky130_fd_sc_hd__nor2_1
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 DAT_O[24] sky130_fd_sc_hd__buf_2
XANTENNA__08489__S net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput95 net95 vssd1 vssd1 vccd1 vccd1 DAT_O[5] sky130_fd_sc_hd__buf_2
XANTENNA__07791__B1 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12116__B1 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_94_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15953_ net2287 _02163_ net1178 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[753\]
+ sky130_fd_sc_hd__dfrtp_1
X_11076_ net3392 net367 _06593_ net324 vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__a22o_1
XANTENNA__16353__RESET_B net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10027_ net408 _05664_ vssd1 vssd1 vccd1 vccd1 _05666_ sky130_fd_sc_hd__nor2_1
XFILLER_64_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15884_ net2218 _02094_ net1078 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[684\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08740__C1 net1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11890__A2 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_127_Left_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_28_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08099__A1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09296__B1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08077__X _03716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11978_ _06535_ net345 net181 net2903 vssd1 vssd1 vccd1 vccd1 _01594_ sky130_fd_sc_hd__a22o_1
XFILLER_16_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16505_ clknet_leaf_49_clk _02667_ net1128 vssd1 vssd1 vccd1 vccd1 top.mmio.mem_data_i\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13717_ net3990 _03062_ _03065_ _07113_ vssd1 vssd1 vccd1 vccd1 _02628_ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_152_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10929_ net3814 net222 _06511_ net464 vssd1 vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__a22o_1
XANTENNA__07846__A1 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11642__A2 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16436_ clknet_leaf_80_clk net2952 net1241 vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09048__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13648_ net3895 _07300_ net664 vssd1 vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_32_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_171_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13395__A2 _07089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14907__1077 clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 net2546 sky130_fd_sc_hd__inv_2
XFILLER_158_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16367_ clknet_leaf_62_clk _02576_ net1160 vssd1 vssd1 vccd1 vccd1 top.CPU.fetch.current_ra\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13579_ net1349 _06228_ vssd1 vssd1 vccd1 vccd1 _03014_ sky130_fd_sc_hd__nand2_1
XFILLER_75_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_167_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07568__S net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09349__A net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11945__A3 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15318_ net1652 _01528_ net1230 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[118\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_132_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16298_ clknet_leaf_108_clk _02507_ net1246 vssd1 vssd1 vccd1 vccd1 top.CPU.data_out\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_172_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_136_Left_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13147__A2 _02738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16243__Q top.CPU.control_unit.instruction\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_47_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15249_ net1583 _01459_ net1189 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11158__B2 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11110__C net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout307 _05158_ vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__clkbuf_2
X_09810_ net733 _05447_ _05448_ net638 vssd1 vssd1 vccd1 vccd1 _05449_ sky130_fd_sc_hd__a31o_1
XFILLER_28_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11818__S net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14835__1005 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 net2474 sky130_fd_sc_hd__inv_2
Xfanout318 net322 vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__buf_2
Xfanout329 _03096_ vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__clkbuf_4
X_14072__242 clknet_leaf_166_clk vssd1 vssd1 vccd1 vccd1 net1711 sky130_fd_sc_hd__inv_2
XFILLER_86_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09741_ top.CPU.registers.data\[443\] top.CPU.registers.data\[411\] net827 vssd1
+ vssd1 vccd1 vccd1 _05380_ sky130_fd_sc_hd__mux2_1
XANTENNA__09084__A net1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14369__539 clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 net2008 sky130_fd_sc_hd__inv_2
XFILLER_39_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08326__A2 net1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12122__A3 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_105_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09672_ net757 _05310_ _05309_ net698 vssd1 vssd1 vccd1 vccd1 _05311_ sky130_fd_sc_hd__o211a_1
XFILLER_27_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10133__A2 _05769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11330__A1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_145_Left_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14113__283 clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 net1752 sky130_fd_sc_hd__inv_2
XFILLER_36_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08623_ top.CPU.registers.data\[654\] net1320 net851 top.CPU.registers.data\[686\]
+ net720 vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__a221o_1
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_19_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__10958__A net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout267_A net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08554_ _04191_ _04192_ vssd1 vssd1 vccd1 vccd1 _04193_ sky130_fd_sc_hd__and2b_1
XANTENNA__09287__B1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07505_ top.CPU.control_unit.instruction\[3\] top.CPU.control_unit.instruction\[1\]
+ top.CPU.control_unit.instruction\[0\] vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__and3b_2
XFILLER_35_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07837__A1 _03474_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08485_ _04122_ _04123_ net455 vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__mux2_1
XANTENNA__11633__A2 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout434_A _06602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1176_A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10841__B1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_1038 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08862__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12892__B top.CPU.alu.program_counter\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout601_A net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14770__940 clknet_leaf_201_clk vssd1 vssd1 vccd1 vccd1 net2409 sky130_fd_sc_hd__inv_2
XANTENNA_fanout222_X net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09106_ net800 _04734_ _04735_ net729 vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__o211a_1
X_09037_ net740 _04668_ _04669_ net766 vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__o211a_1
XFILLER_151_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14811__981 clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 net2450 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_57_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11795__Y _06762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13977__147 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 net1616 sky130_fd_sc_hd__inv_2
XFILLER_117_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold350 top.CPU.registers.data\[409\] vssd1 vssd1 vccd1 vccd1 net2907 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout970_A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold361 top.CPU.registers.data\[534\] vssd1 vssd1 vccd1 vccd1 net2918 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09211__B1 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold372 top.CPU.registers.data\[439\] vssd1 vssd1 vccd1 vccd1 net2929 sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 top.CPU.registers.data\[600\] vssd1 vssd1 vccd1 vccd1 net2940 sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 net61 vssd1 vssd1 vccd1 vccd1 net2951 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_120_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout830 net831 vssd1 vssd1 vccd1 vccd1 net830 sky130_fd_sc_hd__buf_2
XANTENNA__07773__B1 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout841 net854 vssd1 vssd1 vccd1 vccd1 net841 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08970__C1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout852 net853 vssd1 vssd1 vccd1 vccd1 net852 sky130_fd_sc_hd__clkbuf_4
X_09939_ _03859_ _03922_ vssd1 vssd1 vccd1 vccd1 _05578_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout856_X net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout863 net864 vssd1 vssd1 vccd1 vccd1 net863 sky130_fd_sc_hd__clkbuf_4
XFILLER_133_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout874 net877 vssd1 vssd1 vccd1 vccd1 net874 sky130_fd_sc_hd__clkbuf_4
Xfanout885 _03095_ vssd1 vssd1 vccd1 vccd1 net885 sky130_fd_sc_hd__buf_2
Xclkbuf_4_13_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_13_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__11029__A net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout896 _07430_ vssd1 vssd1 vccd1 vccd1 net896 sky130_fd_sc_hd__buf_2
X_12950_ _07389_ vssd1 vssd1 vccd1 vccd1 _07390_ sky130_fd_sc_hd__inv_2
Xhold1050 _02602_ vssd1 vssd1 vccd1 vccd1 net3607 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11321__B2 _06354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1061 top.CPU.registers.data\[995\] vssd1 vssd1 vccd1 vccd1 net3618 sky130_fd_sc_hd__dlygate4sd3_1
X_11901_ net461 _06598_ vssd1 vssd1 vccd1 vccd1 _06771_ sky130_fd_sc_hd__nor2_2
Xhold1072 top.CPU.handler.toreg\[13\] vssd1 vssd1 vccd1 vccd1 net3629 sky130_fd_sc_hd__dlygate4sd3_1
X_12881_ top.CPU.alu.program_counter\[24\] _03646_ vssd1 vssd1 vccd1 vccd1 _07327_
+ sky130_fd_sc_hd__nor2_1
Xhold1083 top.CPU.registers.data\[773\] vssd1 vssd1 vccd1 vccd1 net3640 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1094 top.CPU.registers.data\[996\] vssd1 vssd1 vccd1 vccd1 net3651 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10868__A net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11463__S net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07540__A3 net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11832_ net469 _06663_ net241 net154 net3170 vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__a32o_1
XANTENNA__09278__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07828__A1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10079__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11763_ net470 _06606_ net240 net163 net3266 vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_99_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _04859_ _05275_ _05541_ net370 vssd1 vssd1 vccd1 vccd1 _06329_ sky130_fd_sc_hd__a31o_1
XANTENNA__10832__B1 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13502_ _04593_ _02967_ vssd1 vssd1 vccd1 vccd1 _02971_ sky130_fd_sc_hd__and2_1
XFILLER_9_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11694_ _06522_ net198 net164 net3056 vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__a22o_1
XFILLER_41_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13433_ net3736 _02870_ net120 vssd1 vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__mux2_1
X_16221_ net2555 _02431_ net1112 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[1021\]
+ sky130_fd_sc_hd__dfrtp_1
X_10645_ _06178_ _06262_ net388 vssd1 vssd1 vccd1 vccd1 _06263_ sky130_fd_sc_hd__mux2_1
XANTENNA__11388__A1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16152_ net2486 _02362_ net1150 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[952\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_155_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13364_ net889 _02891_ vssd1 vssd1 vccd1 vccd1 _02892_ sky130_fd_sc_hd__and2_1
XANTENNA__09450__A0 _05084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10576_ _04295_ _04364_ net376 vssd1 vssd1 vccd1 vccd1 _06197_ sky130_fd_sc_hd__mux2_1
XFILLER_5_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15103_ net1485 _01316_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r2_prev\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_12315_ net2593 _05361_ net1238 vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__mux2_1
XANTENNA__11211__B net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16083_ net2417 _02293_ net1177 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[883\]
+ sky130_fd_sc_hd__dfrtp_1
X_13295_ _02837_ vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__inv_2
XFILLER_142_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15034_ clknet_leaf_87_clk _01279_ net1271 vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_110_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12246_ net3457 _05961_ _06599_ vssd1 vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__mux2_1
X_14056__226 clknet_leaf_129_clk vssd1 vssd1 vccd1 vccd1 net1695 sky130_fd_sc_hd__inv_2
XANTENNA__08556__A2 net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13419__A _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12177_ net131 net354 net233 _06856_ vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__a31o_1
XFILLER_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11560__A1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11128_ net516 _06192_ vssd1 vssd1 vccd1 vccd1 _06622_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_147_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13301__A2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15936_ net2270 _02146_ net1090 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[736\]
+ sky130_fd_sc_hd__dfrtp_1
X_11059_ net325 net146 net536 net367 net2813 vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__a32o_1
XFILLER_83_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11312__B2 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15867_ net2201 _02077_ net1214 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[667\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08519__Y _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15798_ net2132 _02008_ net1229 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[598\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07819__A1 net1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14754__924 clknet_leaf_143_clk vssd1 vssd1 vccd1 vccd1 net2393 sky130_fd_sc_hd__inv_2
XFILLER_33_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08270_ top.CPU.registers.data\[694\] top.CPU.registers.data\[662\] net998 vssd1
+ vssd1 vccd1 vccd1 _03909_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16419_ clknet_leaf_55_clk net2625 net1143 vssd1 vssd1 vccd1 vccd1 top.I2C.I2C_state\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10944__C _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08244__A1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13320__C net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12040__A2 _06779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10051__A1 _03148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12932__S net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_8_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_173_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10960__B net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13540__A2 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10305__X _05937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout126 net127 vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10354__A2 _05733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout137 _05771_ vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__buf_2
Xfanout148 _06412_ vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__buf_2
XANTENNA__13828__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout159 _06761_ vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__clkbuf_8
X_07985_ top.CPU.registers.data\[568\] top.CPU.registers.data\[536\] net983 vssd1
+ vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__mux2_1
XFILLER_86_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout384_A net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09724_ _05361_ _05362_ net455 vssd1 vssd1 vccd1 vccd1 _05363_ sky130_fd_sc_hd__mux2_1
XFILLER_86_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11303__B2 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09655_ _05290_ _05292_ _04125_ vssd1 vssd1 vccd1 vccd1 _05294_ sky130_fd_sc_hd__a21o_1
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11854__A2 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout172_X net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout551_A _03172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1293_A _03113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08606_ top.CPU.registers.data\[559\] top.CPU.registers.data\[527\] net974 vssd1
+ vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout649_A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09586_ net619 _05220_ _05224_ _05216_ vssd1 vssd1 vccd1 vccd1 _05225_ sky130_fd_sc_hd__o31a_1
XFILLER_55_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_78 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11067__B1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08537_ net675 _04166_ _04167_ _04175_ net605 vssd1 vssd1 vccd1 vccd1 _04176_ sky130_fd_sc_hd__a311o_1
XANTENNA__15052__Q top.CPU.alu.program_counter\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout437_X net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout816_A net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1179_X net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10814__B1 _05754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11015__C net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08468_ top.CPU.registers.data\[753\] net1383 net988 top.CPU.registers.data\[721\]
+ net913 vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__a221o_1
XANTENNA__08483__B2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14497__667 clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 net2136 sky130_fd_sc_hd__inv_2
XANTENNA__13359__A2 _07089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12016__C1 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08399_ top.CPU.registers.data\[594\] net1292 net1006 top.CPU.registers.data\[626\]
+ net930 vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout604_X net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1346_X net1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10430_ net573 net515 net439 _06057_ vssd1 vssd1 vccd1 vccd1 _06058_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_94_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09432__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10042__A1 top.CPU.alu.immediate\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10361_ net3845 net226 net316 _05991_ vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__a22o_1
XFILLER_136_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12100_ net563 net361 _06633_ net177 top.CPU.registers.data\[102\] vssd1 vssd1 vccd1
+ vccd1 _06818_ sky130_fd_sc_hd__a32o_1
XANTENNA__07994__B1 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13080_ top.CPU.data_out\[15\] net3194 net558 vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__mux2_1
XANTENNA__09717__A net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10292_ _05789_ _05795_ net389 vssd1 vssd1 vccd1 vccd1 _05925_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout973_X net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10870__B _05808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12031_ net139 net3353 net151 vssd1 vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__mux2_1
XANTENNA__08538__A2 net1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold180 top.CPU.fetch.current_ra\[16\] vssd1 vssd1 vccd1 vccd1 net2737 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold191 top.CPU.registers.data\[402\] vssd1 vssd1 vccd1 vccd1 net2748 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07746__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11542__B2 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08943__C1 net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout660 net662 vssd1 vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__buf_4
Xfanout671 _00000_ vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__buf_2
XFILLER_144_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout682 net683 vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__buf_2
XANTENNA__12098__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14906__1076 clknet_leaf_162_clk vssd1 vssd1 vccd1 vccd1 net2545 sky130_fd_sc_hd__inv_2
Xfanout693 net694 vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__buf_2
XANTENNA__12797__B _04189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15721_ net2055 _01931_ net1060 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[521\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12933_ top.CPU.alu.program_counter\[28\] _07374_ net1361 vssd1 vssd1 vccd1 vccd1
+ _01191_ sky130_fd_sc_hd__mux2_1
XANTENNA__11845__A2 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15652_ net1986 _01862_ net1211 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[452\]
+ sky130_fd_sc_hd__dfrtp_1
X_12864_ _07310_ _07311_ vssd1 vssd1 vccd1 vccd1 _07312_ sky130_fd_sc_hd__nor2_1
X_14441__611 clknet_leaf_156_clk vssd1 vssd1 vccd1 vccd1 net2080 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_87_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14738__908 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 net2377 sky130_fd_sc_hd__inv_2
XANTENNA__11058__B1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11815_ net143 net3638 net156 vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__mux2_1
X_12795_ _07249_ _07248_ net128 vssd1 vssd1 vccd1 vccd1 _07250_ sky130_fd_sc_hd__mux2_1
X_15583_ net1917 _01793_ net1222 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[383\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09120__C1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08474__A1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11746_ _06588_ net200 net193 net2730 vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_120_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14834__1004 clknet_leaf_193_clk vssd1 vssd1 vccd1 vccd1 net2473 sky130_fd_sc_hd__inv_2
XFILLER_105_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07700__A _03116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11677_ net465 _06494_ net238 net166 net3040 vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__a32o_1
XFILLER_146_107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16204_ net2538 _02414_ net1069 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[1004\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11222__A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10628_ _05672_ _05873_ _06141_ _05862_ vssd1 vssd1 vccd1 vccd1 _06247_ sky130_fd_sc_hd__a211o_1
X_13416_ top.CPU.control_unit.instruction\[29\] _02929_ net670 vssd1 vssd1 vccd1 vccd1
+ _02463_ sky130_fd_sc_hd__mux2_1
XFILLER_128_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13347_ top.mmio.mem_data_i\[11\] net592 net1343 vssd1 vssd1 vccd1 vccd1 _02879_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__08321__S1 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16135_ net2469 _02345_ net1203 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[935\]
+ sky130_fd_sc_hd__dfrtp_1
X_10559_ _05664_ _05740_ _05760_ _05671_ _06140_ vssd1 vssd1 vccd1 vccd1 _06181_ sky130_fd_sc_hd__o221a_1
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13278_ _07059_ _02824_ _02823_ _07056_ vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_149_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16066_ net2400 _02276_ net1177 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[866\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_149_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10780__B net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13522__A2 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15017_ clknet_leaf_96_clk _01262_ net1247 vssd1 vssd1 vccd1 vccd1 top.SPI.parameters\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13149__A _03118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12229_ _06695_ net245 net170 top.CPU.registers.data\[36\] vssd1 vssd1 vccd1 vccd1
+ _06881_ sky130_fd_sc_hd__a22o_1
XFILLER_97_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_166_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12730__A0 top.CPU.alu.program_counter\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11533__A1 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07770_ top.CPU.control_unit.instruction\[30\] net1046 net899 vssd1 vssd1 vccd1 vccd1
+ _03409_ sky130_fd_sc_hd__o21a_2
XANTENNA__12089__A2 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07581__S net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15919_ net2253 _02129_ net1104 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[719\]
+ sky130_fd_sc_hd__dfrtp_1
X_09440_ net677 _05077_ _05078_ vssd1 vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__and3_1
XANTENNA__08701__A2 net1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10301__A _03167_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14184__354 clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 net1823 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_140_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09371_ net679 _05000_ _05001_ net915 vssd1 vssd1 vccd1 vccd1 _05010_ sky130_fd_sc_hd__o211a_1
XANTENNA__11116__B net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09111__C1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08322_ top.CPU.registers.data\[435\] top.CPU.registers.data\[403\] top.CPU.registers.data\[307\]
+ top.CPU.registers.data\[275\] net988 net913 vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__mux4_1
XFILLER_21_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10955__B _05697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10272__A1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14225__395 clknet_leaf_179_clk vssd1 vssd1 vccd1 vccd1 net1864 sky130_fd_sc_hd__inv_2
XANTENNA__09301__S net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08253_ top.CPU.registers.data\[950\] top.CPU.registers.data\[918\] top.CPU.registers.data\[822\]
+ top.CPU.registers.data\[790\] net993 net917 vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__mux4_1
XFILLER_138_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout132_A _06085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11132__A net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08184_ top.CPU.control_unit.instruction\[23\] net1045 net899 vssd1 vssd1 vccd1 vccd1
+ _03823_ sky130_fd_sc_hd__o21a_2
Xteam_08_1460 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] team_08_1460/LO sky130_fd_sc_hd__conb_1
XFILLER_145_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12662__S net1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10971__A net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1041_A net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13907__77 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 net1546 sky130_fd_sc_hd__inv_2
XFILLER_161_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_560 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10327__A2 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12721__A0 top.CPU.alu.program_counter\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1306_A net1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08925__C1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout766_A net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07968_ net745 _03596_ _03597_ _03606_ vssd1 vssd1 vccd1 vccd1 _03607_ sky130_fd_sc_hd__a31o_1
XFILLER_74_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09707_ top.CPU.registers.data\[601\] net1306 net1029 top.CPU.registers.data\[633\]
+ net946 vssd1 vssd1 vccd1 vccd1 _05346_ sky130_fd_sc_hd__a221o_1
XANTENNA__13506__B _02966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07899_ net800 _03528_ _03529_ net755 vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout933_A net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1296_X net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09638_ _04732_ _04797_ _05276_ vssd1 vssd1 vccd1 vccd1 _05277_ sky130_fd_sc_hd__or3_1
XFILLER_130_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11026__B _06570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09569_ net673 _05202_ _05203_ _05206_ net619 vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__a311o_1
XANTENNA_fanout721_X net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12788__A0 top.CPU.alu.program_counter\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11600_ net136 net3180 net214 vssd1 vssd1 vccd1 vccd1 _01949_ sky130_fd_sc_hd__mux2_1
XANTENNA__09102__C1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12580_ _07062_ _07081_ _07083_ _07084_ vssd1 vssd1 vccd1 vccd1 _00024_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_65_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10799__C1 _06401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10865__B net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11460__A0 _06230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11531_ net3476 net251 _06734_ _06500_ vssd1 vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__a22o_1
XANTENNA__13241__B _02803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11042__A net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11462_ net145 net3819 net264 vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__mux2_1
XFILLER_109_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09405__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13201_ top.I2C.within_byte_counter_reading\[1\] top.I2C.within_byte_counter_reading\[0\]
+ top.I2C.within_byte_counter_reading\[2\] vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__and3b_2
X_10413_ _05942_ _06040_ net392 vssd1 vssd1 vccd1 vccd1 _06041_ sky130_fd_sc_hd__mux2_1
X_11393_ _06515_ net284 net273 net3116 vssd1 vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__a22o_1
XANTENNA__11763__A1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13132_ top.SPI.counter\[0\] net595 _02730_ vssd1 vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__a21o_1
X_10344_ _03613_ _03822_ net374 vssd1 vssd1 vccd1 vccd1 _05975_ sky130_fd_sc_hd__mux2_1
XANTENNA__09447__A net1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09169__C1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13063_ net3280 top.CPU.data_out\[10\] net557 vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__mux2_1
XFILLER_152_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10275_ net3441 net227 net319 _05908_ vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__a22o_1
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08070__B net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1400 top.CPU.control_unit.instruction\[12\] vssd1 vssd1 vccd1 vccd1 net1400
+ sky130_fd_sc_hd__clkbuf_4
X_12014_ net567 _06580_ net364 net151 top.CPU.registers.data\[154\] vssd1 vssd1 vccd1
+ vccd1 _06784_ sky130_fd_sc_hd__a32o_1
Xfanout1411 top.I2C.bit_timer_state\[1\] vssd1 vssd1 vccd1 vccd1 net1411 sky130_fd_sc_hd__clkbuf_2
XFILLER_120_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_109_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13921__91 clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 net1560 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_144_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08931__A2 net1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_6_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout490 net491 vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_161_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_161_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14168__338 clknet_leaf_168_clk vssd1 vssd1 vccd1 vccd1 net1807 sky130_fd_sc_hd__inv_2
XFILLER_0_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09341__C1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15704_ net2038 _01914_ net1148 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[504\]
+ sky130_fd_sc_hd__dfrtp_1
X_12916_ _07356_ _07358_ vssd1 vssd1 vccd1 vccd1 _07359_ sky130_fd_sc_hd__nand2_1
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload8_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_100_Left_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15635_ net1969 _01845_ net1184 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[435\]
+ sky130_fd_sc_hd__dfrtp_1
X_12847_ _07291_ _07295_ vssd1 vssd1 vccd1 vccd1 _07297_ sky130_fd_sc_hd__xnor2_1
X_14209__379 clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 net1848 sky130_fd_sc_hd__inv_2
XFILLER_21_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15566_ net1900 _01776_ net1104 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[366\]
+ sky130_fd_sc_hd__dfrtp_1
X_12778_ _07232_ _07233_ vssd1 vssd1 vccd1 vccd1 _07234_ sky130_fd_sc_hd__nand2_1
XFILLER_14_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11451__A0 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11729_ net138 net539 net500 net194 net2771 vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__a32o_1
XFILLER_119_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15497_ net1831 _01707_ net1061 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[297\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08960__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10006__A1 _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold905 top.CPU.registers.data\[195\] vssd1 vssd1 vccd1 vccd1 net3462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold916 top.SPI.timem\[3\] vssd1 vssd1 vccd1 vccd1 net3473 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_836 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07958__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold927 net98 vssd1 vssd1 vccd1 vccd1 net3484 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16118_ net2452 _02328_ net1228 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[918\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold938 top.CPU.registers.data\[347\] vssd1 vssd1 vccd1 vccd1 net3495 sky130_fd_sc_hd__dlygate4sd3_1
Xhold949 top.CPU.registers.data\[507\] vssd1 vssd1 vccd1 vccd1 net3506 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12054__Y _06796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16251__Q top.CPU.control_unit.instruction\[27\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_171_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08940_ net951 _04575_ _04578_ net626 vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__a211o_1
X_16049_ net2383 _02259_ net1175 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[849\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09791__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08907__C1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12164__D1 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14610__780 clknet_leaf_201_clk vssd1 vssd1 vccd1 vccd1 net2249 sky130_fd_sc_hd__inv_2
X_08871_ top.CPU.registers.data\[235\] net1386 net807 top.CPU.registers.data\[203\]
+ net762 vssd1 vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__a221o_1
XANTENNA__10015__B net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07822_ top.CPU.registers.data\[61\] top.CPU.registers.data\[29\] net817 vssd1 vssd1
+ vccd1 vccd1 _03461_ sky130_fd_sc_hd__mux2_1
XANTENNA__13259__A1 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12511__A _04222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09092__A _04698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07753_ net800 _03391_ vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__or2_1
XANTENNA__08135__B1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09332__C1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07684_ _03270_ _03283_ vssd1 vssd1 vccd1 vccd1 _03323_ sky130_fd_sc_hd__nor2_2
XFILLER_25_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09423_ top.CPU.registers.data\[674\] top.CPU.registers.data\[642\] top.CPU.registers.data\[546\]
+ top.CPU.registers.data\[514\] net986 net911 vssd1 vssd1 vccd1 vccd1 _05062_ sky130_fd_sc_hd__mux4_1
XANTENNA__10493__A1 _04123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12561__A_N _06147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11690__B1 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07894__C1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout347_A net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09354_ top.CPU.registers.data\[387\] net1297 net1018 top.CPU.registers.data\[419\]
+ net915 vssd1 vssd1 vccd1 vccd1 _04993_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1089_A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12234__A2 _06770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08305_ top.CPU.registers.data\[851\] net1324 net855 top.CPU.registers.data\[883\]
+ net748 vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__a221o_1
XFILLER_21_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09285_ top.CPU.registers.data\[292\] top.CPU.registers.data\[260\] net992 vssd1
+ vssd1 vccd1 vccd1 _04924_ sky130_fd_sc_hd__mux2_1
XFILLER_21_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout514_A net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08236_ top.CPU.registers.data\[854\] net1330 net861 top.CPU.registers.data\[886\]
+ net753 vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_60_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13488__S net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14905__1075 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 net2544 sky130_fd_sc_hd__inv_2
X_08167_ top.CPU.registers.data\[759\] net1391 net824 top.CPU.registers.data\[727\]
+ net723 vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__a221o_1
XFILLER_4_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout302_X net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07949__B1 net1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_6 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08098_ net798 _03735_ _03736_ net726 vssd1 vssd1 vccd1 vccd1 _03737_ sky130_fd_sc_hd__o211a_1
XFILLER_134_666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13498__A1 _03369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1309_X net1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10060_ _05509_ _05513_ _05511_ _03445_ vssd1 vssd1 vccd1 vccd1 _05698_ sky130_fd_sc_hd__o211ai_1
XFILLER_121_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout671_X net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14833__1003 clknet_leaf_188_clk vssd1 vssd1 vccd1 vccd1 net2472 sky130_fd_sc_hd__inv_2
XANTENNA__08374__B1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout769_X net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13517__A _04122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout936_X net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09323__C1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11037__A _05808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13750_ top.SPI.timem\[22\] _03085_ vssd1 vssd1 vccd1 vccd1 _03086_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_67_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10962_ _05906_ net545 vssd1 vssd1 vccd1 vccd1 _06532_ sky130_fd_sc_hd__nand2_1
XFILLER_28_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12701_ top.CPU.alu.program_counter\[7\] top.CPU.alu.program_counter\[6\] _07152_
+ vssd1 vssd1 vccd1 vccd1 _07164_ sky130_fd_sc_hd__and3_1
XANTENNA__11681__B1 net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13681_ net2645 net336 vssd1 vssd1 vccd1 vccd1 _02609_ sky130_fd_sc_hd__and2_1
XANTENNA__10876__A net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10893_ net489 _06035_ net437 vssd1 vssd1 vccd1 vccd1 _06490_ sky130_fd_sc_hd__and3_1
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15420_ net1754 _01630_ net1196 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[220\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12632_ net1411 net1341 net2741 vssd1 vssd1 vccd1 vccd1 _00015_ sky130_fd_sc_hd__and3_1
XANTENNA__12225__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13422__B2 _07088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12563_ _06067_ _06081_ _07067_ vssd1 vssd1 vccd1 vccd1 _07068_ sky130_fd_sc_hd__and3_1
XANTENNA__10087__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15351_ net1685 _01561_ net1182 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[151\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11433__B1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11514_ top.CPU.registers.data\[605\] net250 vssd1 vssd1 vccd1 vccd1 _06735_ sky130_fd_sc_hd__and2_1
XFILLER_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12494_ _04952_ _04986_ _05019_ _05054_ vssd1 vssd1 vccd1 vccd1 _07003_ sky130_fd_sc_hd__a22o_1
X_15282_ net1616 _01492_ net1100 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[82\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_22_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14553__723 clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 net2192 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_22_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11445_ net3452 net266 _06722_ net496 vssd1 vssd1 vccd1 vccd1 _02072_ sky130_fd_sc_hd__a22o_1
XFILLER_172_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_931 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08601__A1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08062__C1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11376_ _06491_ net278 net272 net3324 vssd1 vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__a22o_1
XFILLER_4_952 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_156_Right_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13115_ net2729 _02722_ net897 vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__mux2_1
X_10327_ top.CPU.fetch.current_ra\[24\] net1042 net883 top.CPU.handler.toreg\[24\]
+ vssd1 vssd1 vccd1 vccd1 _05959_ sky130_fd_sc_hd__a22o_1
XANTENNA__10116__A net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13489__A1 _05018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_163_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13898__68 clknet_leaf_147_clk vssd1 vssd1 vccd1 vccd1 net1537 sky130_fd_sc_hd__inv_2
X_13046_ net2890 _07448_ net895 vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__mux2_1
XANTENNA__09905__A net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10258_ _05889_ _05891_ net399 vssd1 vssd1 vccd1 vccd1 _05892_ sky130_fd_sc_hd__mux2_2
Xfanout1230 net1232 vssd1 vssd1 vccd1 vccd1 net1230 sky130_fd_sc_hd__clkbuf_4
Xfanout1241 net1242 vssd1 vssd1 vccd1 vccd1 net1241 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09562__C1 net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10189_ _03476_ _03544_ net375 vssd1 vssd1 vccd1 vccd1 _05825_ sky130_fd_sc_hd__mux2_1
Xfanout1252 net1259 vssd1 vssd1 vccd1 vccd1 net1252 sky130_fd_sc_hd__clkbuf_4
Xfanout1263 net1266 vssd1 vssd1 vccd1 vccd1 net1263 sky130_fd_sc_hd__clkbuf_4
Xfanout1274 net1275 vssd1 vssd1 vccd1 vccd1 net1274 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09116__S net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1285 _03114_ vssd1 vssd1 vccd1 vccd1 net1285 sky130_fd_sc_hd__buf_4
XANTENNA__13146__B top.CPU.alu.program_counter\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1296 net1301 vssd1 vssd1 vccd1 vccd1 net1296 sky130_fd_sc_hd__clkbuf_4
X_14997_ clknet_leaf_94_clk _01242_ net1260 vssd1 vssd1 vccd1 vccd1 top.SPI.parameters\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08117__B1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08955__S net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12464__A2 _05361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11672__B1 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07876__C1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15618_ net1952 _01828_ net1172 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[418\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09617__B1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11424__B1 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15549_ net1883 _01759_ net1114 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[349\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_174_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09070_ top.CPU.registers.data\[200\] net1373 net969 top.CPU.registers.data\[232\]
+ net927 vssd1 vssd1 vccd1 vccd1 _04709_ sky130_fd_sc_hd__o221a_1
XFILLER_163_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14296__466 clknet_leaf_174_clk vssd1 vssd1 vccd1 vccd1 net1935 sky130_fd_sc_hd__inv_2
X_08021_ net791 _03654_ _03655_ net719 vssd1 vssd1 vccd1 vccd1 _03660_ sky130_fd_sc_hd__o211a_1
XFILLER_162_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold702 top.CPU.fetch.current_ra\[21\] vssd1 vssd1 vccd1 vccd1 net3259 sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 top.mmio.mem_data_i\[29\] vssd1 vssd1 vccd1 vccd1 net3270 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold724 top.CPU.registers.data\[715\] vssd1 vssd1 vccd1 vccd1 net3281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold735 top.CPU.registers.data\[779\] vssd1 vssd1 vccd1 vccd1 net3292 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_1032 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold746 top.CPU.registers.data\[926\] vssd1 vssd1 vccd1 vccd1 net3303 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold757 top.CPU.registers.data\[870\] vssd1 vssd1 vccd1 vccd1 net3314 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold768 top.CPU.registers.data\[731\] vssd1 vssd1 vccd1 vccd1 net3325 sky130_fd_sc_hd__dlygate4sd3_1
X_09972_ _05602_ _05603_ _03580_ vssd1 vssd1 vccd1 vccd1 _05611_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_123_Right_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold779 top.CPU.registers.data\[516\] vssd1 vssd1 vccd1 vccd1 net3336 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09148__A2 net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08923_ top.CPU.registers.data\[938\] top.CPU.registers.data\[906\] net809 vssd1
+ vssd1 vccd1 vccd1 _04562_ sky130_fd_sc_hd__mux2_1
XFILLER_58_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout297_A _06645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1402 top.mmio.mem_data_i\[15\] vssd1 vssd1 vccd1 vccd1 net3959 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1413 top.CPU.addressnew\[12\] vssd1 vssd1 vccd1 vccd1 net3970 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08854_ top.CPU.registers.data\[459\] net1369 net967 top.CPU.registers.data\[491\]
+ net1364 vssd1 vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__o221a_1
Xhold1424 top.CPU.handler.toreg\[15\] vssd1 vssd1 vccd1 vccd1 net3981 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1004_A net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10702__A2 _05979_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1435 top.I2C.bit_timer_counter\[1\] vssd1 vssd1 vccd1 vccd1 net3992 sky130_fd_sc_hd__dlygate4sd3_1
X_07805_ _03442_ _03443_ vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__and2_1
Xhold1446 top.CPU.registers.data\[85\] vssd1 vssd1 vccd1 vccd1 net4003 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1457 top.SPI.timem\[14\] vssd1 vssd1 vccd1 vccd1 net4014 sky130_fd_sc_hd__dlygate4sd3_1
X_08785_ net789 _04414_ _04415_ net742 vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__o211a_1
Xhold1468 top.SPI.register\[0\] vssd1 vssd1 vccd1 vccd1 net4025 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10032__Y _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout464_A net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07736_ _03374_ vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__inv_2
XFILLER_44_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12455__A2 _03508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09856__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12895__B _05362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10466__A1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07667_ _03298_ _03305_ vssd1 vssd1 vccd1 vccd1 _03306_ sky130_fd_sc_hd__nor2_2
XANTENNA__11663__B1 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10696__A net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout252_X net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1373_A net1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout729_A net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09406_ net708 _05043_ _05044_ _05042_ vssd1 vssd1 vccd1 vccd1 _05045_ sky130_fd_sc_hd__a31o_1
XFILLER_125_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07598_ top.CPU.registers.data\[223\] net1392 net836 top.CPU.registers.data\[255\]
+ net756 vssd1 vssd1 vccd1 vccd1 _03237_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_62_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12207__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14240__410 clknet_leaf_125_clk vssd1 vssd1 vccd1 vccd1 net1879 sky130_fd_sc_hd__inv_2
XANTENNA__10218__B2 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11415__B1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09337_ top.CPU.registers.data\[740\] net1391 net829 top.CPU.registers.data\[708\]
+ net726 vssd1 vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__a221o_1
X_14537__707 clknet_leaf_156_clk vssd1 vssd1 vccd1 vccd1 net2176 sky130_fd_sc_hd__inv_2
XANTENNA_fanout517_X net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1259_X net1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09696__S net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09268_ net676 _04905_ _04906_ vssd1 vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__and3_1
XANTENNA__08453__X _04092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11023__C net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08292__C1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08219_ _03822_ _03855_ vssd1 vssd1 vccd1 vccd1 _03858_ sky130_fd_sc_hd__or2_1
XFILLER_126_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09199_ net930 _04833_ _04834_ net618 vssd1 vssd1 vccd1 vccd1 _04838_ sky130_fd_sc_hd__o211a_1
XFILLER_5_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11230_ net527 _05962_ net544 vssd1 vssd1 vccd1 vccd1 _06670_ sky130_fd_sc_hd__and3_1
XFILLER_135_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09387__A2 net1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11161_ net1405 net576 net525 net131 vssd1 vssd1 vccd1 vccd1 _06641_ sky130_fd_sc_hd__and4_1
XFILLER_136_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12128__D1 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10112_ _03544_ _05399_ net379 vssd1 vssd1 vccd1 vccd1 _05750_ sky130_fd_sc_hd__mux2_1
XANTENNA__09139__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11092_ net486 _06599_ vssd1 vssd1 vccd1 vccd1 _06603_ sky130_fd_sc_hd__nor2_2
XFILLER_121_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11466__S net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10043_ _03315_ _03375_ net410 _05668_ _05681_ vssd1 vssd1 vccd1 vccd1 _05682_ sky130_fd_sc_hd__a221o_1
X_14920_ clknet_leaf_28_clk _01166_ net1149 vssd1 vssd1 vccd1 vccd1 top.CPU.alu.program_counter\[3\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold40 top.CPU.registers.data_out_r2_prev\[3\] vssd1 vssd1 vccd1 vccd1 net2597 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 top.I2C.I2C_state\[13\] vssd1 vssd1 vccd1 vccd1 net2608 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold62 top.CPU.registers.data_out_r1_prev\[31\] vssd1 vssd1 vccd1 vccd1 net2619 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input25_A DAT_I[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold73 top.SPI.timem\[23\] vssd1 vssd1 vccd1 vccd1 net2630 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10159__A2_N net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold84 top.CPU.registers.data\[817\] vssd1 vssd1 vccd1 vccd1 net2641 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1032 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold95 top.CPU.registers.data\[295\] vssd1 vssd1 vccd1 vccd1 net2652 sky130_fd_sc_hd__dlygate4sd3_1
X_13802_ net3815 net333 net326 top.CPU.data_out\[4\] vssd1 vssd1 vccd1 vccd1 _02682_
+ sky130_fd_sc_hd__a22o_1
XFILLER_75_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08775__S net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11994_ _06559_ net342 net180 net2793 vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__a22o_1
X_16521_ clknet_leaf_100_clk _02683_ net1255 vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__dfrtp_1
X_13733_ net3786 _03075_ vssd1 vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__xnor2_1
XFILLER_16_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11654__B1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07858__C1 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10945_ net3580 net223 _06521_ net319 vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__a22o_1
XFILLER_17_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16452_ clknet_leaf_85_clk _02615_ net1242 vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_27_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13664_ _07092_ _07091_ vssd1 vssd1 vccd1 vccd1 _03046_ sky130_fd_sc_hd__and2b_1
X_10876_ net661 _05906_ vssd1 vssd1 vccd1 vccd1 _06478_ sky130_fd_sc_hd__and2_1
X_15403_ net1737 _01613_ net1057 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[203\]
+ sky130_fd_sc_hd__dfrtp_1
X_12615_ _03127_ top.SPI.state\[5\] _07114_ vssd1 vssd1 vccd1 vccd1 _00073_ sky130_fd_sc_hd__a21o_1
XANTENNA__11406__B1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16383_ clknet_leaf_25_clk _02592_ net1155 vssd1 vssd1 vccd1 vccd1 top.CPU.fetch.current_ra\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_156_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13595_ top.CPU.addressnew\[18\] net578 _03022_ _03023_ vssd1 vssd1 vccd1 vccd1 _02548_
+ sky130_fd_sc_hd__a22o_1
XFILLER_169_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15334_ net1668 _01544_ net1081 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[134\]
+ sky130_fd_sc_hd__dfrtp_1
X_12546_ _03133_ top.mmio.m2 top.mmio.m1 top.mmio.s2 _03134_ vssd1 vssd1 vccd1 vccd1
+ _07055_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_117_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14024__194 clknet_leaf_130_clk vssd1 vssd1 vccd1 vccd1 net1663 sky130_fd_sc_hd__inv_2
X_15265_ net1599 _01475_ net1232 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[65\]
+ sky130_fd_sc_hd__dfrtp_1
X_12477_ net451 _03717_ _03955_ _03984_ vssd1 vssd1 vccd1 vccd1 _06986_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_4 net4000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11230__A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08035__C1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08015__S net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11428_ _06571_ net282 net270 net3132 vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__a22o_1
XFILLER_126_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15196_ net1533 _01406_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r1_prev\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11185__A2 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09783__C1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11359_ net3602 net287 net284 _06413_ vssd1 vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__a22o_1
XFILLER_4_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08050__A2 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13029_ top.SPI.parameters\[16\] top.SPI.paroutput\[8\] net1357 vssd1 vssd1 vccd1
+ vccd1 _07440_ sky130_fd_sc_hd__mux2_1
XFILLER_112_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10133__X _05771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08889__A1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1060 net1068 vssd1 vssd1 vccd1 vccd1 net1060 sky130_fd_sc_hd__clkbuf_4
Xfanout1071 net1075 vssd1 vssd1 vccd1 vccd1 net1071 sky130_fd_sc_hd__clkbuf_4
X_14681__851 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 net2320 sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_6_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11893__A0 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1082 net1111 vssd1 vssd1 vccd1 vccd1 net1082 sky130_fd_sc_hd__buf_2
Xfanout1093 net1110 vssd1 vssd1 vccd1 vccd1 net1093 sky130_fd_sc_hd__clkbuf_2
X_14904__1074 clknet_leaf_160_clk vssd1 vssd1 vccd1 vccd1 net2543 sky130_fd_sc_hd__inv_2
X_08570_ top.CPU.registers.data\[847\] net1315 net845 top.CPU.registers.data\[879\]
+ net740 vssd1 vssd1 vccd1 vccd1 _04209_ sky130_fd_sc_hd__a221o_1
XANTENNA__10448__A1 _03986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07521_ net1045 _03159_ vssd1 vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__and2_4
XANTENNA__11645__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14722__892 clknet_leaf_140_clk vssd1 vssd1 vccd1 vccd1 net2361 sky130_fd_sc_hd__inv_2
XANTENNA__08510__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07864__A2 net1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13398__B1 net1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14832__1002 clknet_leaf_196_clk vssd1 vssd1 vccd1 vccd1 net2471 sky130_fd_sc_hd__inv_2
X_09122_ _04757_ _04760_ net1308 vssd1 vssd1 vccd1 vccd1 _04761_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_40_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08274__C1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09053_ net785 _04682_ _04691_ net739 vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout212_A _06752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11140__A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08004_ net952 _03637_ _03639_ _03642_ vssd1 vssd1 vccd1 vccd1 _03643_ sky130_fd_sc_hd__a31o_1
Xhold510 top.CPU.registers.data\[280\] vssd1 vssd1 vccd1 vccd1 net3067 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold521 top.CPU.registers.data\[143\] vssd1 vssd1 vccd1 vccd1 net3078 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08577__B1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold532 top.CPU.registers.data\[405\] vssd1 vssd1 vccd1 vccd1 net3089 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11176__A2 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09774__C1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold543 top.CPU.registers.data\[857\] vssd1 vssd1 vccd1 vccd1 net3100 sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 _02704_ vssd1 vssd1 vccd1 vccd1 net3111 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12670__S net1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold565 top.CPU.registers.data\[359\] vssd1 vssd1 vccd1 vccd1 net3122 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold576 net62 vssd1 vssd1 vccd1 vccd1 net3133 sky130_fd_sc_hd__dlygate4sd3_1
Xhold587 top.CPU.registers.data\[977\] vssd1 vssd1 vccd1 vccd1 net3144 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1219_A net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold598 net96 vssd1 vssd1 vccd1 vccd1 net3155 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11794__B net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09545__A net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09955_ _05575_ _05580_ _05592_ _05593_ vssd1 vssd1 vccd1 vccd1 _05594_ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_38_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08329__B1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout679_A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08906_ net787 _04544_ vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_55_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09264__B net1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09886_ _05524_ vssd1 vssd1 vccd1 vccd1 _05525_ sky130_fd_sc_hd__inv_2
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1210 top.CPU.registers.data\[583\] vssd1 vssd1 vccd1 vccd1 net3767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1221 top.CPU.registers.data\[153\] vssd1 vssd1 vccd1 vccd1 net3778 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1232 top.CPU.registers.data\[930\] vssd1 vssd1 vccd1 vccd1 net3789 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11884__A0 _06212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09541__A2 net1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08837_ _04474_ _04475_ net672 vssd1 vssd1 vccd1 vccd1 _04476_ sky130_fd_sc_hd__o21a_1
Xhold1243 top.CPU.registers.data\[861\] vssd1 vssd1 vccd1 vccd1 net3800 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1254 net70 vssd1 vssd1 vccd1 vccd1 net3811 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout846_A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout467_X net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1265 top.CPU.registers.data\[340\] vssd1 vssd1 vccd1 vccd1 net3822 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09551__Y _05190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1276 top.CPU.registers.data\[1004\] vssd1 vssd1 vccd1 vccd1 net3833 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1287 top.SPI.timem\[4\] vssd1 vssd1 vccd1 vccd1 net3844 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1298 top.CPU.fetch.current_ra\[5\] vssd1 vssd1 vccd1 vccd1 net3855 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09829__B1 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08595__S net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08768_ net746 _04405_ _04406_ net767 vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__o211a_1
XFILLER_82_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08727__S1 net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07719_ top.CPU.registers.data\[511\] top.CPU.registers.data\[479\] top.CPU.registers.data\[447\]
+ top.CPU.registers.data\[415\] net999 net959 vssd1 vssd1 vccd1 vccd1 _03358_ sky130_fd_sc_hd__mux4_1
XANTENNA__11636__B1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout634_X net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08699_ top.CPU.registers.data\[749\] net1386 net807 top.CPU.registers.data\[717\]
+ net714 vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1376_X net1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08501__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10857__C net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10730_ _06262_ _06343_ net388 vssd1 vssd1 vccd1 vccd1 _06344_ sky130_fd_sc_hd__mux2_1
XFILLER_25_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10661_ _04567_ _04634_ net373 vssd1 vssd1 vccd1 vccd1 _06278_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout801_X net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12400_ _03121_ net2627 top.I2C.I2C_state\[22\] vssd1 vssd1 vccd1 vccd1 _00036_ sky130_fd_sc_hd__a21o_1
XANTENNA__09279__X _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13380_ top.CPU.control_unit.instruction\[19\] _02903_ net667 vssd1 vssd1 vccd1 vccd1
+ _02453_ sky130_fd_sc_hd__mux2_1
X_14008__178 clknet_leaf_167_clk vssd1 vssd1 vccd1 vccd1 net1647 sky130_fd_sc_hd__inv_2
XANTENNA__08265__C1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_864 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10592_ net660 net438 _06212_ vssd1 vssd1 vccd1 vccd1 _06213_ sky130_fd_sc_hd__and3_2
XFILLER_12_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12331_ net3124 _04659_ net1234 vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__mux2_1
XFILLER_127_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10592__C _06212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15050_ clknet_leaf_92_clk _01295_ net1269 vssd1 vssd1 vccd1 vccd1 top.SPI.command\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_12262_ net2758 net144 net431 vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__mux2_1
XFILLER_119_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08568__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11213_ net495 _06520_ _06648_ net300 net2953 vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_112_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09765__C1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12193_ net3898 net170 _06863_ _06741_ vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_75_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput41 net41 vssd1 vssd1 vccd1 vccd1 ADR_O[11] sky130_fd_sc_hd__buf_2
Xoutput52 net52 vssd1 vssd1 vccd1 vccd1 ADR_O[21] sky130_fd_sc_hd__buf_2
XANTENNA__10914__A2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11144_ net479 net458 _06631_ net301 net3057 vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__a32o_1
Xoutput63 net63 vssd1 vssd1 vccd1 vccd1 ADR_O[6] sky130_fd_sc_hd__buf_2
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 DAT_O[15] sky130_fd_sc_hd__buf_2
Xoutput85 net85 vssd1 vssd1 vccd1 vccd1 DAT_O[25] sky130_fd_sc_hd__buf_2
XFILLER_122_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13868__38 clknet_leaf_194_clk vssd1 vssd1 vccd1 vccd1 net1507 sky130_fd_sc_hd__inv_2
XANTENNA__12116__A1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput96 net96 vssd1 vssd1 vccd1 vccd1 DAT_O[6] sky130_fd_sc_hd__buf_2
XFILLER_122_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14665__835 clknet_leaf_155_clk vssd1 vssd1 vccd1 vccd1 net2304 sky130_fd_sc_hd__inv_2
XANTENNA__11196__S net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11075_ _06354_ net536 vssd1 vssd1 vccd1 vccd1 _06593_ sky130_fd_sc_hd__and2_1
X_15952_ net2286 _02162_ net1154 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[752\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_163_84 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10026_ _03286_ _03292_ _03321_ vssd1 vssd1 vccd1 vccd1 _05665_ sky130_fd_sc_hd__o21ai_4
XANTENNA__10678__A1 _04634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11875__B1 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09532__A2 net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15883_ net2217 _02093_ net1065 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[683\]
+ sky130_fd_sc_hd__dfrtp_1
X_14706__876 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 net2345 sky130_fd_sc_hd__inv_2
XFILLER_45_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07703__A top.CPU.control_unit.instruction\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11977_ _06534_ net352 net183 net3075 vssd1 vssd1 vccd1 vccd1 _01595_ sky130_fd_sc_hd__a22o_1
X_16504_ clknet_leaf_49_clk _02666_ net1128 vssd1 vssd1 vccd1 vccd1 top.mmio.mem_data_i\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13716_ _03064_ vssd1 vssd1 vccd1 vccd1 _03065_ sky130_fd_sc_hd__inv_2
X_10928_ net487 net518 _06510_ vssd1 vssd1 vccd1 vccd1 _06511_ sky130_fd_sc_hd__and3_1
XFILLER_44_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16435_ clknet_leaf_67_clk net2829 net1168 vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_154_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13647_ top.CPU.fetch.current_ra\[19\] _07289_ net663 vssd1 vssd1 vccd1 vccd1 _02581_
+ sky130_fd_sc_hd__mux2_1
X_10859_ _03170_ _03180_ vssd1 vssd1 vccd1 vccd1 _06466_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_171_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09189__X _04828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07849__S net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16366_ clknet_leaf_60_clk _02575_ net1138 vssd1 vssd1 vccd1 vccd1 top.CPU.fetch.current_ra\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08256__C1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13578_ top.CPU.addressnew\[11\] net578 _03012_ _03013_ vssd1 vssd1 vccd1 vccd1 _02541_
+ sky130_fd_sc_hd__a22o_1
XFILLER_12_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08534__A net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10602__A1 _05667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15317_ net1651 _01527_ net1217 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[117\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10602__B2 _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12529_ _06997_ _07013_ _07033_ _07037_ vssd1 vssd1 vccd1 vccd1 _07038_ sky130_fd_sc_hd__or4b_1
XFILLER_8_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16297_ clknet_leaf_107_clk _02506_ net1248 vssd1 vssd1 vccd1 vccd1 top.CPU.data_out\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_132_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15248_ net1582 _01458_ net1234 vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_172_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11158__A2 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15179_ net1516 _01389_ vssd1 vssd1 vccd1 vccd1 top.CPU.registers.data_out_r1_prev\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_169_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout308 net310 vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09771__A2 net1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout319 net320 vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12503__B _04855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09508__C1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09740_ net799 _05377_ _05378_ net727 vssd1 vssd1 vccd1 vccd1 _05379_ sky130_fd_sc_hd__o211a_1
XANTENNA__10304__A _03650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
.ends

