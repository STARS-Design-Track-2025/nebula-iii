module t07_display(
    input logic clk, nrst, ack,
    output logic [31:0] out
    //output logic delay 
);

    logic [17:0] counter, next_ctr;

    always_ff @(posedge clk, negedge nrst) begin 
        if (~nrst) begin
            counter <= 18'b111111111111111111;
        end else begin
            counter <= next_ctr;
        end
    end

  always_comb begin
    if (ack == 0) begin
        next_ctr = counter + 1;
    end else begin
        next_ctr = counter;
    end

    case (counter) 
        18'd0: out = {16'd3, 16'h80_00}; 
        18'd1: out = {16'd3, 16'h40_00};
        18'd2: out = {16'd3, 16'h80_88};
        18'd3: out = {16'd130, 16'h00_0B};

        18'd4: out = {16'd3, 16'h80_89};
        18'd5: out = {16'd130, 16'h00_02};

        18'd6: out = {16'd3, 16'h80_10};
        18'd7: out = {16'd3, 16'h00_0C};
        18'd8: out = {16'd3, 16'h80_04};
        18'd9: out = {16'd130, 16'h00_81};

        18'd10: out = {16'd3, 16'h80_14};
        18'd11: out = {16'd3, 16'h00_63};
        18'd12: out = {16'd3, 16'h80_15};
        18'd13: out = {16'd3, 16'h00_00};
        18'd14: out = {16'd3, 16'h80_16};
        18'd15: out = {16'd3, 16'h00_03};
        18'd16: out = {16'd3, 16'h80_17};
        18'd17: out = {16'd3, 16'h00_03};
        18'd18: out = {16'd3, 16'h80_18};
        18'd19: out = {16'd3, 16'h00_0B};
        18'd20: out = {16'd3, 16'h80_19};
        18'd21: out = {16'd3, 16'h00_DF};
        18'd22: out = {16'd3, 16'h80_1A};
        18'd23: out = {16'd3, 16'h00_01};
        18'd24: out = {16'd3, 16'h80_1B};
        18'd25: out = {16'd3, 16'h00_1F};
        18'd26: out = {16'd3, 16'h80_1C};
        18'd27: out = {16'd3, 16'h00_00};
        18'd28: out = {16'd3, 16'h80_1D};
        18'd29: out = {16'd3, 16'h00_16};
        18'd30: out = {16'd3, 16'h80_1E};
        18'd31: out = {16'd3, 16'h00_00};
        18'd32: out = {16'd3, 16'h80_1F};
        18'd33: out = {16'd3, 16'h00_01};
        18'd34: out = {16'd3, 16'h80_30};
        18'd35: out = {16'd3, 16'h00_00};
        18'd36: out = {16'd3, 16'h80_31};
        18'd37: out = {16'd3, 16'h00_00};
        18'd38: out = {16'd3, 16'h80_34};
        18'd39: out = {16'd3, 16'h00_1F};
        18'd40: out = {16'd3, 16'h80_35};
        18'd41: out = {16'd3, 16'h00_03};
        18'd42: out = {16'd3, 16'h80_32};
        18'd43: out = {16'd3, 16'h00_00};
        18'd44: out = {16'd3, 16'h80_33};
        18'd45: out = {16'd3, 16'h00_00};
        18'd46: out = {16'd3, 16'h80_36};
        18'd47: out = {16'd3, 16'h00_DF};
        18'd48: out = {16'd3, 16'h80_37};
        18'd49: out = {16'd3, 16'h00_01};
        18'd50: out = {16'd3, 16'h80_8E};
        18'd51: out = {16'd62500, 16'h00_80};


        18'd52: out = {16'd3, 16'h80_01};
        18'd53: out = {16'd3, 16'h00_80};
        18'd54: out = {16'd3, 16'h80_C7};
        18'd55: out = {16'd3, 16'h00_01};
        18'd56: out = {16'd3, 16'h80_8A};
        18'd57: out = {16'd3, 16'h00_8A};
        18'd58: out = {16'd3, 16'h80_8B};
        18'd59: out = {16'd3, 16'h00_80};
        18'd60: out = {16'd3, 16'h80_91};
        18'd61: out = {16'd3, 16'h00_00};
        18'd62: out = {16'd3, 16'h80_92};
        18'd63: out = {16'd3, 16'h00_00};
        18'd64: out = {16'd3, 16'h80_93};
        18'd65: out = {16'd3, 16'h00_00};
        18'd66: out = {16'd3, 16'h80_94};
        18'd67: out = {16'd3, 16'h00_00};
        18'd68: out = {16'd3, 16'h80_95};
        18'd69: out = {16'd3, 16'h00_1F};
        18'd70: out = {16'd3, 16'h80_96};
        18'd71: out = {16'd3, 16'h00_03};
        18'd72: out = {16'd3, 16'h80_97};
        18'd73: out = {16'd3, 16'h00_DF};
        18'd74: out = {16'd3, 16'h80_98};
        18'd75: out = {16'd3, 16'h00_01};
        
        18'd76: out = {16'd3, 16'h80_63};
        18'd77: out = {16'd3, 16'h00_00};
        18'd78: out = {16'd3, 16'h80_64};
        18'd79: out = {16'd3, 16'h00_00};
        18'd80: out = {16'd3, 16'h80_65};
        18'd81: out = {16'd3, 16'h00_00};
        18'd82: out = {16'd3, 16'h80_90};
        18'd83: out = {16'd3, 16'h00_B0};
        18'd84: out = {16'd3, 16'h80_90};
        18'd85: out = {16'd3, 16'h40_00};
        18'd86: out = {16'd3, 16'h80_90};
        18'd87: out = {16'd3, 16'h40_00};
        18'd88: out = {16'd3, 16'h80_90};
        18'd89: out = {16'd3, 16'h40_00};
        18'd90: out = {16'd3, 16'h80_90};
        18'd91: out = {16'd3, 16'h40_00};
        18'd92: out = {16'd3, 16'h80_90};
        18'd93: out = {16'd3, 16'h40_00};
        18'd94: out = {16'd3, 16'h80_90};
        18'd95: out = {16'd3, 16'h40_00};
        18'd96: out = {16'd3, 16'h80_90};
        18'd97: out = {16'd3, 16'h40_00};
        18'd98: out = {16'd3, 16'h80_90};
        18'd99: out = {16'd3, 16'h40_00};
        18'd100: out = {16'd3, 16'h80_90};
        18'd101: out = {16'd3, 16'h40_00};
        18'd102: out = {16'd3, 16'h80_90};
        18'd103: out = {16'd3, 16'h40_00};
        18'd104: out = {16'd3, 16'h80_90};
        18'd105: out = {16'd3, 16'h40_00};
        18'd106: out = {16'd3, 16'h80_90};
        18'd107: out = {16'd3, 16'h40_00};
        18'd108: out = {16'd3, 16'h80_90};
        18'd109: out = {16'd3, 16'h40_00};
        18'd110: out = {16'd3, 16'h80_90};
        18'd111: out = {16'd3, 16'h40_00};
        18'd112: out = {16'd3, 16'h80_90};
        18'd113: out = {16'd3, 16'h40_00};
        18'd114: out = {16'd3, 16'h80_90};
        18'd115: out = {16'd3, 16'h40_00};
        18'd116: out = {16'd3, 16'h80_90};
        18'd117: out = {16'd3, 16'h40_00};
        18'd118: out = {16'd3, 16'h80_90};
        18'd119: out = {16'd3, 16'h40_00};
        18'd120: out = {16'd3, 16'h80_90};
        18'd121: out = {16'd3, 16'h40_00};
        18'd122: out = {16'd3, 16'h80_90};
        18'd123: out = {16'd3, 16'h40_00};
        18'd124: out = {16'd3, 16'h80_90};
        18'd125: out = {16'd3, 16'h40_00};
        18'd126: out = {16'd3, 16'h80_90};
        18'd127: out = {16'd3, 16'h40_00};
        18'd128: out = {16'd3, 16'h80_90};
        18'd129: out = {16'd3, 16'h40_00};
        18'd130: out = {16'd3, 16'h80_90};
        18'd131: out = {16'd3, 16'h40_00};
        18'd132: out = {16'd3, 16'h80_90};
        18'd133: out = {16'd3, 16'h40_00};
        18'd134: out = {16'd3, 16'h80_90};
        18'd135: out = {16'd3, 16'h40_00};
        18'd136: out = {16'd3, 16'h80_90};
        18'd137: out = {16'd3, 16'h40_00};
        18'd138: out = {16'd3, 16'h80_90};
        18'd139: out = {16'd3, 16'h40_00};
        18'd140: out = {16'd3, 16'h80_90};
        18'd141: out = {16'd3, 16'h40_00};
        18'd142: out = {16'd3, 16'h80_90};
        18'd143: out = {16'd3, 16'h40_00};
        18'd144: out = {16'd3, 16'h80_90};
        18'd145: out = {16'd3, 16'h40_00};
        18'd146: out = {16'd3, 16'h80_90};
        18'd147: out = {16'd3, 16'h40_00};
        18'd148: out = {16'd3, 16'h80_90};
        18'd149: out = {16'd3, 16'h40_00};
        18'd150: out = {16'd3, 16'h80_90};
        18'd151: out = {16'd3, 16'h40_00};
        18'd152: out = {16'd3, 16'h80_90};
        18'd153: out = {16'd3, 16'h40_00};
        18'd154: out = {16'd3, 16'h80_90};
        18'd155: out = {16'd3, 16'h40_00};
        18'd156: out = {16'd3, 16'h80_90};
        18'd157: out = {16'd3, 16'h40_00};
        18'd158: out = {16'd3, 16'h80_90};
        18'd159: out = {16'd3, 16'h40_00};
        18'd160: out = {16'd3, 16'h80_90};
        18'd161: out = {16'd3, 16'h40_00};
        18'd162: out = {16'd3, 16'h80_90};
        18'd163: out = {16'd3, 16'h40_00};
        18'd164: out = {16'd3, 16'h80_90};
        18'd165: out = {16'd3, 16'h40_00};
        18'd166: out = {16'd3, 16'h80_90};
        18'd167: out = {16'd3, 16'h40_00};
        18'd168: out = {16'd3, 16'h80_90};
        18'd169: out = {16'd3, 16'h40_00};
        18'd170: out = {16'd3, 16'h80_90};
        18'd171: out = {16'd3, 16'h40_00};
        18'd172: out = {16'd3, 16'h80_90};
        18'd173: out = {16'd3, 16'h40_00};
        18'd174: out = {16'd3, 16'h80_90};
        18'd175: out = {16'd3, 16'h40_00};
        18'd176: out = {16'd3, 16'h80_90};
        18'd177: out = {16'd3, 16'h40_00};
        18'd178: out = {16'd3, 16'h80_90};
        18'd179: out = {16'd3, 16'h40_00};
        18'd180: out = {16'd3, 16'h80_90};
        18'd181: out = {16'd3, 16'h40_00};
        18'd182: out = {16'd3, 16'h80_90};
        18'd183: out = {16'd3, 16'h40_00};
        18'd184: out = {16'd3, 16'h80_90};
        18'd185: out = {16'd3, 16'h40_00};
        18'd186: out = {16'd3, 16'h80_90};
        18'd187: out = {16'd3, 16'h40_00};
        18'd188: out = {16'd3, 16'h80_90};
        18'd189: out = {16'd3, 16'h40_00};
        18'd190: out = {16'd3, 16'h80_90};
        18'd191: out = {16'd3, 16'h40_00};
        18'd192: out = {16'd3, 16'h80_90};
        18'd193: out = {16'd3, 16'h40_00};
        18'd194: out = {16'd3, 16'h80_90};
        18'd195: out = {16'd3, 16'h40_00};
        18'd196: out = {16'd3, 16'h80_90};
        18'd197: out = {16'd3, 16'h40_00};
        18'd198: out = {16'd3, 16'h80_90};
        18'd199: out = {16'd3, 16'h40_00};
        18'd200: out = {16'd3, 16'h80_90};
        18'd201: out = {16'd3, 16'h40_00};
        18'd202: out = {16'd3, 16'h80_90};
        18'd203: out = {16'd3, 16'h40_00};
        18'd204: out = {16'd3, 16'h80_90};
        18'd205: out = {16'd3, 16'h40_00};
        18'd206: out = {16'd3, 16'h80_90};
        18'd207: out = {16'd3, 16'h40_00};
        18'd208: out = {16'd3, 16'h80_90};
        18'd209: out = {16'd3, 16'h40_00};
        18'd210: out = {16'd3, 16'h80_90};
        18'd211: out = {16'd3, 16'h40_00};
        18'd212: out = {16'd3, 16'h80_90};
        18'd213: out = {16'd3, 16'h40_00};
        18'd214: out = {16'd3, 16'h80_90};
        18'd215: out = {16'd3, 16'h40_00};
        18'd216: out = {16'd3, 16'h80_90};
        18'd217: out = {16'd3, 16'h40_00};
        18'd218: out = {16'd3, 16'h80_90};
        18'd219: out = {16'd3, 16'h40_00};
        18'd220: out = {16'd3, 16'h80_90};
        18'd221: out = {16'd3, 16'h40_00};
        18'd222: out = {16'd3, 16'h80_90};
        18'd223: out = {16'd3, 16'h40_00};
        18'd224: out = {16'd3, 16'h80_90};
        18'd225: out = {16'd3, 16'h40_00};
        18'd226: out = {16'd3, 16'h80_90};
        18'd227: out = {16'd3, 16'h40_00};
        18'd228: out = {16'd3, 16'h80_90};
        18'd229: out = {16'd3, 16'h40_00};
        18'd230: out = {16'd3, 16'h80_90};
        18'd231: out = {16'd3, 16'h40_00};
        18'd232: out = {16'd3, 16'h80_90};
        18'd233: out = {16'd3, 16'h40_00};
        18'd234: out = {16'd3, 16'h80_90};
        18'd235: out = {16'd3, 16'h40_00};
        18'd236: out = {16'd3, 16'h80_90};
        18'd237: out = {16'd3, 16'h40_00};
        18'd238: out = {16'd3, 16'h80_90};
        18'd239: out = {16'd3, 16'h40_00};
        18'd240: out = {16'd3, 16'h80_90};
        18'd241: out = {16'd3, 16'h40_00};
        18'd242: out = {16'd3, 16'h80_90};
        18'd243: out = {16'd3, 16'h40_00};
        18'd244: out = {16'd3, 16'h80_90};
        18'd245: out = {16'd3, 16'h40_00};
        18'd246: out = {16'd3, 16'h80_90};
        18'd247: out = {16'd3, 16'h40_00};
        18'd248: out = {16'd3, 16'h80_90};
        18'd249: out = {16'd3, 16'h40_00};
        18'd250: out = {16'd3, 16'h80_90};
        18'd251: out = {16'd3, 16'h40_00};
        18'd252: out = {16'd3, 16'h80_90};
        18'd253: out = {16'd3, 16'h40_00};
        18'd254: out = {16'd3, 16'h80_90};
        18'd255: out = {16'd3, 16'h40_00};
        18'd256: out = {16'd3, 16'h80_90};
        18'd257: out = {16'd3, 16'h40_00};
        18'd258: out = {16'd3, 16'h80_90};
        18'd259: out = {16'd3, 16'h40_00};
        18'd260: out = {16'd3, 16'h80_90};
        18'd261: out = {16'd3, 16'h40_00};
        18'd262: out = {16'd3, 16'h80_90};
        18'd263: out = {16'd3, 16'h40_00};
        18'd264: out = {16'd3, 16'h80_90};
        18'd265: out = {16'd3, 16'h40_00};
        18'd266: out = {16'd3, 16'h80_90};
        18'd267: out = {16'd3, 16'h40_00};
        18'd268: out = {16'd3, 16'h80_90};
        18'd269: out = {16'd3, 16'h40_00};
        18'd270: out = {16'd3, 16'h80_90};
        18'd271: out = {16'd3, 16'h40_00};
        18'd272: out = {16'd3, 16'h80_90};
        18'd273: out = {16'd3, 16'h40_00};
        18'd274: out = {16'd3, 16'h80_90};
        18'd275: out = {16'd3, 16'h40_00};
        18'd276: out = {16'd3, 16'h80_90};
        18'd277: out = {16'd3, 16'h40_00};
        18'd278: out = {16'd3, 16'h80_90};
        18'd279: out = {16'd3, 16'h40_00};
        18'd280: out = {16'd3, 16'h80_90};
        18'd281: out = {16'd3, 16'h40_00};
        18'd282: out = {16'd3, 16'h80_90};
        18'd283: out = {16'd3, 16'h40_00};
        18'd284: out = {16'd3, 16'h80_90};
        18'd285: out = {16'd3, 16'h40_00};
        18'd286: out = {16'd3, 16'h80_90};
        18'd287: out = {16'd3, 16'h40_00};
        18'd288: out = {16'd3, 16'h80_90};
        18'd289: out = {16'd3, 16'h40_00};
        18'd290: out = {16'd3, 16'h80_90};
        18'd291: out = {16'd3, 16'h40_00};
        18'd292: out = {16'd3, 16'h80_90};
        18'd293: out = {16'd3, 16'h40_00};
        18'd294: out = {16'd3, 16'h80_90};
        18'd295: out = {16'd3, 16'h40_00};
        18'd296: out = {16'd3, 16'h80_90};
        18'd297: out = {16'd3, 16'h40_00};
        18'd298: out = {16'd3, 16'h80_90};
        18'd299: out = {16'd3, 16'h40_00};
        18'd300: out = {16'd3, 16'h80_90};
        18'd301: out = {16'd3, 16'h40_00};
        18'd302: out = {16'd3, 16'h80_90};
        18'd303: out = {16'd3, 16'h40_00};
        18'd304: out = {16'd3, 16'h80_90};
        18'd305: out = {16'd3, 16'h40_00};
        18'd306: out = {16'd3, 16'h80_90};
        18'd307: out = {16'd3, 16'h40_00};
        18'd308: out = {16'd3, 16'h80_90};
        18'd309: out = {16'd3, 16'h40_00};
        18'd310: out = {16'd3, 16'h80_90};
        18'd311: out = {16'd3, 16'h40_00};
        18'd312: out = {16'd3, 16'h80_90};
        18'd313: out = {16'd3, 16'h40_00};
        18'd314: out = {16'd3, 16'h80_90};
        18'd315: out = {16'd3, 16'h40_00};
        18'd316: out = {16'd3, 16'h80_90};
        18'd317: out = {16'd3, 16'h40_00};
        18'd318: out = {16'd3, 16'h80_90};
        18'd319: out = {16'd3, 16'h40_00};
        18'd320: out = {16'd3, 16'h80_90};
        18'd321: out = {16'd3, 16'h40_00};
        18'd322: out = {16'd3, 16'h80_90};
        18'd323: out = {16'd3, 16'h40_00};
        18'd324: out = {16'd3, 16'h80_90};
        18'd325: out = {16'd3, 16'h40_00};
        18'd326: out = {16'd3, 16'h80_90};
        18'd327: out = {16'd3, 16'h40_00};
        18'd328: out = {16'd3, 16'h80_90};
        18'd329: out = {16'd3, 16'h40_00};
        18'd330: out = {16'd3, 16'h80_90};
        18'd331: out = {16'd3, 16'h40_00};
        18'd332: out = {16'd3, 16'h80_90};
        18'd333: out = {16'd3, 16'h40_00};
        18'd334: out = {16'd3, 16'h80_90};
        18'd335: out = {16'd3, 16'h40_00};
        18'd336: out = {16'd3, 16'h80_90};
        18'd337: out = {16'd3, 16'h40_00};
        18'd338: out = {16'd3, 16'h80_90};
        18'd339: out = {16'd3, 16'h40_00};
        18'd340: out = {16'd3, 16'h80_90};
        18'd341: out = {16'd3, 16'h40_00};
        18'd342: out = {16'd3, 16'h80_90};
        18'd343: out = {16'd3, 16'h40_00};
        18'd344: out = {16'd3, 16'h80_90};
        18'd345: out = {16'd3, 16'h40_00};
        18'd346: out = {16'd3, 16'h80_90};
        18'd347: out = {16'd3, 16'h40_00};
        18'd348: out = {16'd3, 16'h80_90};
        18'd349: out = {16'd3, 16'h40_00};
        18'd350: out = {16'd3, 16'h80_90};
        18'd351: out = {16'd3, 16'h40_00};
        18'd352: out = {16'd3, 16'h80_90};
        18'd353: out = {16'd3, 16'h40_00};
        18'd354: out = {16'd3, 16'h80_90};
        18'd355: out = {16'd3, 16'h40_00};
        18'd356: out = {16'd3, 16'h80_90};
        18'd357: out = {16'd3, 16'h40_00};
        18'd358: out = {16'd3, 16'h80_90};
        18'd359: out = {16'd3, 16'h40_00};
        18'd360: out = {16'd3, 16'h80_90};
        18'd361: out = {16'd3, 16'h40_00};
        18'd362: out = {16'd3, 16'h80_90};
        18'd363: out = {16'd3, 16'h40_00};
        18'd364: out = {16'd3, 16'h80_90};
        18'd365: out = {16'd3, 16'h40_00};
        18'd366: out = {16'd3, 16'h80_90};
        18'd367: out = {16'd3, 16'h40_00};
        18'd368: out = {16'd3, 16'h80_90};
        18'd369: out = {16'd3, 16'h40_00};
        18'd370: out = {16'd3, 16'h80_90};
        18'd371: out = {16'd3, 16'h40_00};
        18'd372: out = {16'd3, 16'h80_90};
        18'd373: out = {16'd3, 16'h40_00};
        18'd374: out = {16'd3, 16'h80_90};
        18'd375: out = {16'd3, 16'h40_00};
        18'd376: out = {16'd3, 16'h80_90};
        18'd377: out = {16'd3, 16'h40_00};
        18'd378: out = {16'd3, 16'h80_90};
        18'd379: out = {16'd3, 16'h40_00};
        18'd380: out = {16'd3, 16'h80_90};
        18'd381: out = {16'd3, 16'h40_00};
        18'd382: out = {16'd3, 16'h80_90};
        18'd383: out = {16'd3, 16'h40_00};
        18'd384: out = {16'd3, 16'h80_90};
        18'd385: out = {16'd3, 16'h40_00};
        18'd386: out = {16'd3, 16'h80_90};
        18'd387: out = {16'd3, 16'h40_00};
        18'd388: out = {16'd3, 16'h80_90};
        18'd389: out = {16'd3, 16'h40_00};
        18'd390: out = {16'd3, 16'h80_90};
        18'd391: out = {16'd3, 16'h40_00};
        18'd392: out = {16'd3, 16'h80_90};
        18'd393: out = {16'd3, 16'h40_00};
        18'd394: out = {16'd3, 16'h80_90};
        18'd395: out = {16'd3, 16'h40_00};
        18'd396: out = {16'd3, 16'h80_90};
        18'd397: out = {16'd3, 16'h40_00};
        18'd398: out = {16'd3, 16'h80_90};
        18'd399: out = {16'd3, 16'h40_00};
        18'd400: out = {16'd3, 16'h80_90};
        18'd401: out = {16'd3, 16'h40_00};
        18'd402: out = {16'd3, 16'h80_90};
        18'd403: out = {16'd3, 16'h40_00};
        18'd404: out = {16'd3, 16'h80_90};
        18'd405: out = {16'd3, 16'h40_00};
        18'd406: out = {16'd3, 16'h80_90};
        18'd407: out = {16'd3, 16'h40_00};
        18'd408: out = {16'd3, 16'h80_90};
        18'd409: out = {16'd3, 16'h40_00};
        18'd410: out = {16'd3, 16'h80_90};
        18'd411: out = {16'd3, 16'h40_00};
        18'd412: out = {16'd3, 16'h80_90};
        18'd413: out = {16'd3, 16'h40_00};
        18'd414: out = {16'd3, 16'h80_90};
        18'd415: out = {16'd3, 16'h40_00};
        18'd416: out = {16'd3, 16'h80_90};
        18'd417: out = {16'd3, 16'h40_00};
        18'd418: out = {16'd3, 16'h80_90};
        18'd419: out = {16'd3, 16'h40_00};
        18'd420: out = {16'd3, 16'h80_90};
        18'd421: out = {16'd3, 16'h40_00};
        18'd422: out = {16'd3, 16'h80_90};
        18'd423: out = {16'd3, 16'h40_00};
        18'd424: out = {16'd3, 16'h80_90};
        18'd425: out = {16'd3, 16'h40_00};
        18'd426: out = {16'd3, 16'h80_90};
        18'd427: out = {16'd3, 16'h40_00};
        18'd428: out = {16'd3, 16'h80_90};
        18'd429: out = {16'd3, 16'h40_00};
        18'd430: out = {16'd3, 16'h80_90};
        18'd431: out = {16'd3, 16'h40_00};
        18'd432: out = {16'd3, 16'h80_90};
        18'd433: out = {16'd3, 16'h40_00};
        18'd434: out = {16'd3, 16'h80_90};
        18'd435: out = {16'd3, 16'h40_00};
        18'd436: out = {16'd3, 16'h80_90};
        18'd437: out = {16'd3, 16'h40_00};
        18'd438: out = {16'd3, 16'h80_90};
        18'd439: out = {16'd3, 16'h40_00};
        18'd440: out = {16'd3, 16'h80_90};
        18'd441: out = {16'd3, 16'h40_00};
        18'd442: out = {16'd3, 16'h80_90};
        18'd443: out = {16'd3, 16'h40_00};
        18'd444: out = {16'd3, 16'h80_90};
        18'd445: out = {16'd3, 16'h40_00};
        18'd446: out = {16'd3, 16'h80_90};
        18'd447: out = {16'd3, 16'h40_00};
        18'd448: out = {16'd3, 16'h80_90};
        18'd449: out = {16'd3, 16'h40_00};
        18'd450: out = {16'd3, 16'h80_90};
        18'd451: out = {16'd3, 16'h40_00};
        18'd452: out = {16'd3, 16'h80_90};
        18'd453: out = {16'd3, 16'h40_00};
        18'd454: out = {16'd3, 16'h80_90};
        18'd455: out = {16'd3, 16'h40_00};
        18'd456: out = {16'd3, 16'h80_90};
        18'd457: out = {16'd3, 16'h40_00};
        18'd458: out = {16'd3, 16'h80_90};
        18'd459: out = {16'd3, 16'h40_00};
        18'd460: out = {16'd3, 16'h80_90};
        18'd461: out = {16'd3, 16'h40_00};
        18'd462: out = {16'd3, 16'h80_90};
        18'd463: out = {16'd3, 16'h40_00};
        18'd464: out = {16'd3, 16'h80_90};
        18'd465: out = {16'd3, 16'h40_00};
        18'd466: out = {16'd3, 16'h80_90};
        18'd467: out = {16'd3, 16'h40_00};
        18'd468: out = {16'd3, 16'h80_90};
        18'd469: out = {16'd3, 16'h40_00};
        18'd470: out = {16'd3, 16'h80_90};
        18'd471: out = {16'd3, 16'h40_00};
        18'd472: out = {16'd3, 16'h80_90};
        18'd473: out = {16'd3, 16'h40_00};
        18'd474: out = {16'd3, 16'h80_90};
        18'd475: out = {16'd3, 16'h40_00};
        18'd476: out = {16'd3, 16'h80_90};
        18'd477: out = {16'd3, 16'h40_00};
        18'd478: out = {16'd3, 16'h80_90};
        18'd479: out = {16'd3, 16'h40_00};
        18'd480: out = {16'd3, 16'h80_90};
        18'd481: out = {16'd3, 16'h40_00};
        18'd482: out = {16'd3, 16'h80_90};
        18'd483: out = {16'd3, 16'h40_00};
        18'd484: out = {16'd3, 16'h80_90};
        18'd485: out = {16'd3, 16'h40_00};
        18'd486: out = {16'd3, 16'h80_90};
        18'd487: out = {16'd3, 16'h40_00};
        18'd488: out = {16'd3, 16'h80_90};
        18'd489: out = {16'd3, 16'h40_00};
        18'd490: out = {16'd3, 16'h80_90};
        18'd491: out = {16'd3, 16'h40_00};
        18'd492: out = {16'd3, 16'h80_90};
        18'd493: out = {16'd3, 16'h40_00};
        18'd494: out = {16'd3, 16'h80_90};
        18'd495: out = {16'd3, 16'h40_00};
        18'd496: out = {16'd3, 16'h80_90};
        18'd497: out = {16'd3, 16'h40_00};
        18'd498: out = {16'd3, 16'h80_90};
        18'd499: out = {16'd3, 16'h40_00};
        18'd500: out = {16'd3, 16'h80_90};
        18'd501: out = {16'd3, 16'h40_00};
        18'd502: out = {16'd3, 16'h80_90};
        18'd503: out = {16'd3, 16'h40_00};
        18'd504: out = {16'd3, 16'h80_90};
        18'd505: out = {16'd3, 16'h40_00};
        18'd506: out = {16'd3, 16'h80_90};
        18'd507: out = {16'd3, 16'h40_00};
        18'd508: out = {16'd3, 16'h80_90};
        18'd509: out = {16'd3, 16'h40_00};
        18'd510: out = {16'd3, 16'h80_90};
        18'd511: out = {16'd3, 16'h40_00};
        18'd512: out = {16'd3, 16'h80_90};
        18'd513: out = {16'd3, 16'h40_00};
        18'd514: out = {16'd3, 16'h80_90};
        18'd515: out = {16'd3, 16'h40_00};
        18'd516: out = {16'd3, 16'h80_90};
        18'd517: out = {16'd3, 16'h40_00};
        18'd518: out = {16'd3, 16'h80_90};
        18'd519: out = {16'd3, 16'h40_00};
        18'd520: out = {16'd3, 16'h80_90};
        18'd521: out = {16'd3, 16'h40_00};
        18'd522: out = {16'd3, 16'h80_90};
        18'd523: out = {16'd3, 16'h40_00};
        18'd524: out = {16'd3, 16'h80_90};
        18'd525: out = {16'd3, 16'h40_00};
        18'd526: out = {16'd3, 16'h80_90};
        18'd527: out = {16'd3, 16'h40_00};
        18'd528: out = {16'd3, 16'h80_90};
        18'd529: out = {16'd3, 16'h40_00};
        18'd530: out = {16'd3, 16'h80_90};
        18'd531: out = {16'd3, 16'h80_90};
        18'd532: out = {16'd3, 16'h80_90};
        18'd533: out = {16'd3, 16'h40_00};
        18'd534: out = {16'd3, 16'h80_90};
        18'd535: out = {16'd3, 16'h40_00};
        18'd536: out = {16'd3, 16'h80_90};
        18'd537: out = {16'd3, 16'h40_00};
        18'd538: out = {16'd3, 16'h80_90};
        18'd539: out = {16'd3, 16'h40_00};
        18'd540: out = {16'd3, 16'h80_90};
        18'd541: out = {16'd3, 16'h40_00};
        18'd542: out = {16'd3, 16'h80_90};
        18'd543: out = {16'd3, 16'h40_00};
        18'd544: out = {16'd3, 16'h80_90};
        18'd545: out = {16'd3, 16'h40_00};
        18'd546: out = {16'd3, 16'h80_90};
        18'd547: out = {16'd3, 16'h40_00};
        18'd548: out = {16'd3, 16'h80_90};
        18'd549: out = {16'd3, 16'h40_00};
        18'd550: out = {16'd3, 16'h80_90};
        18'd551: out = {16'd3, 16'h40_00};
        18'd552: out = {16'd3, 16'h80_90};
        18'd553: out = {16'd3, 16'h40_00};
        18'd554: out = {16'd3, 16'h80_90};
        18'd555: out = {16'd3, 16'h40_00};
        18'd556: out = {16'd3, 16'h80_90};
        18'd557: out = {16'd3, 16'h40_00};
        18'd558: out = {16'd3, 16'h80_90};
        18'd559: out = {16'd3, 16'h40_00};
        18'd560: out = {16'd3, 16'h80_90};
        18'd561: out = {16'd3, 16'h40_00};
        18'd562: out = {16'd3, 16'h80_90};
        18'd563: out = {16'd3, 16'h40_00};
        18'd564: out = {16'd3, 16'h80_90};
        18'd565: out = {16'd3, 16'h40_00};
        18'd566: out = {16'd3, 16'h80_90};
        18'd567: out = {16'd3, 16'h40_00};
        18'd568: out = {16'd3, 16'h80_90};
        18'd569: out = {16'd3, 16'h40_00};
        18'd570: out = {16'd3, 16'h80_90};
        18'd571: out = {16'd3, 16'h40_00};
        18'd572: out = {16'd3, 16'h80_90};
        18'd573: out = {16'd3, 16'h40_00};
        18'd574: out = {16'd3, 16'h80_90};
        18'd575: out = {16'd3, 16'h40_00};
        18'd576: out = {16'd3, 16'h80_90};
        18'd577: out = {16'd3, 16'h40_00};
        18'd578: out = {16'd3, 16'h80_90};
        18'd579: out = {16'd3, 16'h40_00};
        18'd580: out = {16'd3, 16'h80_90};
        18'd581: out = {16'd3, 16'h40_00};
        18'd582: out = {16'd3, 16'h80_90};
        18'd583: out = {16'd3, 16'h40_00};
        18'd584: out = {16'd3, 16'h80_90};
        18'd585: out = {16'd3, 16'h40_00};
        18'd586: out = {16'd3, 16'h80_90};
        18'd587: out = {16'd3, 16'h40_00};
        18'd588: out = {16'd3, 16'h80_90};
        18'd589: out = {16'd3, 16'h40_00};
        18'd590: out = {16'd3, 16'h80_90};
        18'd591: out = {16'd3, 16'h40_00};
        18'd592: out = {16'd3, 16'h80_90};
        18'd593: out = {16'd3, 16'h40_00};
        18'd594: out = {16'd3, 16'h80_90};
        18'd595: out = {16'd3, 16'h40_00};
        18'd596: out = {16'd3, 16'h80_90};
        18'd597: out = {16'd3, 16'h40_00};
        18'd598: out = {16'd3, 16'h80_90};
        18'd599: out = {16'd3, 16'h40_00};
        18'd600: out = {16'd3, 16'h80_90};
        18'd601: out = {16'd3, 16'h40_00};
        18'd602: out = {16'd3, 16'h80_90};
        18'd603: out = {16'd3, 16'h40_00};
        18'd604: out = {16'd3, 16'h80_90};
        18'd605: out = {16'd3, 16'h40_00};
        18'd606: out = {16'd3, 16'h80_90};
        18'd607: out = {16'd3, 16'h40_00};
        18'd608: out = {16'd3, 16'h80_90};
        18'd609: out = {16'd3, 16'h40_00};
        18'd610: out = {16'd3, 16'h80_90};
        18'd611: out = {16'd3, 16'h40_00};
        18'd612: out = {16'd3, 16'h80_90};
        18'd613: out = {16'd3, 16'h40_00};
        18'd614: out = {16'd3, 16'h80_90};
        18'd615: out = {16'd3, 16'h40_00};
        18'd616: out = {16'd3, 16'h80_90};
        18'd617: out = {16'd3, 16'h40_00};
        18'd618: out = {16'd3, 16'h80_90};
        18'd619: out = {16'd3, 16'h40_00};
        18'd620: out = {16'd3, 16'h80_90};
        18'd621: out = {16'd3, 16'h40_00};
        18'd622: out = {16'd3, 16'h80_90};
        18'd623: out = {16'd3, 16'h40_00};
        18'd624: out = {16'd3, 16'h80_90};
        18'd625: out = {16'd3, 16'h40_00};
        18'd626: out = {16'd3, 16'h80_90};
        18'd627: out = {16'd3, 16'h40_00};
        18'd628: out = {16'd3, 16'h80_90};
        18'd629: out = {16'd3, 16'h40_00};
        18'd630: out = {16'd3, 16'h80_90};
        18'd631: out = {16'd3, 16'h40_00};
        18'd632: out = {16'd3, 16'h80_90};
        18'd633: out = {16'd3, 16'h40_00};
        18'd634: out = {16'd3, 16'h80_90};
        18'd635: out = {16'd3, 16'h40_00};
        18'd636: out = {16'd3, 16'h80_90};
        18'd637: out = {16'd3, 16'h40_00};
        18'd638: out = {16'd3, 16'h80_90};
        18'd639: out = {16'd3, 16'h40_00};
        18'd640: out = {16'd3, 16'h80_90};
        18'd641: out = {16'd3, 16'h40_00};
        18'd642: out = {16'd3, 16'h80_90};
        18'd643: out = {16'd3, 16'h40_00};
        18'd644: out = {16'd3, 16'h80_90};
        18'd645: out = {16'd3, 16'h40_00};
        18'd646: out = {16'd3, 16'h80_90};
        18'd647: out = {16'd3, 16'h40_00};
        18'd648: out = {16'd3, 16'h80_90};
        18'd649: out = {16'd3, 16'h40_00};
        18'd650: out = {16'd3, 16'h80_90};
        18'd651: out = {16'd3, 16'h40_00};
        18'd652: out = {16'd3, 16'h80_90};
        18'd653: out = {16'd3, 16'h40_00};
        18'd654: out = {16'd3, 16'h80_90};
        18'd655: out = {16'd3, 16'h40_00};
        18'd656: out = {16'd3, 16'h80_90};
        18'd657: out = {16'd3, 16'h40_00};
        18'd658: out = {16'd3, 16'h80_90};
        18'd659: out = {16'd3, 16'h40_00};
        18'd670: out = {16'd3, 16'h80_90};
        18'd671: out = {16'd3, 16'h40_00};
        18'd672: out = {16'd3, 16'h80_90};
        18'd673: out = {16'd3, 16'h40_00};
        18'd674: out = {16'd3, 16'h80_90};
        18'd675: out = {16'd3, 16'h40_00};
        18'd676: out = {16'd3, 16'h80_90};
        18'd677: out = {16'd3, 16'h40_00};
        18'd678: out = {16'd3, 16'h80_90};
        18'd679: out = {16'd3, 16'h40_00};
        18'd680: out = {16'd3, 16'h80_90};
        18'd681: out = {16'd3, 16'h40_00};
        18'd682: out = {16'd3, 16'h80_90};
        18'd683: out = {16'd3, 16'h40_00};
        18'd684: out = {16'd3, 16'h80_90};
        18'd685: out = {16'd3, 16'h40_00};
        18'd686: out = {16'd3, 16'h80_90};
        18'd687: out = {16'd3, 16'h40_00};
        18'd688: out = {16'd3, 16'h80_90};
        18'd689: out = {16'd3, 16'h40_00};
        18'd690: out = {16'd3, 16'h80_90};
        18'd691: out = {16'd3, 16'h40_00};
        18'd692: out = {16'd3, 16'h80_90};
        18'd693: out = {16'd3, 16'h40_00};
        18'd694: out = {16'd3, 16'h80_90};
        18'd695: out = {16'd3, 16'h40_00};
        18'd696: out = {16'd3, 16'h80_90};
        18'd697: out = {16'd3, 16'h40_00};
        18'd698: out = {16'd3, 16'h80_90};
        18'd699: out = {16'd3, 16'h40_00};
        18'd700: out = {16'd3, 16'h80_90};
        18'd701: out = {16'd3, 16'h40_00};
        18'd702: out = {16'd3, 16'h80_90};
        18'd703: out = {16'd3, 16'h40_00};
        18'd704: out = {16'd3, 16'h80_90};
        18'd705: out = {16'd3, 16'h40_00};
        18'd706: out = {16'd3, 16'h80_40};
        18'd707: out = {16'd3, 16'h40_00};
        18'd708: out = {16'd3, 16'h00_00};
        18'd709: out = {16'd3, 16'h80_99};
        18'd710: out = {16'd3, 16'h00_90};
        18'd711: out = {16'd3, 16'h80_9A};
        18'd712: out = {16'd3, 16'h00_01};
        18'd713: out = {16'd3, 16'h80_9B};
        18'd714: out = {16'd3, 16'h00_F0};
        18'd715: out = {16'd3, 16'h80_9C};
        18'd716: out = {16'd3, 16'h00_00};
        18'd717: out = {16'd3, 16'h80_9D};
        18'd718: out = {16'd3, 16'h00_32};
        18'd719: out = {16'd3, 16'h80_63};
        18'd720: out = {16'd3, 16'h00_1F};
        18'd721: out = {16'd3, 16'h80_64};
        18'd722: out = {16'd3, 16'h00_00};
        18'd723: out = {16'd3, 16'h80_65};
        18'd724: out = {16'd3, 16'h00_1F};
        18'd725: out = {16'd3, 16'h80_90};
        18'd726: out = {16'd3, 16'h00_60};
        18'd727: out = {16'd3, 16'h80_90};
        18'd728: out = {16'd3, 16'h40_00};
        18'd729: out = {16'd3, 16'h80_90};
        18'd730: out = {16'd3, 16'h40_00};
        18'd731: out = {16'd3, 16'h80_90};
        18'd732: out = {16'd3, 16'h40_00};
        18'd733: out = {16'd3, 16'h80_90};
        18'd734: out = {16'd3, 16'h40_00};
        18'd735: out = {16'd3, 16'h80_90};
        18'd736: out = {16'd3, 16'h40_00};
        18'd737: out = {16'd3, 16'h80_90};
        18'd738: out = {16'd3, 16'h40_00};
        18'd739: out = {16'd3, 16'h80_90};
        18'd740: out = {16'd3, 16'h40_00};
        18'd741: out = {16'd3, 16'h80_90};
        18'd742: out = {16'd3, 16'h40_00};
        18'd743: out = {16'd3, 16'h80_90};
        18'd744: out = {16'd3, 16'h40_00};
        18'd745: out = {16'd3, 16'h80_90};
        18'd746: out = {16'd3, 16'h40_00};
        18'd747: out = {16'd3, 16'h80_90};
        18'd748: out = {16'd3, 16'h40_00};
        18'd749: out = {16'd3, 16'h80_90};
        18'd750: out = {16'd3, 16'h40_00};
        18'd751: out = {16'd3, 16'h80_90};
        18'd752: out = {16'd3, 16'h40_00};
        18'd753: out = {16'd3, 16'h80_90};
        18'd754: out = {16'd3, 16'h40_00};
        18'd755: out = {16'd3, 16'h80_90};
        18'd756: out = {16'd3, 16'h40_00};
        18'd757: out = {16'd3, 16'h80_90};
        18'd758: out = {16'd3, 16'h40_00};
        18'd759: out = {16'd3, 16'h80_90};
        18'd760: out = {16'd3, 16'h40_00};
        18'd761: out = {16'd3, 16'h80_90};
        18'd762: out = {16'd3, 16'h40_00};
        18'd763: out = {16'd3, 16'h80_90};
        18'd764: out = {16'd3, 16'h40_00};
        18'd765: out = {16'd3, 16'h80_90};
        18'd766: out = {16'd3, 16'h40_00};
        18'd767: out = {16'd3, 16'h80_90};
        18'd768: out = {16'd3, 16'h40_00};
        18'd769: out = {16'd3, 16'h80_90};
        18'd770: out = {16'd3, 16'h40_00};
        18'd771: out = {16'd3, 16'h80_90};
        18'd772: out = {16'd3, 16'h40_00};
        18'd773: out = {16'd3, 16'h80_90};
        18'd774: out = {16'd3, 16'h40_00};
        18'd775: out = {16'd3, 16'h80_90};
        18'd776: out = {16'd3, 16'h40_00};
        18'd777: out = {16'd3, 16'h80_90};
        18'd778: out = {16'd3, 16'h40_00};
        18'd779: out = {16'd3, 16'h80_90};
        18'd780: out = {16'd3, 16'h40_00};
        18'd781: out = {16'd3, 16'h80_90};
        18'd782: out = {16'd3, 16'h40_00};
        18'd783: out = {16'd3, 16'h80_90};
        18'd784: out = {16'd3, 16'h40_00};
        18'd785: out = {16'd3, 16'h80_90};
        18'd786: out = {16'd3, 16'h40_00};
        18'd787: out = {16'd3, 16'h80_90};
        18'd788: out = {16'd3, 16'h40_00};
        18'd789: out = {16'd3, 16'h80_90};
        18'd790: out = {16'd3, 16'h40_00};
        18'd791: out = {16'd3, 16'h80_90};
        18'd792: out = {16'd3, 16'h40_00};
        18'd793: out = {16'd3, 16'h80_90};
        18'd794: out = {16'd3, 16'h40_00};
        18'd795: out = {16'd3, 16'h80_90};
        18'd796: out = {16'd3, 16'h40_00};
        18'd797: out = {16'd3, 16'h80_90};
        18'd798: out = {16'd3, 16'h40_00};
        18'd799: out = {16'd3, 16'h80_90};
        18'd800: out = {16'd3, 16'h40_00};
        18'd801: out = {16'd3, 16'h80_90};
        18'd802: out = {16'd3, 16'h40_00};
        18'd803: out = {16'd3, 16'h80_90};
        18'd804: out = {16'd3, 16'h40_00};
        18'd805: out = {16'd3, 16'h80_90};
        18'd806: out = {16'd3, 16'h40_00};
        18'd807: out = {16'd3, 16'h80_90};
        18'd808: out = {16'd3, 16'h40_00};
        18'd809: out = {16'd3, 16'h80_90};
        18'd810: out = {16'd3, 16'h40_00};
        18'd811: out = {16'd3, 16'h80_90};
        18'd812: out = {16'd3, 16'h40_00};
        18'd813: out = {16'd3, 16'h80_90};
        18'd814: out = {16'd3, 16'h40_00};
        18'd815: out = {16'd3, 16'h80_90};
        18'd816: out = {16'd3, 16'h40_00};
        18'd817: out = {16'd3, 16'h80_90};
        18'd818: out = {16'd3, 16'h40_00};
        18'd819: out = {16'd3, 16'h80_90};
        18'd820: out = {16'd3, 16'h40_00};
        18'd821: out = {16'd3, 16'h80_90};
        18'd822: out = {16'd3, 16'h40_00};
        18'd823: out = {16'd3, 16'h80_90};
        18'd824: out = {16'd3, 16'h40_00};
        18'd825: out = {16'd3, 16'h80_90};
        18'd826: out = {16'd3, 16'h40_00};
        18'd827: out = {16'd3, 16'h80_90};
        18'd828: out = {16'd3, 16'h40_00};
        18'd829: out = {16'd3, 16'h80_90};
        18'd830: out = {16'd3, 16'h40_00};
        18'd831: out = {16'd3, 16'h80_90};
        18'd832: out = {16'd3, 16'h40_00};
        18'd833: out = {16'd3, 16'h80_90};
        18'd834: out = {16'd3, 16'h40_00};
        18'd835: out = {16'd3, 16'h80_90};
        18'd836: out = {16'd3, 16'h40_00};
        18'd837: out = {16'd3, 16'h80_90};
        18'd838: out = {16'd3, 16'h40_00};
        18'd839: out = {16'd3, 16'h80_90};
        18'd840: out = {16'd3, 16'h40_00};
        18'd841: out = {16'd3, 16'h80_90};
        18'd842: out = {16'd3, 16'h40_00};
        18'd843: out = {16'd3, 16'h80_90};
        18'd844: out = {16'd3, 16'h40_00};
        18'd845: out = {16'd3, 16'h80_90};
        18'd846: out = {16'd3, 16'h40_00};
        
        default: begin
            // delay = 1;
            out = '0;
        end 
    endcase
  end
endmodule





        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_40};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h00_00};
        // 18'd: out = {16'd3, 16'h80_99};
        // 18'd: out = {16'd3, 16'h00_90};
        // 18'd: out = {16'd3, 16'h80_9A};
        // 18'd: out = {16'd3, 16'h00_01};
        // 18'd: out = {16'd3, 16'h80_9B};
        // 18'd: out = {16'd3, 16'h00_F0};
        // 18'd: out = {16'd3, 16'h80_9C};
        // 18'd: out = {16'd3, 16'h00_00};
        // 18'd: out = {16'd3, 16'h80_9D};
        // 18'd: out = {16'd3, 16'h00_32};
        // 18'd: out = {16'd3, 16'h80_63};
        // 18'd: out = {16'd3, 16'h00_1F};
        // 18'd: out = {16'd3, 16'h80_64};
        // 18'd: out = {16'd3, 16'h00_00};
        // 18'd: out = {16'd3, 16'h80_65};
        // 18'd: out = {16'd3, 16'h00_1F};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h00_60};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};
        // 18'd: out = {16'd3, 16'h80_90};
        // 18'd: out = {16'd3, 16'h40_00};


